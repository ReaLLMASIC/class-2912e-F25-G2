magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< metal1 >>
rect -44 11968 200 12000
rect -44 11916 0 11968
rect 156 11916 200 11968
rect -44 11844 200 11916
rect -44 11792 0 11844
rect 156 11792 200 11844
rect -44 11720 200 11792
rect -44 11668 0 11720
rect 156 11668 200 11720
rect -44 11596 200 11668
rect -44 11544 0 11596
rect 156 11544 200 11596
rect -44 11472 200 11544
rect -44 11420 0 11472
rect 156 11420 200 11472
rect -44 11348 200 11420
rect -44 11296 0 11348
rect 156 11296 200 11348
rect -44 11224 200 11296
rect -44 11172 0 11224
rect 156 11172 200 11224
rect -44 11100 200 11172
rect -44 11048 0 11100
rect 156 11048 200 11100
rect -44 10976 200 11048
rect -44 10924 0 10976
rect 156 10924 200 10976
rect -44 10852 200 10924
rect -44 10800 0 10852
rect 156 10800 200 10852
rect -44 10728 200 10800
rect -44 10676 0 10728
rect 156 10676 200 10728
rect -44 10604 200 10676
rect -44 10552 0 10604
rect 156 10552 200 10604
rect -44 10480 200 10552
rect -44 10428 0 10480
rect 156 10428 200 10480
rect -44 10356 200 10428
rect -44 10304 0 10356
rect 156 10304 200 10356
rect -44 10232 200 10304
rect -44 10180 0 10232
rect 156 10180 200 10232
rect -44 10108 200 10180
rect -44 10056 0 10108
rect 156 10056 200 10108
rect -44 9984 200 10056
rect -44 9932 0 9984
rect 156 9932 200 9984
rect -44 9860 200 9932
rect -44 9808 0 9860
rect 156 9808 200 9860
rect -44 9736 200 9808
rect -44 9684 0 9736
rect 156 9684 200 9736
rect -44 9612 200 9684
rect -44 9560 0 9612
rect 156 9560 200 9612
rect -44 9488 200 9560
rect -44 9436 0 9488
rect 156 9436 200 9488
rect -44 9364 200 9436
rect -44 9312 0 9364
rect 156 9312 200 9364
rect -44 9240 200 9312
rect -44 9188 0 9240
rect 156 9188 200 9240
rect -44 9116 200 9188
rect -44 9064 0 9116
rect 156 9064 200 9116
rect -44 8992 200 9064
rect -44 8940 0 8992
rect 156 8940 200 8992
rect -44 8868 200 8940
rect -44 8816 0 8868
rect 156 8816 200 8868
rect -44 8744 200 8816
rect -44 8692 0 8744
rect 156 8692 200 8744
rect -44 8620 200 8692
rect -44 8568 0 8620
rect 156 8568 200 8620
rect -44 8496 200 8568
rect -44 8444 0 8496
rect 156 8444 200 8496
rect -44 8372 200 8444
rect -44 8320 0 8372
rect 156 8320 200 8372
rect -44 8248 200 8320
rect -44 8196 0 8248
rect 156 8196 200 8248
rect -44 8124 200 8196
rect -44 8072 0 8124
rect 156 8072 200 8124
rect -44 8000 200 8072
rect -44 7948 0 8000
rect 156 7948 200 8000
rect -44 7876 200 7948
rect -44 7824 0 7876
rect 156 7824 200 7876
rect -44 7752 200 7824
rect -44 7700 0 7752
rect 156 7700 200 7752
rect -44 7628 200 7700
rect -44 7576 0 7628
rect 156 7576 200 7628
rect -44 7504 200 7576
rect -44 7452 0 7504
rect 156 7452 200 7504
rect -44 7380 200 7452
rect -44 7328 0 7380
rect 156 7328 200 7380
rect -44 7256 200 7328
rect -44 7204 0 7256
rect 156 7204 200 7256
rect -44 7132 200 7204
rect -44 7080 0 7132
rect 156 7080 200 7132
rect -44 7008 200 7080
rect -44 6956 0 7008
rect 156 6956 200 7008
rect -44 6884 200 6956
rect -44 6832 0 6884
rect 156 6832 200 6884
rect -44 6760 200 6832
rect -44 6708 0 6760
rect 156 6708 200 6760
rect -44 6636 200 6708
rect -44 6584 0 6636
rect 156 6584 200 6636
rect -44 6512 200 6584
rect -44 6460 0 6512
rect 156 6460 200 6512
rect -44 6388 200 6460
rect -44 6336 0 6388
rect 156 6336 200 6388
rect -44 6264 200 6336
rect -44 6212 0 6264
rect 156 6212 200 6264
rect -44 6140 200 6212
rect -44 6088 0 6140
rect 156 6088 200 6140
rect -44 6016 200 6088
rect -44 5964 0 6016
rect 156 5964 200 6016
rect -44 5892 200 5964
rect -44 5840 0 5892
rect 156 5840 200 5892
rect -44 5768 200 5840
rect -44 5716 0 5768
rect 156 5716 200 5768
rect -44 5644 200 5716
rect -44 5592 0 5644
rect 156 5592 200 5644
rect -44 5520 200 5592
rect -44 5468 0 5520
rect 156 5468 200 5520
rect -44 5396 200 5468
rect -44 5344 0 5396
rect 156 5344 200 5396
rect -44 5272 200 5344
rect -44 5220 0 5272
rect 156 5220 200 5272
rect -44 5148 200 5220
rect -44 5096 0 5148
rect 156 5096 200 5148
rect -44 5024 200 5096
rect -44 4972 0 5024
rect 156 4972 200 5024
rect -44 4900 200 4972
rect -44 4848 0 4900
rect 156 4848 200 4900
rect -44 4776 200 4848
rect -44 4724 0 4776
rect 156 4724 200 4776
rect -44 4652 200 4724
rect -44 4600 0 4652
rect 156 4600 200 4652
rect -44 4528 200 4600
rect -44 4476 0 4528
rect 156 4476 200 4528
rect -44 4404 200 4476
rect -44 4352 0 4404
rect 156 4352 200 4404
rect -44 4280 200 4352
rect -44 4228 0 4280
rect 156 4228 200 4280
rect -44 4156 200 4228
rect -44 4104 0 4156
rect 156 4104 200 4156
rect -44 4032 200 4104
rect -44 3980 0 4032
rect 156 3980 200 4032
rect -44 3908 200 3980
rect -44 3856 0 3908
rect 156 3856 200 3908
rect -44 3784 200 3856
rect -44 3732 0 3784
rect 156 3732 200 3784
rect -44 3660 200 3732
rect -44 3608 0 3660
rect 156 3608 200 3660
rect -44 3536 200 3608
rect -44 3484 0 3536
rect 156 3484 200 3536
rect -44 3412 200 3484
rect -44 3360 0 3412
rect 156 3360 200 3412
rect -44 3288 200 3360
rect -44 3236 0 3288
rect 156 3236 200 3288
rect -44 3164 200 3236
rect -44 3112 0 3164
rect 156 3112 200 3164
rect -44 3040 200 3112
rect -44 2988 0 3040
rect 156 2988 200 3040
rect -44 2916 200 2988
rect -44 2864 0 2916
rect 156 2864 200 2916
rect -44 2792 200 2864
rect -44 2740 0 2792
rect 156 2740 200 2792
rect -44 2668 200 2740
rect -44 2616 0 2668
rect 156 2616 200 2668
rect -44 2544 200 2616
rect -44 2492 0 2544
rect 156 2492 200 2544
rect -44 2420 200 2492
rect -44 2368 0 2420
rect 156 2368 200 2420
rect -44 2296 200 2368
rect -44 2244 0 2296
rect 156 2244 200 2296
rect -44 2172 200 2244
rect -44 2120 0 2172
rect 156 2120 200 2172
rect -44 2048 200 2120
rect -44 1996 0 2048
rect 156 1996 200 2048
rect -44 1924 200 1996
rect -44 1872 0 1924
rect 156 1872 200 1924
rect -44 1800 200 1872
rect -44 1748 0 1800
rect 156 1748 200 1800
rect -44 1676 200 1748
rect -44 1624 0 1676
rect 156 1624 200 1676
rect -44 1552 200 1624
rect -44 1500 0 1552
rect 156 1500 200 1552
rect -44 1428 200 1500
rect -44 1376 0 1428
rect 156 1376 200 1428
rect -44 1304 200 1376
rect -44 1252 0 1304
rect 156 1252 200 1304
rect -44 1180 200 1252
rect -44 1128 0 1180
rect 156 1128 200 1180
rect -44 1056 200 1128
rect -44 1004 0 1056
rect 156 1004 200 1056
rect -44 932 200 1004
rect -44 880 0 932
rect 156 880 200 932
rect -44 808 200 880
rect -44 756 0 808
rect 156 756 200 808
rect -44 684 200 756
rect -44 632 0 684
rect 156 632 200 684
rect -44 560 200 632
rect -44 508 0 560
rect 156 508 200 560
rect -44 436 200 508
rect -44 384 0 436
rect 156 384 200 436
rect -44 312 200 384
rect -44 260 0 312
rect 156 260 200 312
rect -44 188 200 260
rect -44 136 0 188
rect 156 136 200 188
rect -44 64 200 136
rect -44 12 0 64
rect 156 12 200 64
rect -44 0 200 12
rect 340 11968 1584 12000
rect 340 11916 378 11968
rect 430 11916 502 11968
rect 554 11916 626 11968
rect 678 11916 750 11968
rect 802 11916 874 11968
rect 926 11916 998 11968
rect 1050 11916 1122 11968
rect 1174 11916 1246 11968
rect 1298 11916 1370 11968
rect 1422 11916 1494 11968
rect 1546 11916 1584 11968
rect 340 11844 1584 11916
rect 340 11792 378 11844
rect 430 11792 502 11844
rect 554 11792 626 11844
rect 678 11792 750 11844
rect 802 11792 874 11844
rect 926 11792 998 11844
rect 1050 11792 1122 11844
rect 1174 11792 1246 11844
rect 1298 11792 1370 11844
rect 1422 11792 1494 11844
rect 1546 11792 1584 11844
rect 340 11720 1584 11792
rect 340 11668 378 11720
rect 430 11668 502 11720
rect 554 11668 626 11720
rect 678 11668 750 11720
rect 802 11668 874 11720
rect 926 11668 998 11720
rect 1050 11668 1122 11720
rect 1174 11668 1246 11720
rect 1298 11668 1370 11720
rect 1422 11668 1494 11720
rect 1546 11668 1584 11720
rect 340 11596 1584 11668
rect 340 11544 378 11596
rect 430 11544 502 11596
rect 554 11544 626 11596
rect 678 11544 750 11596
rect 802 11544 874 11596
rect 926 11544 998 11596
rect 1050 11544 1122 11596
rect 1174 11544 1246 11596
rect 1298 11544 1370 11596
rect 1422 11544 1494 11596
rect 1546 11544 1584 11596
rect 340 11472 1584 11544
rect 340 11420 378 11472
rect 430 11420 502 11472
rect 554 11420 626 11472
rect 678 11420 750 11472
rect 802 11420 874 11472
rect 926 11420 998 11472
rect 1050 11420 1122 11472
rect 1174 11420 1246 11472
rect 1298 11420 1370 11472
rect 1422 11420 1494 11472
rect 1546 11420 1584 11472
rect 340 11348 1584 11420
rect 340 11296 378 11348
rect 430 11296 502 11348
rect 554 11296 626 11348
rect 678 11296 750 11348
rect 802 11296 874 11348
rect 926 11296 998 11348
rect 1050 11296 1122 11348
rect 1174 11296 1246 11348
rect 1298 11296 1370 11348
rect 1422 11296 1494 11348
rect 1546 11296 1584 11348
rect 340 11224 1584 11296
rect 340 11172 378 11224
rect 430 11172 502 11224
rect 554 11172 626 11224
rect 678 11172 750 11224
rect 802 11172 874 11224
rect 926 11172 998 11224
rect 1050 11172 1122 11224
rect 1174 11172 1246 11224
rect 1298 11172 1370 11224
rect 1422 11172 1494 11224
rect 1546 11172 1584 11224
rect 340 11100 1584 11172
rect 340 11048 378 11100
rect 430 11048 502 11100
rect 554 11048 626 11100
rect 678 11048 750 11100
rect 802 11048 874 11100
rect 926 11048 998 11100
rect 1050 11048 1122 11100
rect 1174 11048 1246 11100
rect 1298 11048 1370 11100
rect 1422 11048 1494 11100
rect 1546 11048 1584 11100
rect 340 10976 1584 11048
rect 340 10924 378 10976
rect 430 10924 502 10976
rect 554 10924 626 10976
rect 678 10924 750 10976
rect 802 10924 874 10976
rect 926 10924 998 10976
rect 1050 10924 1122 10976
rect 1174 10924 1246 10976
rect 1298 10924 1370 10976
rect 1422 10924 1494 10976
rect 1546 10924 1584 10976
rect 340 10852 1584 10924
rect 340 10800 378 10852
rect 430 10800 502 10852
rect 554 10800 626 10852
rect 678 10800 750 10852
rect 802 10800 874 10852
rect 926 10800 998 10852
rect 1050 10800 1122 10852
rect 1174 10800 1246 10852
rect 1298 10800 1370 10852
rect 1422 10800 1494 10852
rect 1546 10800 1584 10852
rect 340 10728 1584 10800
rect 340 10676 378 10728
rect 430 10676 502 10728
rect 554 10676 626 10728
rect 678 10676 750 10728
rect 802 10676 874 10728
rect 926 10676 998 10728
rect 1050 10676 1122 10728
rect 1174 10676 1246 10728
rect 1298 10676 1370 10728
rect 1422 10676 1494 10728
rect 1546 10676 1584 10728
rect 340 10604 1584 10676
rect 340 10552 378 10604
rect 430 10552 502 10604
rect 554 10552 626 10604
rect 678 10552 750 10604
rect 802 10552 874 10604
rect 926 10552 998 10604
rect 1050 10552 1122 10604
rect 1174 10552 1246 10604
rect 1298 10552 1370 10604
rect 1422 10552 1494 10604
rect 1546 10552 1584 10604
rect 340 10480 1584 10552
rect 340 10428 378 10480
rect 430 10428 502 10480
rect 554 10428 626 10480
rect 678 10428 750 10480
rect 802 10428 874 10480
rect 926 10428 998 10480
rect 1050 10428 1122 10480
rect 1174 10428 1246 10480
rect 1298 10428 1370 10480
rect 1422 10428 1494 10480
rect 1546 10428 1584 10480
rect 340 10356 1584 10428
rect 340 10304 378 10356
rect 430 10304 502 10356
rect 554 10304 626 10356
rect 678 10304 750 10356
rect 802 10304 874 10356
rect 926 10304 998 10356
rect 1050 10304 1122 10356
rect 1174 10304 1246 10356
rect 1298 10304 1370 10356
rect 1422 10304 1494 10356
rect 1546 10304 1584 10356
rect 340 10232 1584 10304
rect 340 10180 378 10232
rect 430 10180 502 10232
rect 554 10180 626 10232
rect 678 10180 750 10232
rect 802 10180 874 10232
rect 926 10180 998 10232
rect 1050 10180 1122 10232
rect 1174 10180 1246 10232
rect 1298 10180 1370 10232
rect 1422 10180 1494 10232
rect 1546 10180 1584 10232
rect 340 10108 1584 10180
rect 340 10056 378 10108
rect 430 10056 502 10108
rect 554 10056 626 10108
rect 678 10056 750 10108
rect 802 10056 874 10108
rect 926 10056 998 10108
rect 1050 10056 1122 10108
rect 1174 10056 1246 10108
rect 1298 10056 1370 10108
rect 1422 10056 1494 10108
rect 1546 10056 1584 10108
rect 340 9984 1584 10056
rect 340 9932 378 9984
rect 430 9932 502 9984
rect 554 9932 626 9984
rect 678 9932 750 9984
rect 802 9932 874 9984
rect 926 9932 998 9984
rect 1050 9932 1122 9984
rect 1174 9932 1246 9984
rect 1298 9932 1370 9984
rect 1422 9932 1494 9984
rect 1546 9932 1584 9984
rect 340 9860 1584 9932
rect 340 9808 378 9860
rect 430 9808 502 9860
rect 554 9808 626 9860
rect 678 9808 750 9860
rect 802 9808 874 9860
rect 926 9808 998 9860
rect 1050 9808 1122 9860
rect 1174 9808 1246 9860
rect 1298 9808 1370 9860
rect 1422 9808 1494 9860
rect 1546 9808 1584 9860
rect 340 9736 1584 9808
rect 340 9684 378 9736
rect 430 9684 502 9736
rect 554 9684 626 9736
rect 678 9684 750 9736
rect 802 9684 874 9736
rect 926 9684 998 9736
rect 1050 9684 1122 9736
rect 1174 9684 1246 9736
rect 1298 9684 1370 9736
rect 1422 9684 1494 9736
rect 1546 9684 1584 9736
rect 340 9612 1584 9684
rect 340 9560 378 9612
rect 430 9560 502 9612
rect 554 9560 626 9612
rect 678 9560 750 9612
rect 802 9560 874 9612
rect 926 9560 998 9612
rect 1050 9560 1122 9612
rect 1174 9560 1246 9612
rect 1298 9560 1370 9612
rect 1422 9560 1494 9612
rect 1546 9560 1584 9612
rect 340 9488 1584 9560
rect 340 9436 378 9488
rect 430 9436 502 9488
rect 554 9436 626 9488
rect 678 9436 750 9488
rect 802 9436 874 9488
rect 926 9436 998 9488
rect 1050 9436 1122 9488
rect 1174 9436 1246 9488
rect 1298 9436 1370 9488
rect 1422 9436 1494 9488
rect 1546 9436 1584 9488
rect 340 9364 1584 9436
rect 340 9312 378 9364
rect 430 9312 502 9364
rect 554 9312 626 9364
rect 678 9312 750 9364
rect 802 9312 874 9364
rect 926 9312 998 9364
rect 1050 9312 1122 9364
rect 1174 9312 1246 9364
rect 1298 9312 1370 9364
rect 1422 9312 1494 9364
rect 1546 9312 1584 9364
rect 340 9240 1584 9312
rect 340 9188 378 9240
rect 430 9188 502 9240
rect 554 9188 626 9240
rect 678 9188 750 9240
rect 802 9188 874 9240
rect 926 9188 998 9240
rect 1050 9188 1122 9240
rect 1174 9188 1246 9240
rect 1298 9188 1370 9240
rect 1422 9188 1494 9240
rect 1546 9188 1584 9240
rect 340 9116 1584 9188
rect 340 9064 378 9116
rect 430 9064 502 9116
rect 554 9064 626 9116
rect 678 9064 750 9116
rect 802 9064 874 9116
rect 926 9064 998 9116
rect 1050 9064 1122 9116
rect 1174 9064 1246 9116
rect 1298 9064 1370 9116
rect 1422 9064 1494 9116
rect 1546 9064 1584 9116
rect 340 8992 1584 9064
rect 340 8940 378 8992
rect 430 8940 502 8992
rect 554 8940 626 8992
rect 678 8940 750 8992
rect 802 8940 874 8992
rect 926 8940 998 8992
rect 1050 8940 1122 8992
rect 1174 8940 1246 8992
rect 1298 8940 1370 8992
rect 1422 8940 1494 8992
rect 1546 8940 1584 8992
rect 340 8868 1584 8940
rect 340 8816 378 8868
rect 430 8816 502 8868
rect 554 8816 626 8868
rect 678 8816 750 8868
rect 802 8816 874 8868
rect 926 8816 998 8868
rect 1050 8816 1122 8868
rect 1174 8816 1246 8868
rect 1298 8816 1370 8868
rect 1422 8816 1494 8868
rect 1546 8816 1584 8868
rect 340 8744 1584 8816
rect 340 8692 378 8744
rect 430 8692 502 8744
rect 554 8692 626 8744
rect 678 8692 750 8744
rect 802 8692 874 8744
rect 926 8692 998 8744
rect 1050 8692 1122 8744
rect 1174 8692 1246 8744
rect 1298 8692 1370 8744
rect 1422 8692 1494 8744
rect 1546 8692 1584 8744
rect 340 8620 1584 8692
rect 340 8568 378 8620
rect 430 8568 502 8620
rect 554 8568 626 8620
rect 678 8568 750 8620
rect 802 8568 874 8620
rect 926 8568 998 8620
rect 1050 8568 1122 8620
rect 1174 8568 1246 8620
rect 1298 8568 1370 8620
rect 1422 8568 1494 8620
rect 1546 8568 1584 8620
rect 340 8496 1584 8568
rect 340 8444 378 8496
rect 430 8444 502 8496
rect 554 8444 626 8496
rect 678 8444 750 8496
rect 802 8444 874 8496
rect 926 8444 998 8496
rect 1050 8444 1122 8496
rect 1174 8444 1246 8496
rect 1298 8444 1370 8496
rect 1422 8444 1494 8496
rect 1546 8444 1584 8496
rect 340 8372 1584 8444
rect 340 8320 378 8372
rect 430 8320 502 8372
rect 554 8320 626 8372
rect 678 8320 750 8372
rect 802 8320 874 8372
rect 926 8320 998 8372
rect 1050 8320 1122 8372
rect 1174 8320 1246 8372
rect 1298 8320 1370 8372
rect 1422 8320 1494 8372
rect 1546 8320 1584 8372
rect 340 8248 1584 8320
rect 340 8196 378 8248
rect 430 8196 502 8248
rect 554 8196 626 8248
rect 678 8196 750 8248
rect 802 8196 874 8248
rect 926 8196 998 8248
rect 1050 8196 1122 8248
rect 1174 8196 1246 8248
rect 1298 8196 1370 8248
rect 1422 8196 1494 8248
rect 1546 8196 1584 8248
rect 340 8124 1584 8196
rect 340 8072 378 8124
rect 430 8072 502 8124
rect 554 8072 626 8124
rect 678 8072 750 8124
rect 802 8072 874 8124
rect 926 8072 998 8124
rect 1050 8072 1122 8124
rect 1174 8072 1246 8124
rect 1298 8072 1370 8124
rect 1422 8072 1494 8124
rect 1546 8072 1584 8124
rect 340 8000 1584 8072
rect 340 7948 378 8000
rect 430 7948 502 8000
rect 554 7948 626 8000
rect 678 7948 750 8000
rect 802 7948 874 8000
rect 926 7948 998 8000
rect 1050 7948 1122 8000
rect 1174 7948 1246 8000
rect 1298 7948 1370 8000
rect 1422 7948 1494 8000
rect 1546 7948 1584 8000
rect 340 7876 1584 7948
rect 340 7824 378 7876
rect 430 7824 502 7876
rect 554 7824 626 7876
rect 678 7824 750 7876
rect 802 7824 874 7876
rect 926 7824 998 7876
rect 1050 7824 1122 7876
rect 1174 7824 1246 7876
rect 1298 7824 1370 7876
rect 1422 7824 1494 7876
rect 1546 7824 1584 7876
rect 340 7752 1584 7824
rect 340 7700 378 7752
rect 430 7700 502 7752
rect 554 7700 626 7752
rect 678 7700 750 7752
rect 802 7700 874 7752
rect 926 7700 998 7752
rect 1050 7700 1122 7752
rect 1174 7700 1246 7752
rect 1298 7700 1370 7752
rect 1422 7700 1494 7752
rect 1546 7700 1584 7752
rect 340 7628 1584 7700
rect 340 7576 378 7628
rect 430 7576 502 7628
rect 554 7576 626 7628
rect 678 7576 750 7628
rect 802 7576 874 7628
rect 926 7576 998 7628
rect 1050 7576 1122 7628
rect 1174 7576 1246 7628
rect 1298 7576 1370 7628
rect 1422 7576 1494 7628
rect 1546 7576 1584 7628
rect 340 7504 1584 7576
rect 340 7452 378 7504
rect 430 7452 502 7504
rect 554 7452 626 7504
rect 678 7452 750 7504
rect 802 7452 874 7504
rect 926 7452 998 7504
rect 1050 7452 1122 7504
rect 1174 7452 1246 7504
rect 1298 7452 1370 7504
rect 1422 7452 1494 7504
rect 1546 7452 1584 7504
rect 340 7380 1584 7452
rect 340 7328 378 7380
rect 430 7328 502 7380
rect 554 7328 626 7380
rect 678 7328 750 7380
rect 802 7328 874 7380
rect 926 7328 998 7380
rect 1050 7328 1122 7380
rect 1174 7328 1246 7380
rect 1298 7328 1370 7380
rect 1422 7328 1494 7380
rect 1546 7328 1584 7380
rect 340 7256 1584 7328
rect 340 7204 378 7256
rect 430 7204 502 7256
rect 554 7204 626 7256
rect 678 7204 750 7256
rect 802 7204 874 7256
rect 926 7204 998 7256
rect 1050 7204 1122 7256
rect 1174 7204 1246 7256
rect 1298 7204 1370 7256
rect 1422 7204 1494 7256
rect 1546 7204 1584 7256
rect 340 7132 1584 7204
rect 340 7080 378 7132
rect 430 7080 502 7132
rect 554 7080 626 7132
rect 678 7080 750 7132
rect 802 7080 874 7132
rect 926 7080 998 7132
rect 1050 7080 1122 7132
rect 1174 7080 1246 7132
rect 1298 7080 1370 7132
rect 1422 7080 1494 7132
rect 1546 7080 1584 7132
rect 340 7008 1584 7080
rect 340 6956 378 7008
rect 430 6956 502 7008
rect 554 6956 626 7008
rect 678 6956 750 7008
rect 802 6956 874 7008
rect 926 6956 998 7008
rect 1050 6956 1122 7008
rect 1174 6956 1246 7008
rect 1298 6956 1370 7008
rect 1422 6956 1494 7008
rect 1546 6956 1584 7008
rect 340 6884 1584 6956
rect 340 6832 378 6884
rect 430 6832 502 6884
rect 554 6832 626 6884
rect 678 6832 750 6884
rect 802 6832 874 6884
rect 926 6832 998 6884
rect 1050 6832 1122 6884
rect 1174 6832 1246 6884
rect 1298 6832 1370 6884
rect 1422 6832 1494 6884
rect 1546 6832 1584 6884
rect 340 6760 1584 6832
rect 340 6708 378 6760
rect 430 6708 502 6760
rect 554 6708 626 6760
rect 678 6708 750 6760
rect 802 6708 874 6760
rect 926 6708 998 6760
rect 1050 6708 1122 6760
rect 1174 6708 1246 6760
rect 1298 6708 1370 6760
rect 1422 6708 1494 6760
rect 1546 6708 1584 6760
rect 340 6636 1584 6708
rect 340 6584 378 6636
rect 430 6584 502 6636
rect 554 6584 626 6636
rect 678 6584 750 6636
rect 802 6584 874 6636
rect 926 6584 998 6636
rect 1050 6584 1122 6636
rect 1174 6584 1246 6636
rect 1298 6584 1370 6636
rect 1422 6584 1494 6636
rect 1546 6584 1584 6636
rect 340 6512 1584 6584
rect 340 6460 378 6512
rect 430 6460 502 6512
rect 554 6460 626 6512
rect 678 6460 750 6512
rect 802 6460 874 6512
rect 926 6460 998 6512
rect 1050 6460 1122 6512
rect 1174 6460 1246 6512
rect 1298 6460 1370 6512
rect 1422 6460 1494 6512
rect 1546 6460 1584 6512
rect 340 6388 1584 6460
rect 340 6336 378 6388
rect 430 6336 502 6388
rect 554 6336 626 6388
rect 678 6336 750 6388
rect 802 6336 874 6388
rect 926 6336 998 6388
rect 1050 6336 1122 6388
rect 1174 6336 1246 6388
rect 1298 6336 1370 6388
rect 1422 6336 1494 6388
rect 1546 6336 1584 6388
rect 340 6264 1584 6336
rect 340 6212 378 6264
rect 430 6212 502 6264
rect 554 6212 626 6264
rect 678 6212 750 6264
rect 802 6212 874 6264
rect 926 6212 998 6264
rect 1050 6212 1122 6264
rect 1174 6212 1246 6264
rect 1298 6212 1370 6264
rect 1422 6212 1494 6264
rect 1546 6212 1584 6264
rect 340 6140 1584 6212
rect 340 6088 378 6140
rect 430 6088 502 6140
rect 554 6088 626 6140
rect 678 6088 750 6140
rect 802 6088 874 6140
rect 926 6088 998 6140
rect 1050 6088 1122 6140
rect 1174 6088 1246 6140
rect 1298 6088 1370 6140
rect 1422 6088 1494 6140
rect 1546 6088 1584 6140
rect 340 6016 1584 6088
rect 340 5964 378 6016
rect 430 5964 502 6016
rect 554 5964 626 6016
rect 678 5964 750 6016
rect 802 5964 874 6016
rect 926 5964 998 6016
rect 1050 5964 1122 6016
rect 1174 5964 1246 6016
rect 1298 5964 1370 6016
rect 1422 5964 1494 6016
rect 1546 5964 1584 6016
rect 340 5892 1584 5964
rect 340 5840 378 5892
rect 430 5840 502 5892
rect 554 5840 626 5892
rect 678 5840 750 5892
rect 802 5840 874 5892
rect 926 5840 998 5892
rect 1050 5840 1122 5892
rect 1174 5840 1246 5892
rect 1298 5840 1370 5892
rect 1422 5840 1494 5892
rect 1546 5840 1584 5892
rect 340 5768 1584 5840
rect 340 5716 378 5768
rect 430 5716 502 5768
rect 554 5716 626 5768
rect 678 5716 750 5768
rect 802 5716 874 5768
rect 926 5716 998 5768
rect 1050 5716 1122 5768
rect 1174 5716 1246 5768
rect 1298 5716 1370 5768
rect 1422 5716 1494 5768
rect 1546 5716 1584 5768
rect 340 5644 1584 5716
rect 340 5592 378 5644
rect 430 5592 502 5644
rect 554 5592 626 5644
rect 678 5592 750 5644
rect 802 5592 874 5644
rect 926 5592 998 5644
rect 1050 5592 1122 5644
rect 1174 5592 1246 5644
rect 1298 5592 1370 5644
rect 1422 5592 1494 5644
rect 1546 5592 1584 5644
rect 340 5520 1584 5592
rect 340 5468 378 5520
rect 430 5468 502 5520
rect 554 5468 626 5520
rect 678 5468 750 5520
rect 802 5468 874 5520
rect 926 5468 998 5520
rect 1050 5468 1122 5520
rect 1174 5468 1246 5520
rect 1298 5468 1370 5520
rect 1422 5468 1494 5520
rect 1546 5468 1584 5520
rect 340 5396 1584 5468
rect 340 5344 378 5396
rect 430 5344 502 5396
rect 554 5344 626 5396
rect 678 5344 750 5396
rect 802 5344 874 5396
rect 926 5344 998 5396
rect 1050 5344 1122 5396
rect 1174 5344 1246 5396
rect 1298 5344 1370 5396
rect 1422 5344 1494 5396
rect 1546 5344 1584 5396
rect 340 5272 1584 5344
rect 340 5220 378 5272
rect 430 5220 502 5272
rect 554 5220 626 5272
rect 678 5220 750 5272
rect 802 5220 874 5272
rect 926 5220 998 5272
rect 1050 5220 1122 5272
rect 1174 5220 1246 5272
rect 1298 5220 1370 5272
rect 1422 5220 1494 5272
rect 1546 5220 1584 5272
rect 340 5148 1584 5220
rect 340 5096 378 5148
rect 430 5096 502 5148
rect 554 5096 626 5148
rect 678 5096 750 5148
rect 802 5096 874 5148
rect 926 5096 998 5148
rect 1050 5096 1122 5148
rect 1174 5096 1246 5148
rect 1298 5096 1370 5148
rect 1422 5096 1494 5148
rect 1546 5096 1584 5148
rect 340 5024 1584 5096
rect 340 4972 378 5024
rect 430 4972 502 5024
rect 554 4972 626 5024
rect 678 4972 750 5024
rect 802 4972 874 5024
rect 926 4972 998 5024
rect 1050 4972 1122 5024
rect 1174 4972 1246 5024
rect 1298 4972 1370 5024
rect 1422 4972 1494 5024
rect 1546 4972 1584 5024
rect 340 4900 1584 4972
rect 340 4848 378 4900
rect 430 4848 502 4900
rect 554 4848 626 4900
rect 678 4848 750 4900
rect 802 4848 874 4900
rect 926 4848 998 4900
rect 1050 4848 1122 4900
rect 1174 4848 1246 4900
rect 1298 4848 1370 4900
rect 1422 4848 1494 4900
rect 1546 4848 1584 4900
rect 340 4776 1584 4848
rect 340 4724 378 4776
rect 430 4724 502 4776
rect 554 4724 626 4776
rect 678 4724 750 4776
rect 802 4724 874 4776
rect 926 4724 998 4776
rect 1050 4724 1122 4776
rect 1174 4724 1246 4776
rect 1298 4724 1370 4776
rect 1422 4724 1494 4776
rect 1546 4724 1584 4776
rect 340 4652 1584 4724
rect 340 4600 378 4652
rect 430 4600 502 4652
rect 554 4600 626 4652
rect 678 4600 750 4652
rect 802 4600 874 4652
rect 926 4600 998 4652
rect 1050 4600 1122 4652
rect 1174 4600 1246 4652
rect 1298 4600 1370 4652
rect 1422 4600 1494 4652
rect 1546 4600 1584 4652
rect 340 4528 1584 4600
rect 340 4476 378 4528
rect 430 4476 502 4528
rect 554 4476 626 4528
rect 678 4476 750 4528
rect 802 4476 874 4528
rect 926 4476 998 4528
rect 1050 4476 1122 4528
rect 1174 4476 1246 4528
rect 1298 4476 1370 4528
rect 1422 4476 1494 4528
rect 1546 4476 1584 4528
rect 340 4404 1584 4476
rect 340 4352 378 4404
rect 430 4352 502 4404
rect 554 4352 626 4404
rect 678 4352 750 4404
rect 802 4352 874 4404
rect 926 4352 998 4404
rect 1050 4352 1122 4404
rect 1174 4352 1246 4404
rect 1298 4352 1370 4404
rect 1422 4352 1494 4404
rect 1546 4352 1584 4404
rect 340 4280 1584 4352
rect 340 4228 378 4280
rect 430 4228 502 4280
rect 554 4228 626 4280
rect 678 4228 750 4280
rect 802 4228 874 4280
rect 926 4228 998 4280
rect 1050 4228 1122 4280
rect 1174 4228 1246 4280
rect 1298 4228 1370 4280
rect 1422 4228 1494 4280
rect 1546 4228 1584 4280
rect 340 4156 1584 4228
rect 340 4104 378 4156
rect 430 4104 502 4156
rect 554 4104 626 4156
rect 678 4104 750 4156
rect 802 4104 874 4156
rect 926 4104 998 4156
rect 1050 4104 1122 4156
rect 1174 4104 1246 4156
rect 1298 4104 1370 4156
rect 1422 4104 1494 4156
rect 1546 4104 1584 4156
rect 340 4032 1584 4104
rect 340 3980 378 4032
rect 430 3980 502 4032
rect 554 3980 626 4032
rect 678 3980 750 4032
rect 802 3980 874 4032
rect 926 3980 998 4032
rect 1050 3980 1122 4032
rect 1174 3980 1246 4032
rect 1298 3980 1370 4032
rect 1422 3980 1494 4032
rect 1546 3980 1584 4032
rect 340 3908 1584 3980
rect 340 3856 378 3908
rect 430 3856 502 3908
rect 554 3856 626 3908
rect 678 3856 750 3908
rect 802 3856 874 3908
rect 926 3856 998 3908
rect 1050 3856 1122 3908
rect 1174 3856 1246 3908
rect 1298 3856 1370 3908
rect 1422 3856 1494 3908
rect 1546 3856 1584 3908
rect 340 3784 1584 3856
rect 340 3732 378 3784
rect 430 3732 502 3784
rect 554 3732 626 3784
rect 678 3732 750 3784
rect 802 3732 874 3784
rect 926 3732 998 3784
rect 1050 3732 1122 3784
rect 1174 3732 1246 3784
rect 1298 3732 1370 3784
rect 1422 3732 1494 3784
rect 1546 3732 1584 3784
rect 340 3660 1584 3732
rect 340 3608 378 3660
rect 430 3608 502 3660
rect 554 3608 626 3660
rect 678 3608 750 3660
rect 802 3608 874 3660
rect 926 3608 998 3660
rect 1050 3608 1122 3660
rect 1174 3608 1246 3660
rect 1298 3608 1370 3660
rect 1422 3608 1494 3660
rect 1546 3608 1584 3660
rect 340 3536 1584 3608
rect 340 3484 378 3536
rect 430 3484 502 3536
rect 554 3484 626 3536
rect 678 3484 750 3536
rect 802 3484 874 3536
rect 926 3484 998 3536
rect 1050 3484 1122 3536
rect 1174 3484 1246 3536
rect 1298 3484 1370 3536
rect 1422 3484 1494 3536
rect 1546 3484 1584 3536
rect 340 3412 1584 3484
rect 340 3360 378 3412
rect 430 3360 502 3412
rect 554 3360 626 3412
rect 678 3360 750 3412
rect 802 3360 874 3412
rect 926 3360 998 3412
rect 1050 3360 1122 3412
rect 1174 3360 1246 3412
rect 1298 3360 1370 3412
rect 1422 3360 1494 3412
rect 1546 3360 1584 3412
rect 340 3288 1584 3360
rect 340 3236 378 3288
rect 430 3236 502 3288
rect 554 3236 626 3288
rect 678 3236 750 3288
rect 802 3236 874 3288
rect 926 3236 998 3288
rect 1050 3236 1122 3288
rect 1174 3236 1246 3288
rect 1298 3236 1370 3288
rect 1422 3236 1494 3288
rect 1546 3236 1584 3288
rect 340 3164 1584 3236
rect 340 3112 378 3164
rect 430 3112 502 3164
rect 554 3112 626 3164
rect 678 3112 750 3164
rect 802 3112 874 3164
rect 926 3112 998 3164
rect 1050 3112 1122 3164
rect 1174 3112 1246 3164
rect 1298 3112 1370 3164
rect 1422 3112 1494 3164
rect 1546 3112 1584 3164
rect 340 3040 1584 3112
rect 340 2988 378 3040
rect 430 2988 502 3040
rect 554 2988 626 3040
rect 678 2988 750 3040
rect 802 2988 874 3040
rect 926 2988 998 3040
rect 1050 2988 1122 3040
rect 1174 2988 1246 3040
rect 1298 2988 1370 3040
rect 1422 2988 1494 3040
rect 1546 2988 1584 3040
rect 340 2916 1584 2988
rect 340 2864 378 2916
rect 430 2864 502 2916
rect 554 2864 626 2916
rect 678 2864 750 2916
rect 802 2864 874 2916
rect 926 2864 998 2916
rect 1050 2864 1122 2916
rect 1174 2864 1246 2916
rect 1298 2864 1370 2916
rect 1422 2864 1494 2916
rect 1546 2864 1584 2916
rect 340 2792 1584 2864
rect 340 2740 378 2792
rect 430 2740 502 2792
rect 554 2740 626 2792
rect 678 2740 750 2792
rect 802 2740 874 2792
rect 926 2740 998 2792
rect 1050 2740 1122 2792
rect 1174 2740 1246 2792
rect 1298 2740 1370 2792
rect 1422 2740 1494 2792
rect 1546 2740 1584 2792
rect 340 2668 1584 2740
rect 340 2616 378 2668
rect 430 2616 502 2668
rect 554 2616 626 2668
rect 678 2616 750 2668
rect 802 2616 874 2668
rect 926 2616 998 2668
rect 1050 2616 1122 2668
rect 1174 2616 1246 2668
rect 1298 2616 1370 2668
rect 1422 2616 1494 2668
rect 1546 2616 1584 2668
rect 340 2544 1584 2616
rect 340 2492 378 2544
rect 430 2492 502 2544
rect 554 2492 626 2544
rect 678 2492 750 2544
rect 802 2492 874 2544
rect 926 2492 998 2544
rect 1050 2492 1122 2544
rect 1174 2492 1246 2544
rect 1298 2492 1370 2544
rect 1422 2492 1494 2544
rect 1546 2492 1584 2544
rect 340 2420 1584 2492
rect 340 2368 378 2420
rect 430 2368 502 2420
rect 554 2368 626 2420
rect 678 2368 750 2420
rect 802 2368 874 2420
rect 926 2368 998 2420
rect 1050 2368 1122 2420
rect 1174 2368 1246 2420
rect 1298 2368 1370 2420
rect 1422 2368 1494 2420
rect 1546 2368 1584 2420
rect 340 2296 1584 2368
rect 340 2244 378 2296
rect 430 2244 502 2296
rect 554 2244 626 2296
rect 678 2244 750 2296
rect 802 2244 874 2296
rect 926 2244 998 2296
rect 1050 2244 1122 2296
rect 1174 2244 1246 2296
rect 1298 2244 1370 2296
rect 1422 2244 1494 2296
rect 1546 2244 1584 2296
rect 340 2172 1584 2244
rect 340 2120 378 2172
rect 430 2120 502 2172
rect 554 2120 626 2172
rect 678 2120 750 2172
rect 802 2120 874 2172
rect 926 2120 998 2172
rect 1050 2120 1122 2172
rect 1174 2120 1246 2172
rect 1298 2120 1370 2172
rect 1422 2120 1494 2172
rect 1546 2120 1584 2172
rect 340 2048 1584 2120
rect 340 1996 378 2048
rect 430 1996 502 2048
rect 554 1996 626 2048
rect 678 1996 750 2048
rect 802 1996 874 2048
rect 926 1996 998 2048
rect 1050 1996 1122 2048
rect 1174 1996 1246 2048
rect 1298 1996 1370 2048
rect 1422 1996 1494 2048
rect 1546 1996 1584 2048
rect 340 1924 1584 1996
rect 340 1872 378 1924
rect 430 1872 502 1924
rect 554 1872 626 1924
rect 678 1872 750 1924
rect 802 1872 874 1924
rect 926 1872 998 1924
rect 1050 1872 1122 1924
rect 1174 1872 1246 1924
rect 1298 1872 1370 1924
rect 1422 1872 1494 1924
rect 1546 1872 1584 1924
rect 340 1800 1584 1872
rect 340 1748 378 1800
rect 430 1748 502 1800
rect 554 1748 626 1800
rect 678 1748 750 1800
rect 802 1748 874 1800
rect 926 1748 998 1800
rect 1050 1748 1122 1800
rect 1174 1748 1246 1800
rect 1298 1748 1370 1800
rect 1422 1748 1494 1800
rect 1546 1748 1584 1800
rect 340 1676 1584 1748
rect 340 1624 378 1676
rect 430 1624 502 1676
rect 554 1624 626 1676
rect 678 1624 750 1676
rect 802 1624 874 1676
rect 926 1624 998 1676
rect 1050 1624 1122 1676
rect 1174 1624 1246 1676
rect 1298 1624 1370 1676
rect 1422 1624 1494 1676
rect 1546 1624 1584 1676
rect 340 1552 1584 1624
rect 340 1500 378 1552
rect 430 1500 502 1552
rect 554 1500 626 1552
rect 678 1500 750 1552
rect 802 1500 874 1552
rect 926 1500 998 1552
rect 1050 1500 1122 1552
rect 1174 1500 1246 1552
rect 1298 1500 1370 1552
rect 1422 1500 1494 1552
rect 1546 1500 1584 1552
rect 340 1428 1584 1500
rect 340 1376 378 1428
rect 430 1376 502 1428
rect 554 1376 626 1428
rect 678 1376 750 1428
rect 802 1376 874 1428
rect 926 1376 998 1428
rect 1050 1376 1122 1428
rect 1174 1376 1246 1428
rect 1298 1376 1370 1428
rect 1422 1376 1494 1428
rect 1546 1376 1584 1428
rect 340 1304 1584 1376
rect 340 1252 378 1304
rect 430 1252 502 1304
rect 554 1252 626 1304
rect 678 1252 750 1304
rect 802 1252 874 1304
rect 926 1252 998 1304
rect 1050 1252 1122 1304
rect 1174 1252 1246 1304
rect 1298 1252 1370 1304
rect 1422 1252 1494 1304
rect 1546 1252 1584 1304
rect 340 1180 1584 1252
rect 340 1128 378 1180
rect 430 1128 502 1180
rect 554 1128 626 1180
rect 678 1128 750 1180
rect 802 1128 874 1180
rect 926 1128 998 1180
rect 1050 1128 1122 1180
rect 1174 1128 1246 1180
rect 1298 1128 1370 1180
rect 1422 1128 1494 1180
rect 1546 1128 1584 1180
rect 340 1056 1584 1128
rect 340 1004 378 1056
rect 430 1004 502 1056
rect 554 1004 626 1056
rect 678 1004 750 1056
rect 802 1004 874 1056
rect 926 1004 998 1056
rect 1050 1004 1122 1056
rect 1174 1004 1246 1056
rect 1298 1004 1370 1056
rect 1422 1004 1494 1056
rect 1546 1004 1584 1056
rect 340 932 1584 1004
rect 340 880 378 932
rect 430 880 502 932
rect 554 880 626 932
rect 678 880 750 932
rect 802 880 874 932
rect 926 880 998 932
rect 1050 880 1122 932
rect 1174 880 1246 932
rect 1298 880 1370 932
rect 1422 880 1494 932
rect 1546 880 1584 932
rect 340 808 1584 880
rect 340 756 378 808
rect 430 756 502 808
rect 554 756 626 808
rect 678 756 750 808
rect 802 756 874 808
rect 926 756 998 808
rect 1050 756 1122 808
rect 1174 756 1246 808
rect 1298 756 1370 808
rect 1422 756 1494 808
rect 1546 756 1584 808
rect 340 684 1584 756
rect 340 632 378 684
rect 430 632 502 684
rect 554 632 626 684
rect 678 632 750 684
rect 802 632 874 684
rect 926 632 998 684
rect 1050 632 1122 684
rect 1174 632 1246 684
rect 1298 632 1370 684
rect 1422 632 1494 684
rect 1546 632 1584 684
rect 340 560 1584 632
rect 340 508 378 560
rect 430 508 502 560
rect 554 508 626 560
rect 678 508 750 560
rect 802 508 874 560
rect 926 508 998 560
rect 1050 508 1122 560
rect 1174 508 1246 560
rect 1298 508 1370 560
rect 1422 508 1494 560
rect 1546 508 1584 560
rect 340 436 1584 508
rect 340 384 378 436
rect 430 384 502 436
rect 554 384 626 436
rect 678 384 750 436
rect 802 384 874 436
rect 926 384 998 436
rect 1050 384 1122 436
rect 1174 384 1246 436
rect 1298 384 1370 436
rect 1422 384 1494 436
rect 1546 384 1584 436
rect 340 312 1584 384
rect 340 260 378 312
rect 430 260 502 312
rect 554 260 626 312
rect 678 260 750 312
rect 802 260 874 312
rect 926 260 998 312
rect 1050 260 1122 312
rect 1174 260 1246 312
rect 1298 260 1370 312
rect 1422 260 1494 312
rect 1546 260 1584 312
rect 340 188 1584 260
rect 340 136 378 188
rect 430 136 502 188
rect 554 136 626 188
rect 678 136 750 188
rect 802 136 874 188
rect 926 136 998 188
rect 1050 136 1122 188
rect 1174 136 1246 188
rect 1298 136 1370 188
rect 1422 136 1494 188
rect 1546 136 1584 188
rect 340 64 1584 136
rect 340 12 378 64
rect 430 12 502 64
rect 554 12 626 64
rect 678 12 750 64
rect 802 12 874 64
rect 926 12 998 64
rect 1050 12 1122 64
rect 1174 12 1246 64
rect 1298 12 1370 64
rect 1422 12 1494 64
rect 1546 12 1584 64
rect 340 0 1584 12
<< via1 >>
rect 0 11916 156 11968
rect 0 11792 156 11844
rect 0 11668 156 11720
rect 0 11544 156 11596
rect 0 11420 156 11472
rect 0 11296 156 11348
rect 0 11172 156 11224
rect 0 11048 156 11100
rect 0 10924 156 10976
rect 0 10800 156 10852
rect 0 10676 156 10728
rect 0 10552 156 10604
rect 0 10428 156 10480
rect 0 10304 156 10356
rect 0 10180 156 10232
rect 0 10056 156 10108
rect 0 9932 156 9984
rect 0 9808 156 9860
rect 0 9684 156 9736
rect 0 9560 156 9612
rect 0 9436 156 9488
rect 0 9312 156 9364
rect 0 9188 156 9240
rect 0 9064 156 9116
rect 0 8940 156 8992
rect 0 8816 156 8868
rect 0 8692 156 8744
rect 0 8568 156 8620
rect 0 8444 156 8496
rect 0 8320 156 8372
rect 0 8196 156 8248
rect 0 8072 156 8124
rect 0 7948 156 8000
rect 0 7824 156 7876
rect 0 7700 156 7752
rect 0 7576 156 7628
rect 0 7452 156 7504
rect 0 7328 156 7380
rect 0 7204 156 7256
rect 0 7080 156 7132
rect 0 6956 156 7008
rect 0 6832 156 6884
rect 0 6708 156 6760
rect 0 6584 156 6636
rect 0 6460 156 6512
rect 0 6336 156 6388
rect 0 6212 156 6264
rect 0 6088 156 6140
rect 0 5964 156 6016
rect 0 5840 156 5892
rect 0 5716 156 5768
rect 0 5592 156 5644
rect 0 5468 156 5520
rect 0 5344 156 5396
rect 0 5220 156 5272
rect 0 5096 156 5148
rect 0 4972 156 5024
rect 0 4848 156 4900
rect 0 4724 156 4776
rect 0 4600 156 4652
rect 0 4476 156 4528
rect 0 4352 156 4404
rect 0 4228 156 4280
rect 0 4104 156 4156
rect 0 3980 156 4032
rect 0 3856 156 3908
rect 0 3732 156 3784
rect 0 3608 156 3660
rect 0 3484 156 3536
rect 0 3360 156 3412
rect 0 3236 156 3288
rect 0 3112 156 3164
rect 0 2988 156 3040
rect 0 2864 156 2916
rect 0 2740 156 2792
rect 0 2616 156 2668
rect 0 2492 156 2544
rect 0 2368 156 2420
rect 0 2244 156 2296
rect 0 2120 156 2172
rect 0 1996 156 2048
rect 0 1872 156 1924
rect 0 1748 156 1800
rect 0 1624 156 1676
rect 0 1500 156 1552
rect 0 1376 156 1428
rect 0 1252 156 1304
rect 0 1128 156 1180
rect 0 1004 156 1056
rect 0 880 156 932
rect 0 756 156 808
rect 0 632 156 684
rect 0 508 156 560
rect 0 384 156 436
rect 0 260 156 312
rect 0 136 156 188
rect 0 12 156 64
rect 378 11916 430 11968
rect 502 11916 554 11968
rect 626 11916 678 11968
rect 750 11916 802 11968
rect 874 11916 926 11968
rect 998 11916 1050 11968
rect 1122 11916 1174 11968
rect 1246 11916 1298 11968
rect 1370 11916 1422 11968
rect 1494 11916 1546 11968
rect 378 11792 430 11844
rect 502 11792 554 11844
rect 626 11792 678 11844
rect 750 11792 802 11844
rect 874 11792 926 11844
rect 998 11792 1050 11844
rect 1122 11792 1174 11844
rect 1246 11792 1298 11844
rect 1370 11792 1422 11844
rect 1494 11792 1546 11844
rect 378 11668 430 11720
rect 502 11668 554 11720
rect 626 11668 678 11720
rect 750 11668 802 11720
rect 874 11668 926 11720
rect 998 11668 1050 11720
rect 1122 11668 1174 11720
rect 1246 11668 1298 11720
rect 1370 11668 1422 11720
rect 1494 11668 1546 11720
rect 378 11544 430 11596
rect 502 11544 554 11596
rect 626 11544 678 11596
rect 750 11544 802 11596
rect 874 11544 926 11596
rect 998 11544 1050 11596
rect 1122 11544 1174 11596
rect 1246 11544 1298 11596
rect 1370 11544 1422 11596
rect 1494 11544 1546 11596
rect 378 11420 430 11472
rect 502 11420 554 11472
rect 626 11420 678 11472
rect 750 11420 802 11472
rect 874 11420 926 11472
rect 998 11420 1050 11472
rect 1122 11420 1174 11472
rect 1246 11420 1298 11472
rect 1370 11420 1422 11472
rect 1494 11420 1546 11472
rect 378 11296 430 11348
rect 502 11296 554 11348
rect 626 11296 678 11348
rect 750 11296 802 11348
rect 874 11296 926 11348
rect 998 11296 1050 11348
rect 1122 11296 1174 11348
rect 1246 11296 1298 11348
rect 1370 11296 1422 11348
rect 1494 11296 1546 11348
rect 378 11172 430 11224
rect 502 11172 554 11224
rect 626 11172 678 11224
rect 750 11172 802 11224
rect 874 11172 926 11224
rect 998 11172 1050 11224
rect 1122 11172 1174 11224
rect 1246 11172 1298 11224
rect 1370 11172 1422 11224
rect 1494 11172 1546 11224
rect 378 11048 430 11100
rect 502 11048 554 11100
rect 626 11048 678 11100
rect 750 11048 802 11100
rect 874 11048 926 11100
rect 998 11048 1050 11100
rect 1122 11048 1174 11100
rect 1246 11048 1298 11100
rect 1370 11048 1422 11100
rect 1494 11048 1546 11100
rect 378 10924 430 10976
rect 502 10924 554 10976
rect 626 10924 678 10976
rect 750 10924 802 10976
rect 874 10924 926 10976
rect 998 10924 1050 10976
rect 1122 10924 1174 10976
rect 1246 10924 1298 10976
rect 1370 10924 1422 10976
rect 1494 10924 1546 10976
rect 378 10800 430 10852
rect 502 10800 554 10852
rect 626 10800 678 10852
rect 750 10800 802 10852
rect 874 10800 926 10852
rect 998 10800 1050 10852
rect 1122 10800 1174 10852
rect 1246 10800 1298 10852
rect 1370 10800 1422 10852
rect 1494 10800 1546 10852
rect 378 10676 430 10728
rect 502 10676 554 10728
rect 626 10676 678 10728
rect 750 10676 802 10728
rect 874 10676 926 10728
rect 998 10676 1050 10728
rect 1122 10676 1174 10728
rect 1246 10676 1298 10728
rect 1370 10676 1422 10728
rect 1494 10676 1546 10728
rect 378 10552 430 10604
rect 502 10552 554 10604
rect 626 10552 678 10604
rect 750 10552 802 10604
rect 874 10552 926 10604
rect 998 10552 1050 10604
rect 1122 10552 1174 10604
rect 1246 10552 1298 10604
rect 1370 10552 1422 10604
rect 1494 10552 1546 10604
rect 378 10428 430 10480
rect 502 10428 554 10480
rect 626 10428 678 10480
rect 750 10428 802 10480
rect 874 10428 926 10480
rect 998 10428 1050 10480
rect 1122 10428 1174 10480
rect 1246 10428 1298 10480
rect 1370 10428 1422 10480
rect 1494 10428 1546 10480
rect 378 10304 430 10356
rect 502 10304 554 10356
rect 626 10304 678 10356
rect 750 10304 802 10356
rect 874 10304 926 10356
rect 998 10304 1050 10356
rect 1122 10304 1174 10356
rect 1246 10304 1298 10356
rect 1370 10304 1422 10356
rect 1494 10304 1546 10356
rect 378 10180 430 10232
rect 502 10180 554 10232
rect 626 10180 678 10232
rect 750 10180 802 10232
rect 874 10180 926 10232
rect 998 10180 1050 10232
rect 1122 10180 1174 10232
rect 1246 10180 1298 10232
rect 1370 10180 1422 10232
rect 1494 10180 1546 10232
rect 378 10056 430 10108
rect 502 10056 554 10108
rect 626 10056 678 10108
rect 750 10056 802 10108
rect 874 10056 926 10108
rect 998 10056 1050 10108
rect 1122 10056 1174 10108
rect 1246 10056 1298 10108
rect 1370 10056 1422 10108
rect 1494 10056 1546 10108
rect 378 9932 430 9984
rect 502 9932 554 9984
rect 626 9932 678 9984
rect 750 9932 802 9984
rect 874 9932 926 9984
rect 998 9932 1050 9984
rect 1122 9932 1174 9984
rect 1246 9932 1298 9984
rect 1370 9932 1422 9984
rect 1494 9932 1546 9984
rect 378 9808 430 9860
rect 502 9808 554 9860
rect 626 9808 678 9860
rect 750 9808 802 9860
rect 874 9808 926 9860
rect 998 9808 1050 9860
rect 1122 9808 1174 9860
rect 1246 9808 1298 9860
rect 1370 9808 1422 9860
rect 1494 9808 1546 9860
rect 378 9684 430 9736
rect 502 9684 554 9736
rect 626 9684 678 9736
rect 750 9684 802 9736
rect 874 9684 926 9736
rect 998 9684 1050 9736
rect 1122 9684 1174 9736
rect 1246 9684 1298 9736
rect 1370 9684 1422 9736
rect 1494 9684 1546 9736
rect 378 9560 430 9612
rect 502 9560 554 9612
rect 626 9560 678 9612
rect 750 9560 802 9612
rect 874 9560 926 9612
rect 998 9560 1050 9612
rect 1122 9560 1174 9612
rect 1246 9560 1298 9612
rect 1370 9560 1422 9612
rect 1494 9560 1546 9612
rect 378 9436 430 9488
rect 502 9436 554 9488
rect 626 9436 678 9488
rect 750 9436 802 9488
rect 874 9436 926 9488
rect 998 9436 1050 9488
rect 1122 9436 1174 9488
rect 1246 9436 1298 9488
rect 1370 9436 1422 9488
rect 1494 9436 1546 9488
rect 378 9312 430 9364
rect 502 9312 554 9364
rect 626 9312 678 9364
rect 750 9312 802 9364
rect 874 9312 926 9364
rect 998 9312 1050 9364
rect 1122 9312 1174 9364
rect 1246 9312 1298 9364
rect 1370 9312 1422 9364
rect 1494 9312 1546 9364
rect 378 9188 430 9240
rect 502 9188 554 9240
rect 626 9188 678 9240
rect 750 9188 802 9240
rect 874 9188 926 9240
rect 998 9188 1050 9240
rect 1122 9188 1174 9240
rect 1246 9188 1298 9240
rect 1370 9188 1422 9240
rect 1494 9188 1546 9240
rect 378 9064 430 9116
rect 502 9064 554 9116
rect 626 9064 678 9116
rect 750 9064 802 9116
rect 874 9064 926 9116
rect 998 9064 1050 9116
rect 1122 9064 1174 9116
rect 1246 9064 1298 9116
rect 1370 9064 1422 9116
rect 1494 9064 1546 9116
rect 378 8940 430 8992
rect 502 8940 554 8992
rect 626 8940 678 8992
rect 750 8940 802 8992
rect 874 8940 926 8992
rect 998 8940 1050 8992
rect 1122 8940 1174 8992
rect 1246 8940 1298 8992
rect 1370 8940 1422 8992
rect 1494 8940 1546 8992
rect 378 8816 430 8868
rect 502 8816 554 8868
rect 626 8816 678 8868
rect 750 8816 802 8868
rect 874 8816 926 8868
rect 998 8816 1050 8868
rect 1122 8816 1174 8868
rect 1246 8816 1298 8868
rect 1370 8816 1422 8868
rect 1494 8816 1546 8868
rect 378 8692 430 8744
rect 502 8692 554 8744
rect 626 8692 678 8744
rect 750 8692 802 8744
rect 874 8692 926 8744
rect 998 8692 1050 8744
rect 1122 8692 1174 8744
rect 1246 8692 1298 8744
rect 1370 8692 1422 8744
rect 1494 8692 1546 8744
rect 378 8568 430 8620
rect 502 8568 554 8620
rect 626 8568 678 8620
rect 750 8568 802 8620
rect 874 8568 926 8620
rect 998 8568 1050 8620
rect 1122 8568 1174 8620
rect 1246 8568 1298 8620
rect 1370 8568 1422 8620
rect 1494 8568 1546 8620
rect 378 8444 430 8496
rect 502 8444 554 8496
rect 626 8444 678 8496
rect 750 8444 802 8496
rect 874 8444 926 8496
rect 998 8444 1050 8496
rect 1122 8444 1174 8496
rect 1246 8444 1298 8496
rect 1370 8444 1422 8496
rect 1494 8444 1546 8496
rect 378 8320 430 8372
rect 502 8320 554 8372
rect 626 8320 678 8372
rect 750 8320 802 8372
rect 874 8320 926 8372
rect 998 8320 1050 8372
rect 1122 8320 1174 8372
rect 1246 8320 1298 8372
rect 1370 8320 1422 8372
rect 1494 8320 1546 8372
rect 378 8196 430 8248
rect 502 8196 554 8248
rect 626 8196 678 8248
rect 750 8196 802 8248
rect 874 8196 926 8248
rect 998 8196 1050 8248
rect 1122 8196 1174 8248
rect 1246 8196 1298 8248
rect 1370 8196 1422 8248
rect 1494 8196 1546 8248
rect 378 8072 430 8124
rect 502 8072 554 8124
rect 626 8072 678 8124
rect 750 8072 802 8124
rect 874 8072 926 8124
rect 998 8072 1050 8124
rect 1122 8072 1174 8124
rect 1246 8072 1298 8124
rect 1370 8072 1422 8124
rect 1494 8072 1546 8124
rect 378 7948 430 8000
rect 502 7948 554 8000
rect 626 7948 678 8000
rect 750 7948 802 8000
rect 874 7948 926 8000
rect 998 7948 1050 8000
rect 1122 7948 1174 8000
rect 1246 7948 1298 8000
rect 1370 7948 1422 8000
rect 1494 7948 1546 8000
rect 378 7824 430 7876
rect 502 7824 554 7876
rect 626 7824 678 7876
rect 750 7824 802 7876
rect 874 7824 926 7876
rect 998 7824 1050 7876
rect 1122 7824 1174 7876
rect 1246 7824 1298 7876
rect 1370 7824 1422 7876
rect 1494 7824 1546 7876
rect 378 7700 430 7752
rect 502 7700 554 7752
rect 626 7700 678 7752
rect 750 7700 802 7752
rect 874 7700 926 7752
rect 998 7700 1050 7752
rect 1122 7700 1174 7752
rect 1246 7700 1298 7752
rect 1370 7700 1422 7752
rect 1494 7700 1546 7752
rect 378 7576 430 7628
rect 502 7576 554 7628
rect 626 7576 678 7628
rect 750 7576 802 7628
rect 874 7576 926 7628
rect 998 7576 1050 7628
rect 1122 7576 1174 7628
rect 1246 7576 1298 7628
rect 1370 7576 1422 7628
rect 1494 7576 1546 7628
rect 378 7452 430 7504
rect 502 7452 554 7504
rect 626 7452 678 7504
rect 750 7452 802 7504
rect 874 7452 926 7504
rect 998 7452 1050 7504
rect 1122 7452 1174 7504
rect 1246 7452 1298 7504
rect 1370 7452 1422 7504
rect 1494 7452 1546 7504
rect 378 7328 430 7380
rect 502 7328 554 7380
rect 626 7328 678 7380
rect 750 7328 802 7380
rect 874 7328 926 7380
rect 998 7328 1050 7380
rect 1122 7328 1174 7380
rect 1246 7328 1298 7380
rect 1370 7328 1422 7380
rect 1494 7328 1546 7380
rect 378 7204 430 7256
rect 502 7204 554 7256
rect 626 7204 678 7256
rect 750 7204 802 7256
rect 874 7204 926 7256
rect 998 7204 1050 7256
rect 1122 7204 1174 7256
rect 1246 7204 1298 7256
rect 1370 7204 1422 7256
rect 1494 7204 1546 7256
rect 378 7080 430 7132
rect 502 7080 554 7132
rect 626 7080 678 7132
rect 750 7080 802 7132
rect 874 7080 926 7132
rect 998 7080 1050 7132
rect 1122 7080 1174 7132
rect 1246 7080 1298 7132
rect 1370 7080 1422 7132
rect 1494 7080 1546 7132
rect 378 6956 430 7008
rect 502 6956 554 7008
rect 626 6956 678 7008
rect 750 6956 802 7008
rect 874 6956 926 7008
rect 998 6956 1050 7008
rect 1122 6956 1174 7008
rect 1246 6956 1298 7008
rect 1370 6956 1422 7008
rect 1494 6956 1546 7008
rect 378 6832 430 6884
rect 502 6832 554 6884
rect 626 6832 678 6884
rect 750 6832 802 6884
rect 874 6832 926 6884
rect 998 6832 1050 6884
rect 1122 6832 1174 6884
rect 1246 6832 1298 6884
rect 1370 6832 1422 6884
rect 1494 6832 1546 6884
rect 378 6708 430 6760
rect 502 6708 554 6760
rect 626 6708 678 6760
rect 750 6708 802 6760
rect 874 6708 926 6760
rect 998 6708 1050 6760
rect 1122 6708 1174 6760
rect 1246 6708 1298 6760
rect 1370 6708 1422 6760
rect 1494 6708 1546 6760
rect 378 6584 430 6636
rect 502 6584 554 6636
rect 626 6584 678 6636
rect 750 6584 802 6636
rect 874 6584 926 6636
rect 998 6584 1050 6636
rect 1122 6584 1174 6636
rect 1246 6584 1298 6636
rect 1370 6584 1422 6636
rect 1494 6584 1546 6636
rect 378 6460 430 6512
rect 502 6460 554 6512
rect 626 6460 678 6512
rect 750 6460 802 6512
rect 874 6460 926 6512
rect 998 6460 1050 6512
rect 1122 6460 1174 6512
rect 1246 6460 1298 6512
rect 1370 6460 1422 6512
rect 1494 6460 1546 6512
rect 378 6336 430 6388
rect 502 6336 554 6388
rect 626 6336 678 6388
rect 750 6336 802 6388
rect 874 6336 926 6388
rect 998 6336 1050 6388
rect 1122 6336 1174 6388
rect 1246 6336 1298 6388
rect 1370 6336 1422 6388
rect 1494 6336 1546 6388
rect 378 6212 430 6264
rect 502 6212 554 6264
rect 626 6212 678 6264
rect 750 6212 802 6264
rect 874 6212 926 6264
rect 998 6212 1050 6264
rect 1122 6212 1174 6264
rect 1246 6212 1298 6264
rect 1370 6212 1422 6264
rect 1494 6212 1546 6264
rect 378 6088 430 6140
rect 502 6088 554 6140
rect 626 6088 678 6140
rect 750 6088 802 6140
rect 874 6088 926 6140
rect 998 6088 1050 6140
rect 1122 6088 1174 6140
rect 1246 6088 1298 6140
rect 1370 6088 1422 6140
rect 1494 6088 1546 6140
rect 378 5964 430 6016
rect 502 5964 554 6016
rect 626 5964 678 6016
rect 750 5964 802 6016
rect 874 5964 926 6016
rect 998 5964 1050 6016
rect 1122 5964 1174 6016
rect 1246 5964 1298 6016
rect 1370 5964 1422 6016
rect 1494 5964 1546 6016
rect 378 5840 430 5892
rect 502 5840 554 5892
rect 626 5840 678 5892
rect 750 5840 802 5892
rect 874 5840 926 5892
rect 998 5840 1050 5892
rect 1122 5840 1174 5892
rect 1246 5840 1298 5892
rect 1370 5840 1422 5892
rect 1494 5840 1546 5892
rect 378 5716 430 5768
rect 502 5716 554 5768
rect 626 5716 678 5768
rect 750 5716 802 5768
rect 874 5716 926 5768
rect 998 5716 1050 5768
rect 1122 5716 1174 5768
rect 1246 5716 1298 5768
rect 1370 5716 1422 5768
rect 1494 5716 1546 5768
rect 378 5592 430 5644
rect 502 5592 554 5644
rect 626 5592 678 5644
rect 750 5592 802 5644
rect 874 5592 926 5644
rect 998 5592 1050 5644
rect 1122 5592 1174 5644
rect 1246 5592 1298 5644
rect 1370 5592 1422 5644
rect 1494 5592 1546 5644
rect 378 5468 430 5520
rect 502 5468 554 5520
rect 626 5468 678 5520
rect 750 5468 802 5520
rect 874 5468 926 5520
rect 998 5468 1050 5520
rect 1122 5468 1174 5520
rect 1246 5468 1298 5520
rect 1370 5468 1422 5520
rect 1494 5468 1546 5520
rect 378 5344 430 5396
rect 502 5344 554 5396
rect 626 5344 678 5396
rect 750 5344 802 5396
rect 874 5344 926 5396
rect 998 5344 1050 5396
rect 1122 5344 1174 5396
rect 1246 5344 1298 5396
rect 1370 5344 1422 5396
rect 1494 5344 1546 5396
rect 378 5220 430 5272
rect 502 5220 554 5272
rect 626 5220 678 5272
rect 750 5220 802 5272
rect 874 5220 926 5272
rect 998 5220 1050 5272
rect 1122 5220 1174 5272
rect 1246 5220 1298 5272
rect 1370 5220 1422 5272
rect 1494 5220 1546 5272
rect 378 5096 430 5148
rect 502 5096 554 5148
rect 626 5096 678 5148
rect 750 5096 802 5148
rect 874 5096 926 5148
rect 998 5096 1050 5148
rect 1122 5096 1174 5148
rect 1246 5096 1298 5148
rect 1370 5096 1422 5148
rect 1494 5096 1546 5148
rect 378 4972 430 5024
rect 502 4972 554 5024
rect 626 4972 678 5024
rect 750 4972 802 5024
rect 874 4972 926 5024
rect 998 4972 1050 5024
rect 1122 4972 1174 5024
rect 1246 4972 1298 5024
rect 1370 4972 1422 5024
rect 1494 4972 1546 5024
rect 378 4848 430 4900
rect 502 4848 554 4900
rect 626 4848 678 4900
rect 750 4848 802 4900
rect 874 4848 926 4900
rect 998 4848 1050 4900
rect 1122 4848 1174 4900
rect 1246 4848 1298 4900
rect 1370 4848 1422 4900
rect 1494 4848 1546 4900
rect 378 4724 430 4776
rect 502 4724 554 4776
rect 626 4724 678 4776
rect 750 4724 802 4776
rect 874 4724 926 4776
rect 998 4724 1050 4776
rect 1122 4724 1174 4776
rect 1246 4724 1298 4776
rect 1370 4724 1422 4776
rect 1494 4724 1546 4776
rect 378 4600 430 4652
rect 502 4600 554 4652
rect 626 4600 678 4652
rect 750 4600 802 4652
rect 874 4600 926 4652
rect 998 4600 1050 4652
rect 1122 4600 1174 4652
rect 1246 4600 1298 4652
rect 1370 4600 1422 4652
rect 1494 4600 1546 4652
rect 378 4476 430 4528
rect 502 4476 554 4528
rect 626 4476 678 4528
rect 750 4476 802 4528
rect 874 4476 926 4528
rect 998 4476 1050 4528
rect 1122 4476 1174 4528
rect 1246 4476 1298 4528
rect 1370 4476 1422 4528
rect 1494 4476 1546 4528
rect 378 4352 430 4404
rect 502 4352 554 4404
rect 626 4352 678 4404
rect 750 4352 802 4404
rect 874 4352 926 4404
rect 998 4352 1050 4404
rect 1122 4352 1174 4404
rect 1246 4352 1298 4404
rect 1370 4352 1422 4404
rect 1494 4352 1546 4404
rect 378 4228 430 4280
rect 502 4228 554 4280
rect 626 4228 678 4280
rect 750 4228 802 4280
rect 874 4228 926 4280
rect 998 4228 1050 4280
rect 1122 4228 1174 4280
rect 1246 4228 1298 4280
rect 1370 4228 1422 4280
rect 1494 4228 1546 4280
rect 378 4104 430 4156
rect 502 4104 554 4156
rect 626 4104 678 4156
rect 750 4104 802 4156
rect 874 4104 926 4156
rect 998 4104 1050 4156
rect 1122 4104 1174 4156
rect 1246 4104 1298 4156
rect 1370 4104 1422 4156
rect 1494 4104 1546 4156
rect 378 3980 430 4032
rect 502 3980 554 4032
rect 626 3980 678 4032
rect 750 3980 802 4032
rect 874 3980 926 4032
rect 998 3980 1050 4032
rect 1122 3980 1174 4032
rect 1246 3980 1298 4032
rect 1370 3980 1422 4032
rect 1494 3980 1546 4032
rect 378 3856 430 3908
rect 502 3856 554 3908
rect 626 3856 678 3908
rect 750 3856 802 3908
rect 874 3856 926 3908
rect 998 3856 1050 3908
rect 1122 3856 1174 3908
rect 1246 3856 1298 3908
rect 1370 3856 1422 3908
rect 1494 3856 1546 3908
rect 378 3732 430 3784
rect 502 3732 554 3784
rect 626 3732 678 3784
rect 750 3732 802 3784
rect 874 3732 926 3784
rect 998 3732 1050 3784
rect 1122 3732 1174 3784
rect 1246 3732 1298 3784
rect 1370 3732 1422 3784
rect 1494 3732 1546 3784
rect 378 3608 430 3660
rect 502 3608 554 3660
rect 626 3608 678 3660
rect 750 3608 802 3660
rect 874 3608 926 3660
rect 998 3608 1050 3660
rect 1122 3608 1174 3660
rect 1246 3608 1298 3660
rect 1370 3608 1422 3660
rect 1494 3608 1546 3660
rect 378 3484 430 3536
rect 502 3484 554 3536
rect 626 3484 678 3536
rect 750 3484 802 3536
rect 874 3484 926 3536
rect 998 3484 1050 3536
rect 1122 3484 1174 3536
rect 1246 3484 1298 3536
rect 1370 3484 1422 3536
rect 1494 3484 1546 3536
rect 378 3360 430 3412
rect 502 3360 554 3412
rect 626 3360 678 3412
rect 750 3360 802 3412
rect 874 3360 926 3412
rect 998 3360 1050 3412
rect 1122 3360 1174 3412
rect 1246 3360 1298 3412
rect 1370 3360 1422 3412
rect 1494 3360 1546 3412
rect 378 3236 430 3288
rect 502 3236 554 3288
rect 626 3236 678 3288
rect 750 3236 802 3288
rect 874 3236 926 3288
rect 998 3236 1050 3288
rect 1122 3236 1174 3288
rect 1246 3236 1298 3288
rect 1370 3236 1422 3288
rect 1494 3236 1546 3288
rect 378 3112 430 3164
rect 502 3112 554 3164
rect 626 3112 678 3164
rect 750 3112 802 3164
rect 874 3112 926 3164
rect 998 3112 1050 3164
rect 1122 3112 1174 3164
rect 1246 3112 1298 3164
rect 1370 3112 1422 3164
rect 1494 3112 1546 3164
rect 378 2988 430 3040
rect 502 2988 554 3040
rect 626 2988 678 3040
rect 750 2988 802 3040
rect 874 2988 926 3040
rect 998 2988 1050 3040
rect 1122 2988 1174 3040
rect 1246 2988 1298 3040
rect 1370 2988 1422 3040
rect 1494 2988 1546 3040
rect 378 2864 430 2916
rect 502 2864 554 2916
rect 626 2864 678 2916
rect 750 2864 802 2916
rect 874 2864 926 2916
rect 998 2864 1050 2916
rect 1122 2864 1174 2916
rect 1246 2864 1298 2916
rect 1370 2864 1422 2916
rect 1494 2864 1546 2916
rect 378 2740 430 2792
rect 502 2740 554 2792
rect 626 2740 678 2792
rect 750 2740 802 2792
rect 874 2740 926 2792
rect 998 2740 1050 2792
rect 1122 2740 1174 2792
rect 1246 2740 1298 2792
rect 1370 2740 1422 2792
rect 1494 2740 1546 2792
rect 378 2616 430 2668
rect 502 2616 554 2668
rect 626 2616 678 2668
rect 750 2616 802 2668
rect 874 2616 926 2668
rect 998 2616 1050 2668
rect 1122 2616 1174 2668
rect 1246 2616 1298 2668
rect 1370 2616 1422 2668
rect 1494 2616 1546 2668
rect 378 2492 430 2544
rect 502 2492 554 2544
rect 626 2492 678 2544
rect 750 2492 802 2544
rect 874 2492 926 2544
rect 998 2492 1050 2544
rect 1122 2492 1174 2544
rect 1246 2492 1298 2544
rect 1370 2492 1422 2544
rect 1494 2492 1546 2544
rect 378 2368 430 2420
rect 502 2368 554 2420
rect 626 2368 678 2420
rect 750 2368 802 2420
rect 874 2368 926 2420
rect 998 2368 1050 2420
rect 1122 2368 1174 2420
rect 1246 2368 1298 2420
rect 1370 2368 1422 2420
rect 1494 2368 1546 2420
rect 378 2244 430 2296
rect 502 2244 554 2296
rect 626 2244 678 2296
rect 750 2244 802 2296
rect 874 2244 926 2296
rect 998 2244 1050 2296
rect 1122 2244 1174 2296
rect 1246 2244 1298 2296
rect 1370 2244 1422 2296
rect 1494 2244 1546 2296
rect 378 2120 430 2172
rect 502 2120 554 2172
rect 626 2120 678 2172
rect 750 2120 802 2172
rect 874 2120 926 2172
rect 998 2120 1050 2172
rect 1122 2120 1174 2172
rect 1246 2120 1298 2172
rect 1370 2120 1422 2172
rect 1494 2120 1546 2172
rect 378 1996 430 2048
rect 502 1996 554 2048
rect 626 1996 678 2048
rect 750 1996 802 2048
rect 874 1996 926 2048
rect 998 1996 1050 2048
rect 1122 1996 1174 2048
rect 1246 1996 1298 2048
rect 1370 1996 1422 2048
rect 1494 1996 1546 2048
rect 378 1872 430 1924
rect 502 1872 554 1924
rect 626 1872 678 1924
rect 750 1872 802 1924
rect 874 1872 926 1924
rect 998 1872 1050 1924
rect 1122 1872 1174 1924
rect 1246 1872 1298 1924
rect 1370 1872 1422 1924
rect 1494 1872 1546 1924
rect 378 1748 430 1800
rect 502 1748 554 1800
rect 626 1748 678 1800
rect 750 1748 802 1800
rect 874 1748 926 1800
rect 998 1748 1050 1800
rect 1122 1748 1174 1800
rect 1246 1748 1298 1800
rect 1370 1748 1422 1800
rect 1494 1748 1546 1800
rect 378 1624 430 1676
rect 502 1624 554 1676
rect 626 1624 678 1676
rect 750 1624 802 1676
rect 874 1624 926 1676
rect 998 1624 1050 1676
rect 1122 1624 1174 1676
rect 1246 1624 1298 1676
rect 1370 1624 1422 1676
rect 1494 1624 1546 1676
rect 378 1500 430 1552
rect 502 1500 554 1552
rect 626 1500 678 1552
rect 750 1500 802 1552
rect 874 1500 926 1552
rect 998 1500 1050 1552
rect 1122 1500 1174 1552
rect 1246 1500 1298 1552
rect 1370 1500 1422 1552
rect 1494 1500 1546 1552
rect 378 1376 430 1428
rect 502 1376 554 1428
rect 626 1376 678 1428
rect 750 1376 802 1428
rect 874 1376 926 1428
rect 998 1376 1050 1428
rect 1122 1376 1174 1428
rect 1246 1376 1298 1428
rect 1370 1376 1422 1428
rect 1494 1376 1546 1428
rect 378 1252 430 1304
rect 502 1252 554 1304
rect 626 1252 678 1304
rect 750 1252 802 1304
rect 874 1252 926 1304
rect 998 1252 1050 1304
rect 1122 1252 1174 1304
rect 1246 1252 1298 1304
rect 1370 1252 1422 1304
rect 1494 1252 1546 1304
rect 378 1128 430 1180
rect 502 1128 554 1180
rect 626 1128 678 1180
rect 750 1128 802 1180
rect 874 1128 926 1180
rect 998 1128 1050 1180
rect 1122 1128 1174 1180
rect 1246 1128 1298 1180
rect 1370 1128 1422 1180
rect 1494 1128 1546 1180
rect 378 1004 430 1056
rect 502 1004 554 1056
rect 626 1004 678 1056
rect 750 1004 802 1056
rect 874 1004 926 1056
rect 998 1004 1050 1056
rect 1122 1004 1174 1056
rect 1246 1004 1298 1056
rect 1370 1004 1422 1056
rect 1494 1004 1546 1056
rect 378 880 430 932
rect 502 880 554 932
rect 626 880 678 932
rect 750 880 802 932
rect 874 880 926 932
rect 998 880 1050 932
rect 1122 880 1174 932
rect 1246 880 1298 932
rect 1370 880 1422 932
rect 1494 880 1546 932
rect 378 756 430 808
rect 502 756 554 808
rect 626 756 678 808
rect 750 756 802 808
rect 874 756 926 808
rect 998 756 1050 808
rect 1122 756 1174 808
rect 1246 756 1298 808
rect 1370 756 1422 808
rect 1494 756 1546 808
rect 378 632 430 684
rect 502 632 554 684
rect 626 632 678 684
rect 750 632 802 684
rect 874 632 926 684
rect 998 632 1050 684
rect 1122 632 1174 684
rect 1246 632 1298 684
rect 1370 632 1422 684
rect 1494 632 1546 684
rect 378 508 430 560
rect 502 508 554 560
rect 626 508 678 560
rect 750 508 802 560
rect 874 508 926 560
rect 998 508 1050 560
rect 1122 508 1174 560
rect 1246 508 1298 560
rect 1370 508 1422 560
rect 1494 508 1546 560
rect 378 384 430 436
rect 502 384 554 436
rect 626 384 678 436
rect 750 384 802 436
rect 874 384 926 436
rect 998 384 1050 436
rect 1122 384 1174 436
rect 1246 384 1298 436
rect 1370 384 1422 436
rect 1494 384 1546 436
rect 378 260 430 312
rect 502 260 554 312
rect 626 260 678 312
rect 750 260 802 312
rect 874 260 926 312
rect 998 260 1050 312
rect 1122 260 1174 312
rect 1246 260 1298 312
rect 1370 260 1422 312
rect 1494 260 1546 312
rect 378 136 430 188
rect 502 136 554 188
rect 626 136 678 188
rect 750 136 802 188
rect 874 136 926 188
rect 998 136 1050 188
rect 1122 136 1174 188
rect 1246 136 1298 188
rect 1370 136 1422 188
rect 1494 136 1546 188
rect 378 12 430 64
rect 502 12 554 64
rect 626 12 678 64
rect 750 12 802 64
rect 874 12 926 64
rect 998 12 1050 64
rect 1122 12 1174 64
rect 1246 12 1298 64
rect 1370 12 1422 64
rect 1494 12 1546 64
<< metal2 >>
rect -44 11968 200 12000
rect -44 11938 0 11968
rect 156 11938 200 11968
rect -44 11882 -22 11938
rect 34 11882 120 11916
rect 176 11882 200 11938
rect -44 11844 200 11882
rect -44 11796 0 11844
rect 156 11796 200 11844
rect -44 11740 -22 11796
rect 34 11740 120 11792
rect 176 11740 200 11796
rect -44 11720 200 11740
rect -44 11668 0 11720
rect 156 11668 200 11720
rect -44 11654 200 11668
rect -44 11598 -22 11654
rect 34 11598 120 11654
rect 176 11598 200 11654
rect -44 11596 200 11598
rect -44 11544 0 11596
rect 156 11544 200 11596
rect -44 11512 200 11544
rect -44 11456 -22 11512
rect 34 11472 120 11512
rect 176 11456 200 11512
rect -44 11420 0 11456
rect 156 11420 200 11456
rect -44 11370 200 11420
rect -44 11314 -22 11370
rect 34 11348 120 11370
rect 176 11314 200 11370
rect -44 11296 0 11314
rect 156 11296 200 11314
rect -44 11228 200 11296
rect -44 11172 -22 11228
rect 34 11224 120 11228
rect 176 11172 200 11228
rect -44 11100 200 11172
rect -44 11086 0 11100
rect 156 11086 200 11100
rect -44 11030 -22 11086
rect 34 11030 120 11048
rect 176 11030 200 11086
rect -44 10976 200 11030
rect -44 10944 0 10976
rect 156 10944 200 10976
rect -44 10888 -22 10944
rect 34 10888 120 10924
rect 176 10888 200 10944
rect -44 10852 200 10888
rect -44 10802 0 10852
rect 156 10802 200 10852
rect -44 10746 -22 10802
rect 34 10746 120 10800
rect 176 10746 200 10802
rect -44 10728 200 10746
rect -44 10676 0 10728
rect 156 10676 200 10728
rect -44 10660 200 10676
rect -44 10604 -22 10660
rect 34 10604 120 10660
rect 176 10604 200 10660
rect -44 10552 0 10604
rect 156 10552 200 10604
rect -44 10518 200 10552
rect -44 10462 -22 10518
rect 34 10480 120 10518
rect 176 10462 200 10518
rect -44 10428 0 10462
rect 156 10428 200 10462
rect -44 10376 200 10428
rect -44 10320 -22 10376
rect 34 10356 120 10376
rect 176 10320 200 10376
rect -44 10304 0 10320
rect 156 10304 200 10320
rect -44 10234 200 10304
rect -44 10178 -22 10234
rect 34 10232 120 10234
rect 34 10178 120 10180
rect 176 10178 200 10234
rect -44 10108 200 10178
rect -44 10092 0 10108
rect 156 10092 200 10108
rect -44 10036 -22 10092
rect 34 10036 120 10056
rect 176 10036 200 10092
rect -44 9984 200 10036
rect -44 9950 0 9984
rect 156 9950 200 9984
rect -44 9894 -22 9950
rect 34 9894 120 9932
rect 176 9894 200 9950
rect -44 9860 200 9894
rect -44 9808 0 9860
rect 156 9808 200 9860
rect -44 9752 -22 9808
rect 34 9752 120 9808
rect 176 9752 200 9808
rect -44 9736 200 9752
rect -44 9684 0 9736
rect 156 9684 200 9736
rect -44 9612 200 9684
rect -44 9560 0 9612
rect 156 9560 200 9612
rect -44 9488 200 9560
rect -44 9436 0 9488
rect 156 9436 200 9488
rect -44 9426 200 9436
rect -44 9370 -22 9426
rect 34 9370 120 9426
rect 176 9370 200 9426
rect -44 9364 200 9370
rect -44 9312 0 9364
rect 156 9312 200 9364
rect -44 9284 200 9312
rect -44 9228 -22 9284
rect 34 9240 120 9284
rect 176 9228 200 9284
rect -44 9188 0 9228
rect 156 9188 200 9228
rect -44 9142 200 9188
rect -44 9086 -22 9142
rect 34 9116 120 9142
rect 176 9086 200 9142
rect -44 9064 0 9086
rect 156 9064 200 9086
rect -44 9000 200 9064
rect -44 8944 -22 9000
rect 34 8992 120 9000
rect 176 8944 200 9000
rect -44 8940 0 8944
rect 156 8940 200 8944
rect -44 8868 200 8940
rect -44 8858 0 8868
rect 156 8858 200 8868
rect -44 8802 -22 8858
rect 34 8802 120 8816
rect 176 8802 200 8858
rect -44 8744 200 8802
rect -44 8716 0 8744
rect 156 8716 200 8744
rect -44 8660 -22 8716
rect 34 8660 120 8692
rect 176 8660 200 8716
rect -44 8620 200 8660
rect -44 8574 0 8620
rect 156 8574 200 8620
rect -44 8518 -22 8574
rect 34 8518 120 8568
rect 176 8518 200 8574
rect -44 8496 200 8518
rect -44 8444 0 8496
rect 156 8444 200 8496
rect -44 8432 200 8444
rect -44 8376 -22 8432
rect 34 8376 120 8432
rect 176 8376 200 8432
rect -44 8372 200 8376
rect -44 8320 0 8372
rect 156 8320 200 8372
rect -44 8290 200 8320
rect -44 8234 -22 8290
rect 34 8248 120 8290
rect 176 8234 200 8290
rect -44 8196 0 8234
rect 156 8196 200 8234
rect -44 8148 200 8196
rect -44 8092 -22 8148
rect 34 8124 120 8148
rect 176 8092 200 8148
rect -44 8072 0 8092
rect 156 8072 200 8092
rect -44 8006 200 8072
rect -44 7950 -22 8006
rect 34 8000 120 8006
rect 176 7950 200 8006
rect -44 7948 0 7950
rect 156 7948 200 7950
rect -44 7876 200 7948
rect -44 7864 0 7876
rect 156 7864 200 7876
rect -44 7808 -22 7864
rect 34 7808 120 7824
rect 176 7808 200 7864
rect -44 7752 200 7808
rect -44 7722 0 7752
rect 156 7722 200 7752
rect -44 7666 -22 7722
rect 34 7666 120 7700
rect 176 7666 200 7722
rect -44 7628 200 7666
rect -44 7580 0 7628
rect 156 7580 200 7628
rect -44 7524 -22 7580
rect 34 7524 120 7576
rect 176 7524 200 7580
rect -44 7504 200 7524
rect -44 7452 0 7504
rect 156 7452 200 7504
rect -44 7438 200 7452
rect -44 7382 -22 7438
rect 34 7382 120 7438
rect 176 7382 200 7438
rect -44 7380 200 7382
rect -44 7328 0 7380
rect 156 7328 200 7380
rect -44 7296 200 7328
rect -44 7240 -22 7296
rect 34 7256 120 7296
rect 176 7240 200 7296
rect -44 7204 0 7240
rect 156 7204 200 7240
rect -44 7154 200 7204
rect -44 7098 -22 7154
rect 34 7132 120 7154
rect 176 7098 200 7154
rect -44 7080 0 7098
rect 156 7080 200 7098
rect -44 7012 200 7080
rect -44 6956 -22 7012
rect 34 7008 120 7012
rect 176 6956 200 7012
rect -44 6884 200 6956
rect -44 6870 0 6884
rect 156 6870 200 6884
rect -44 6814 -22 6870
rect 34 6814 120 6832
rect 176 6814 200 6870
rect -44 6760 200 6814
rect -44 6728 0 6760
rect 156 6728 200 6760
rect -44 6672 -22 6728
rect 34 6672 120 6708
rect 176 6672 200 6728
rect -44 6636 200 6672
rect -44 6586 0 6636
rect 156 6586 200 6636
rect -44 6530 -22 6586
rect 34 6530 120 6584
rect 176 6530 200 6586
rect -44 6512 200 6530
rect -44 6460 0 6512
rect 156 6460 200 6512
rect -44 6388 200 6460
rect -44 6336 0 6388
rect 156 6336 200 6388
rect -44 6264 200 6336
rect -44 6239 0 6264
rect 156 6239 200 6264
rect -44 6183 -22 6239
rect 34 6183 120 6212
rect 176 6183 200 6239
rect -44 6140 200 6183
rect -44 6097 0 6140
rect 156 6097 200 6140
rect -44 6041 -22 6097
rect 34 6041 120 6088
rect 176 6041 200 6097
rect -44 6016 200 6041
rect -44 5964 0 6016
rect 156 5964 200 6016
rect -44 5955 200 5964
rect -44 5899 -22 5955
rect 34 5899 120 5955
rect 176 5899 200 5955
rect -44 5892 200 5899
rect -44 5840 0 5892
rect 156 5840 200 5892
rect -44 5813 200 5840
rect -44 5757 -22 5813
rect 34 5768 120 5813
rect 176 5757 200 5813
rect -44 5716 0 5757
rect 156 5716 200 5757
rect -44 5671 200 5716
rect -44 5615 -22 5671
rect 34 5644 120 5671
rect 176 5615 200 5671
rect -44 5592 0 5615
rect 156 5592 200 5615
rect -44 5529 200 5592
rect -44 5473 -22 5529
rect 34 5520 120 5529
rect 176 5473 200 5529
rect -44 5468 0 5473
rect 156 5468 200 5473
rect -44 5396 200 5468
rect -44 5387 0 5396
rect 156 5387 200 5396
rect -44 5331 -22 5387
rect 34 5331 120 5344
rect 176 5331 200 5387
rect -44 5272 200 5331
rect -44 5245 0 5272
rect 156 5245 200 5272
rect -44 5189 -22 5245
rect 34 5189 120 5220
rect 176 5189 200 5245
rect -44 5148 200 5189
rect -44 5103 0 5148
rect 156 5103 200 5148
rect -44 5047 -22 5103
rect 34 5047 120 5096
rect 176 5047 200 5103
rect -44 5024 200 5047
rect -44 4972 0 5024
rect 156 4972 200 5024
rect -44 4961 200 4972
rect -44 4905 -22 4961
rect 34 4905 120 4961
rect 176 4905 200 4961
rect -44 4900 200 4905
rect -44 4848 0 4900
rect 156 4848 200 4900
rect -44 4819 200 4848
rect -44 4763 -22 4819
rect 34 4776 120 4819
rect 176 4763 200 4819
rect -44 4724 0 4763
rect 156 4724 200 4763
rect -44 4677 200 4724
rect -44 4621 -22 4677
rect 34 4652 120 4677
rect 176 4621 200 4677
rect -44 4600 0 4621
rect 156 4600 200 4621
rect -44 4535 200 4600
rect -44 4479 -22 4535
rect 34 4528 120 4535
rect 176 4479 200 4535
rect -44 4476 0 4479
rect 156 4476 200 4479
rect -44 4404 200 4476
rect -44 4393 0 4404
rect 156 4393 200 4404
rect -44 4337 -22 4393
rect 34 4337 120 4352
rect 176 4337 200 4393
rect -44 4280 200 4337
rect -44 4251 0 4280
rect 156 4251 200 4280
rect -44 4195 -22 4251
rect 34 4195 120 4228
rect 176 4195 200 4251
rect -44 4156 200 4195
rect -44 4109 0 4156
rect 156 4109 200 4156
rect -44 4053 -22 4109
rect 34 4053 120 4104
rect 176 4053 200 4109
rect -44 4032 200 4053
rect -44 3980 0 4032
rect 156 3980 200 4032
rect -44 3967 200 3980
rect -44 3911 -22 3967
rect 34 3911 120 3967
rect 176 3911 200 3967
rect -44 3908 200 3911
rect -44 3856 0 3908
rect 156 3856 200 3908
rect -44 3825 200 3856
rect -44 3769 -22 3825
rect 34 3784 120 3825
rect 176 3769 200 3825
rect -44 3732 0 3769
rect 156 3732 200 3769
rect -44 3683 200 3732
rect -44 3627 -22 3683
rect 34 3660 120 3683
rect 176 3627 200 3683
rect -44 3608 0 3627
rect 156 3608 200 3627
rect -44 3541 200 3608
rect -44 3485 -22 3541
rect 34 3536 120 3541
rect 176 3485 200 3541
rect -44 3484 0 3485
rect 156 3484 200 3485
rect -44 3412 200 3484
rect -44 3399 0 3412
rect 156 3399 200 3412
rect -44 3343 -22 3399
rect 34 3343 120 3360
rect 176 3343 200 3399
rect -44 3288 200 3343
rect -44 3236 0 3288
rect 156 3236 200 3288
rect -44 3164 200 3236
rect -44 3112 0 3164
rect 156 3112 200 3164
rect -44 3051 200 3112
rect -44 2995 -22 3051
rect 34 3040 120 3051
rect 176 2995 200 3051
rect -44 2988 0 2995
rect 156 2988 200 2995
rect -44 2916 200 2988
rect -44 2909 0 2916
rect 156 2909 200 2916
rect -44 2853 -22 2909
rect 34 2853 120 2864
rect 176 2853 200 2909
rect -44 2792 200 2853
rect -44 2767 0 2792
rect 156 2767 200 2792
rect -44 2711 -22 2767
rect 34 2711 120 2740
rect 176 2711 200 2767
rect -44 2668 200 2711
rect -44 2625 0 2668
rect 156 2625 200 2668
rect -44 2569 -22 2625
rect 34 2569 120 2616
rect 176 2569 200 2625
rect -44 2544 200 2569
rect -44 2492 0 2544
rect 156 2492 200 2544
rect -44 2483 200 2492
rect -44 2427 -22 2483
rect 34 2427 120 2483
rect 176 2427 200 2483
rect -44 2420 200 2427
rect -44 2368 0 2420
rect 156 2368 200 2420
rect -44 2341 200 2368
rect -44 2285 -22 2341
rect 34 2296 120 2341
rect 176 2285 200 2341
rect -44 2244 0 2285
rect 156 2244 200 2285
rect -44 2199 200 2244
rect -44 2143 -22 2199
rect 34 2172 120 2199
rect 176 2143 200 2199
rect -44 2120 0 2143
rect 156 2120 200 2143
rect -44 2057 200 2120
rect -44 2001 -22 2057
rect 34 2048 120 2057
rect 176 2001 200 2057
rect -44 1996 0 2001
rect 156 1996 200 2001
rect -44 1924 200 1996
rect -44 1915 0 1924
rect 156 1915 200 1924
rect -44 1859 -22 1915
rect 34 1859 120 1872
rect 176 1859 200 1915
rect -44 1800 200 1859
rect -44 1773 0 1800
rect 156 1773 200 1800
rect -44 1717 -22 1773
rect 34 1717 120 1748
rect 176 1717 200 1773
rect -44 1676 200 1717
rect -44 1631 0 1676
rect 156 1631 200 1676
rect -44 1575 -22 1631
rect 34 1575 120 1624
rect 176 1575 200 1631
rect -44 1552 200 1575
rect -44 1500 0 1552
rect 156 1500 200 1552
rect -44 1489 200 1500
rect -44 1433 -22 1489
rect 34 1433 120 1489
rect 176 1433 200 1489
rect -44 1428 200 1433
rect -44 1376 0 1428
rect 156 1376 200 1428
rect -44 1347 200 1376
rect -44 1291 -22 1347
rect 34 1304 120 1347
rect 176 1291 200 1347
rect -44 1252 0 1291
rect 156 1252 200 1291
rect -44 1205 200 1252
rect -44 1149 -22 1205
rect 34 1180 120 1205
rect 176 1149 200 1205
rect -44 1128 0 1149
rect 156 1128 200 1149
rect -44 1063 200 1128
rect -44 1007 -22 1063
rect 34 1056 120 1063
rect 176 1007 200 1063
rect -44 1004 0 1007
rect 156 1004 200 1007
rect -44 932 200 1004
rect -44 921 0 932
rect 156 921 200 932
rect -44 865 -22 921
rect 34 865 120 880
rect 176 865 200 921
rect -44 808 200 865
rect -44 779 0 808
rect 156 779 200 808
rect -44 723 -22 779
rect 34 723 120 756
rect 176 723 200 779
rect -44 684 200 723
rect -44 637 0 684
rect 156 637 200 684
rect -44 581 -22 637
rect 34 581 120 632
rect 176 581 200 637
rect -44 560 200 581
rect -44 508 0 560
rect 156 508 200 560
rect -44 495 200 508
rect -44 439 -22 495
rect 34 439 120 495
rect 176 439 200 495
rect -44 436 200 439
rect -44 384 0 436
rect 156 384 200 436
rect -44 353 200 384
rect -44 297 -22 353
rect 34 312 120 353
rect 176 297 200 353
rect -44 260 0 297
rect 156 260 200 297
rect -44 211 200 260
rect -44 155 -22 211
rect 34 188 120 211
rect 176 155 200 211
rect -44 136 0 155
rect 156 136 200 155
rect -44 64 200 136
rect -44 12 0 64
rect 156 12 200 64
rect -44 0 200 12
rect 340 11968 1584 12000
rect 340 11916 378 11968
rect 430 11916 502 11968
rect 554 11916 626 11968
rect 678 11916 750 11968
rect 802 11916 874 11968
rect 926 11916 998 11968
rect 1050 11916 1122 11968
rect 1174 11916 1246 11968
rect 1298 11916 1370 11968
rect 1422 11916 1494 11968
rect 1546 11916 1584 11968
rect 340 11844 1584 11916
rect 340 11792 378 11844
rect 430 11792 502 11844
rect 554 11792 626 11844
rect 678 11792 750 11844
rect 802 11792 874 11844
rect 926 11792 998 11844
rect 1050 11792 1122 11844
rect 1174 11792 1246 11844
rect 1298 11792 1370 11844
rect 1422 11792 1494 11844
rect 1546 11792 1584 11844
rect 340 11720 1584 11792
rect 340 11668 378 11720
rect 430 11668 502 11720
rect 554 11668 626 11720
rect 678 11668 750 11720
rect 802 11668 874 11720
rect 926 11668 998 11720
rect 1050 11668 1122 11720
rect 1174 11668 1246 11720
rect 1298 11668 1370 11720
rect 1422 11668 1494 11720
rect 1546 11668 1584 11720
rect 340 11596 1584 11668
rect 340 11544 378 11596
rect 430 11544 502 11596
rect 554 11544 626 11596
rect 678 11544 750 11596
rect 802 11544 874 11596
rect 926 11544 998 11596
rect 1050 11544 1122 11596
rect 1174 11544 1246 11596
rect 1298 11544 1370 11596
rect 1422 11544 1494 11596
rect 1546 11544 1584 11596
rect 340 11472 1584 11544
rect 340 11420 378 11472
rect 430 11420 502 11472
rect 554 11420 626 11472
rect 678 11420 750 11472
rect 802 11420 874 11472
rect 926 11420 998 11472
rect 1050 11420 1122 11472
rect 1174 11420 1246 11472
rect 1298 11420 1370 11472
rect 1422 11420 1494 11472
rect 1546 11420 1584 11472
rect 340 11348 1584 11420
rect 340 11296 378 11348
rect 430 11296 502 11348
rect 554 11296 626 11348
rect 678 11296 750 11348
rect 802 11296 874 11348
rect 926 11296 998 11348
rect 1050 11296 1122 11348
rect 1174 11296 1246 11348
rect 1298 11296 1370 11348
rect 1422 11296 1494 11348
rect 1546 11296 1584 11348
rect 340 11224 1584 11296
rect 340 11172 378 11224
rect 430 11172 502 11224
rect 554 11172 626 11224
rect 678 11172 750 11224
rect 802 11172 874 11224
rect 926 11172 998 11224
rect 1050 11172 1122 11224
rect 1174 11172 1246 11224
rect 1298 11172 1370 11224
rect 1422 11172 1494 11224
rect 1546 11172 1584 11224
rect 340 11100 1584 11172
rect 340 11048 378 11100
rect 430 11048 502 11100
rect 554 11048 626 11100
rect 678 11048 750 11100
rect 802 11048 874 11100
rect 926 11048 998 11100
rect 1050 11048 1122 11100
rect 1174 11048 1246 11100
rect 1298 11048 1370 11100
rect 1422 11048 1494 11100
rect 1546 11048 1584 11100
rect 340 10976 1584 11048
rect 340 10924 378 10976
rect 430 10924 502 10976
rect 554 10924 626 10976
rect 678 10924 750 10976
rect 802 10924 874 10976
rect 926 10924 998 10976
rect 1050 10924 1122 10976
rect 1174 10924 1246 10976
rect 1298 10924 1370 10976
rect 1422 10924 1494 10976
rect 1546 10924 1584 10976
rect 340 10852 1584 10924
rect 340 10800 378 10852
rect 430 10800 502 10852
rect 554 10800 626 10852
rect 678 10800 750 10852
rect 802 10800 874 10852
rect 926 10800 998 10852
rect 1050 10800 1122 10852
rect 1174 10800 1246 10852
rect 1298 10800 1370 10852
rect 1422 10800 1494 10852
rect 1546 10800 1584 10852
rect 340 10728 1584 10800
rect 340 10676 378 10728
rect 430 10676 502 10728
rect 554 10676 626 10728
rect 678 10676 750 10728
rect 802 10676 874 10728
rect 926 10676 998 10728
rect 1050 10676 1122 10728
rect 1174 10676 1246 10728
rect 1298 10676 1370 10728
rect 1422 10676 1494 10728
rect 1546 10676 1584 10728
rect 340 10604 1584 10676
rect 340 10552 378 10604
rect 430 10552 502 10604
rect 554 10552 626 10604
rect 678 10552 750 10604
rect 802 10552 874 10604
rect 926 10552 998 10604
rect 1050 10552 1122 10604
rect 1174 10552 1246 10604
rect 1298 10552 1370 10604
rect 1422 10552 1494 10604
rect 1546 10552 1584 10604
rect 340 10480 1584 10552
rect 340 10428 378 10480
rect 430 10428 502 10480
rect 554 10428 626 10480
rect 678 10428 750 10480
rect 802 10428 874 10480
rect 926 10428 998 10480
rect 1050 10428 1122 10480
rect 1174 10428 1246 10480
rect 1298 10428 1370 10480
rect 1422 10428 1494 10480
rect 1546 10428 1584 10480
rect 340 10356 1584 10428
rect 340 10304 378 10356
rect 430 10304 502 10356
rect 554 10304 626 10356
rect 678 10304 750 10356
rect 802 10304 874 10356
rect 926 10304 998 10356
rect 1050 10304 1122 10356
rect 1174 10304 1246 10356
rect 1298 10304 1370 10356
rect 1422 10304 1494 10356
rect 1546 10304 1584 10356
rect 340 10232 1584 10304
rect 340 10180 378 10232
rect 430 10180 502 10232
rect 554 10180 626 10232
rect 678 10180 750 10232
rect 802 10180 874 10232
rect 926 10180 998 10232
rect 1050 10180 1122 10232
rect 1174 10180 1246 10232
rect 1298 10180 1370 10232
rect 1422 10180 1494 10232
rect 1546 10180 1584 10232
rect 340 10108 1584 10180
rect 340 10056 378 10108
rect 430 10056 502 10108
rect 554 10056 626 10108
rect 678 10056 750 10108
rect 802 10056 874 10108
rect 926 10056 998 10108
rect 1050 10056 1122 10108
rect 1174 10056 1246 10108
rect 1298 10056 1370 10108
rect 1422 10056 1494 10108
rect 1546 10056 1584 10108
rect 340 9984 1584 10056
rect 340 9932 378 9984
rect 430 9932 502 9984
rect 554 9932 626 9984
rect 678 9932 750 9984
rect 802 9932 874 9984
rect 926 9932 998 9984
rect 1050 9932 1122 9984
rect 1174 9932 1246 9984
rect 1298 9932 1370 9984
rect 1422 9932 1494 9984
rect 1546 9932 1584 9984
rect 340 9860 1584 9932
rect 340 9808 378 9860
rect 430 9808 502 9860
rect 554 9808 626 9860
rect 678 9808 750 9860
rect 802 9808 874 9860
rect 926 9808 998 9860
rect 1050 9808 1122 9860
rect 1174 9808 1246 9860
rect 1298 9808 1370 9860
rect 1422 9808 1494 9860
rect 1546 9808 1584 9860
rect 340 9736 1584 9808
rect 340 9684 378 9736
rect 430 9684 502 9736
rect 554 9684 626 9736
rect 678 9684 750 9736
rect 802 9684 874 9736
rect 926 9684 998 9736
rect 1050 9684 1122 9736
rect 1174 9684 1246 9736
rect 1298 9684 1370 9736
rect 1422 9684 1494 9736
rect 1546 9684 1584 9736
rect 340 9612 1584 9684
rect 340 9560 378 9612
rect 430 9560 502 9612
rect 554 9560 626 9612
rect 678 9560 750 9612
rect 802 9560 874 9612
rect 926 9560 998 9612
rect 1050 9560 1122 9612
rect 1174 9560 1246 9612
rect 1298 9560 1370 9612
rect 1422 9560 1494 9612
rect 1546 9560 1584 9612
rect 340 9488 1584 9560
rect 340 9436 378 9488
rect 430 9436 502 9488
rect 554 9436 626 9488
rect 678 9436 750 9488
rect 802 9436 874 9488
rect 926 9436 998 9488
rect 1050 9436 1122 9488
rect 1174 9436 1246 9488
rect 1298 9436 1370 9488
rect 1422 9436 1494 9488
rect 1546 9436 1584 9488
rect 340 9364 1584 9436
rect 340 9312 378 9364
rect 430 9312 502 9364
rect 554 9312 626 9364
rect 678 9312 750 9364
rect 802 9312 874 9364
rect 926 9312 998 9364
rect 1050 9312 1122 9364
rect 1174 9312 1246 9364
rect 1298 9312 1370 9364
rect 1422 9312 1494 9364
rect 1546 9312 1584 9364
rect 340 9240 1584 9312
rect 340 9188 378 9240
rect 430 9188 502 9240
rect 554 9188 626 9240
rect 678 9188 750 9240
rect 802 9188 874 9240
rect 926 9188 998 9240
rect 1050 9188 1122 9240
rect 1174 9188 1246 9240
rect 1298 9188 1370 9240
rect 1422 9188 1494 9240
rect 1546 9188 1584 9240
rect 340 9116 1584 9188
rect 340 9064 378 9116
rect 430 9064 502 9116
rect 554 9064 626 9116
rect 678 9064 750 9116
rect 802 9064 874 9116
rect 926 9064 998 9116
rect 1050 9064 1122 9116
rect 1174 9064 1246 9116
rect 1298 9064 1370 9116
rect 1422 9064 1494 9116
rect 1546 9064 1584 9116
rect 340 8992 1584 9064
rect 340 8940 378 8992
rect 430 8940 502 8992
rect 554 8940 626 8992
rect 678 8940 750 8992
rect 802 8940 874 8992
rect 926 8940 998 8992
rect 1050 8940 1122 8992
rect 1174 8940 1246 8992
rect 1298 8940 1370 8992
rect 1422 8940 1494 8992
rect 1546 8940 1584 8992
rect 340 8868 1584 8940
rect 340 8816 378 8868
rect 430 8816 502 8868
rect 554 8816 626 8868
rect 678 8816 750 8868
rect 802 8816 874 8868
rect 926 8816 998 8868
rect 1050 8816 1122 8868
rect 1174 8816 1246 8868
rect 1298 8816 1370 8868
rect 1422 8816 1494 8868
rect 1546 8816 1584 8868
rect 340 8744 1584 8816
rect 340 8692 378 8744
rect 430 8692 502 8744
rect 554 8692 626 8744
rect 678 8692 750 8744
rect 802 8692 874 8744
rect 926 8692 998 8744
rect 1050 8692 1122 8744
rect 1174 8692 1246 8744
rect 1298 8692 1370 8744
rect 1422 8692 1494 8744
rect 1546 8692 1584 8744
rect 340 8620 1584 8692
rect 340 8568 378 8620
rect 430 8568 502 8620
rect 554 8568 626 8620
rect 678 8568 750 8620
rect 802 8568 874 8620
rect 926 8568 998 8620
rect 1050 8568 1122 8620
rect 1174 8568 1246 8620
rect 1298 8568 1370 8620
rect 1422 8568 1494 8620
rect 1546 8568 1584 8620
rect 340 8496 1584 8568
rect 340 8444 378 8496
rect 430 8444 502 8496
rect 554 8444 626 8496
rect 678 8444 750 8496
rect 802 8444 874 8496
rect 926 8444 998 8496
rect 1050 8444 1122 8496
rect 1174 8444 1246 8496
rect 1298 8444 1370 8496
rect 1422 8444 1494 8496
rect 1546 8444 1584 8496
rect 340 8372 1584 8444
rect 340 8320 378 8372
rect 430 8320 502 8372
rect 554 8320 626 8372
rect 678 8320 750 8372
rect 802 8320 874 8372
rect 926 8320 998 8372
rect 1050 8320 1122 8372
rect 1174 8320 1246 8372
rect 1298 8320 1370 8372
rect 1422 8320 1494 8372
rect 1546 8320 1584 8372
rect 340 8248 1584 8320
rect 340 8196 378 8248
rect 430 8196 502 8248
rect 554 8196 626 8248
rect 678 8196 750 8248
rect 802 8196 874 8248
rect 926 8196 998 8248
rect 1050 8196 1122 8248
rect 1174 8196 1246 8248
rect 1298 8196 1370 8248
rect 1422 8196 1494 8248
rect 1546 8196 1584 8248
rect 340 8124 1584 8196
rect 340 8072 378 8124
rect 430 8072 502 8124
rect 554 8072 626 8124
rect 678 8072 750 8124
rect 802 8072 874 8124
rect 926 8072 998 8124
rect 1050 8072 1122 8124
rect 1174 8072 1246 8124
rect 1298 8072 1370 8124
rect 1422 8072 1494 8124
rect 1546 8072 1584 8124
rect 340 8000 1584 8072
rect 340 7948 378 8000
rect 430 7948 502 8000
rect 554 7948 626 8000
rect 678 7948 750 8000
rect 802 7948 874 8000
rect 926 7948 998 8000
rect 1050 7948 1122 8000
rect 1174 7948 1246 8000
rect 1298 7948 1370 8000
rect 1422 7948 1494 8000
rect 1546 7948 1584 8000
rect 340 7876 1584 7948
rect 340 7824 378 7876
rect 430 7824 502 7876
rect 554 7824 626 7876
rect 678 7824 750 7876
rect 802 7824 874 7876
rect 926 7824 998 7876
rect 1050 7824 1122 7876
rect 1174 7824 1246 7876
rect 1298 7824 1370 7876
rect 1422 7824 1494 7876
rect 1546 7824 1584 7876
rect 340 7752 1584 7824
rect 340 7700 378 7752
rect 430 7700 502 7752
rect 554 7700 626 7752
rect 678 7700 750 7752
rect 802 7700 874 7752
rect 926 7700 998 7752
rect 1050 7700 1122 7752
rect 1174 7700 1246 7752
rect 1298 7700 1370 7752
rect 1422 7700 1494 7752
rect 1546 7700 1584 7752
rect 340 7628 1584 7700
rect 340 7576 378 7628
rect 430 7576 502 7628
rect 554 7576 626 7628
rect 678 7576 750 7628
rect 802 7576 874 7628
rect 926 7576 998 7628
rect 1050 7576 1122 7628
rect 1174 7576 1246 7628
rect 1298 7576 1370 7628
rect 1422 7576 1494 7628
rect 1546 7576 1584 7628
rect 340 7504 1584 7576
rect 340 7452 378 7504
rect 430 7452 502 7504
rect 554 7452 626 7504
rect 678 7452 750 7504
rect 802 7452 874 7504
rect 926 7452 998 7504
rect 1050 7452 1122 7504
rect 1174 7452 1246 7504
rect 1298 7452 1370 7504
rect 1422 7452 1494 7504
rect 1546 7452 1584 7504
rect 340 7380 1584 7452
rect 340 7328 378 7380
rect 430 7328 502 7380
rect 554 7328 626 7380
rect 678 7328 750 7380
rect 802 7328 874 7380
rect 926 7328 998 7380
rect 1050 7328 1122 7380
rect 1174 7328 1246 7380
rect 1298 7328 1370 7380
rect 1422 7328 1494 7380
rect 1546 7328 1584 7380
rect 340 7256 1584 7328
rect 340 7204 378 7256
rect 430 7204 502 7256
rect 554 7204 626 7256
rect 678 7204 750 7256
rect 802 7204 874 7256
rect 926 7204 998 7256
rect 1050 7204 1122 7256
rect 1174 7204 1246 7256
rect 1298 7204 1370 7256
rect 1422 7204 1494 7256
rect 1546 7204 1584 7256
rect 340 7132 1584 7204
rect 340 7080 378 7132
rect 430 7080 502 7132
rect 554 7080 626 7132
rect 678 7080 750 7132
rect 802 7080 874 7132
rect 926 7080 998 7132
rect 1050 7080 1122 7132
rect 1174 7080 1246 7132
rect 1298 7080 1370 7132
rect 1422 7080 1494 7132
rect 1546 7080 1584 7132
rect 340 7008 1584 7080
rect 340 6956 378 7008
rect 430 6956 502 7008
rect 554 6956 626 7008
rect 678 6956 750 7008
rect 802 6956 874 7008
rect 926 6956 998 7008
rect 1050 6956 1122 7008
rect 1174 6956 1246 7008
rect 1298 6956 1370 7008
rect 1422 6956 1494 7008
rect 1546 6956 1584 7008
rect 340 6884 1584 6956
rect 340 6832 378 6884
rect 430 6832 502 6884
rect 554 6832 626 6884
rect 678 6832 750 6884
rect 802 6832 874 6884
rect 926 6832 998 6884
rect 1050 6832 1122 6884
rect 1174 6832 1246 6884
rect 1298 6832 1370 6884
rect 1422 6832 1494 6884
rect 1546 6832 1584 6884
rect 340 6760 1584 6832
rect 340 6708 378 6760
rect 430 6708 502 6760
rect 554 6708 626 6760
rect 678 6708 750 6760
rect 802 6708 874 6760
rect 926 6708 998 6760
rect 1050 6708 1122 6760
rect 1174 6708 1246 6760
rect 1298 6708 1370 6760
rect 1422 6708 1494 6760
rect 1546 6708 1584 6760
rect 340 6636 1584 6708
rect 340 6584 378 6636
rect 430 6584 502 6636
rect 554 6584 626 6636
rect 678 6584 750 6636
rect 802 6584 874 6636
rect 926 6584 998 6636
rect 1050 6584 1122 6636
rect 1174 6584 1246 6636
rect 1298 6584 1370 6636
rect 1422 6584 1494 6636
rect 1546 6584 1584 6636
rect 340 6512 1584 6584
rect 340 6460 378 6512
rect 430 6460 502 6512
rect 554 6460 626 6512
rect 678 6460 750 6512
rect 802 6460 874 6512
rect 926 6460 998 6512
rect 1050 6460 1122 6512
rect 1174 6460 1246 6512
rect 1298 6460 1370 6512
rect 1422 6460 1494 6512
rect 1546 6460 1584 6512
rect 340 6388 1584 6460
rect 340 6336 378 6388
rect 430 6336 502 6388
rect 554 6336 626 6388
rect 678 6336 750 6388
rect 802 6336 874 6388
rect 926 6336 998 6388
rect 1050 6336 1122 6388
rect 1174 6336 1246 6388
rect 1298 6336 1370 6388
rect 1422 6336 1494 6388
rect 1546 6336 1584 6388
rect 340 6264 1584 6336
rect 340 6212 378 6264
rect 430 6212 502 6264
rect 554 6212 626 6264
rect 678 6212 750 6264
rect 802 6212 874 6264
rect 926 6212 998 6264
rect 1050 6212 1122 6264
rect 1174 6212 1246 6264
rect 1298 6212 1370 6264
rect 1422 6212 1494 6264
rect 1546 6212 1584 6264
rect 340 6140 1584 6212
rect 340 6088 378 6140
rect 430 6088 502 6140
rect 554 6088 626 6140
rect 678 6088 750 6140
rect 802 6088 874 6140
rect 926 6088 998 6140
rect 1050 6088 1122 6140
rect 1174 6088 1246 6140
rect 1298 6088 1370 6140
rect 1422 6088 1494 6140
rect 1546 6088 1584 6140
rect 340 6016 1584 6088
rect 340 5964 378 6016
rect 430 5964 502 6016
rect 554 5964 626 6016
rect 678 5964 750 6016
rect 802 5964 874 6016
rect 926 5964 998 6016
rect 1050 5964 1122 6016
rect 1174 5964 1246 6016
rect 1298 5964 1370 6016
rect 1422 5964 1494 6016
rect 1546 5964 1584 6016
rect 340 5892 1584 5964
rect 340 5840 378 5892
rect 430 5840 502 5892
rect 554 5840 626 5892
rect 678 5840 750 5892
rect 802 5840 874 5892
rect 926 5840 998 5892
rect 1050 5840 1122 5892
rect 1174 5840 1246 5892
rect 1298 5840 1370 5892
rect 1422 5840 1494 5892
rect 1546 5840 1584 5892
rect 340 5768 1584 5840
rect 340 5716 378 5768
rect 430 5716 502 5768
rect 554 5716 626 5768
rect 678 5716 750 5768
rect 802 5716 874 5768
rect 926 5716 998 5768
rect 1050 5716 1122 5768
rect 1174 5716 1246 5768
rect 1298 5716 1370 5768
rect 1422 5716 1494 5768
rect 1546 5716 1584 5768
rect 340 5644 1584 5716
rect 340 5592 378 5644
rect 430 5592 502 5644
rect 554 5592 626 5644
rect 678 5592 750 5644
rect 802 5592 874 5644
rect 926 5592 998 5644
rect 1050 5592 1122 5644
rect 1174 5592 1246 5644
rect 1298 5592 1370 5644
rect 1422 5592 1494 5644
rect 1546 5592 1584 5644
rect 340 5520 1584 5592
rect 340 5468 378 5520
rect 430 5468 502 5520
rect 554 5468 626 5520
rect 678 5468 750 5520
rect 802 5468 874 5520
rect 926 5468 998 5520
rect 1050 5468 1122 5520
rect 1174 5468 1246 5520
rect 1298 5468 1370 5520
rect 1422 5468 1494 5520
rect 1546 5468 1584 5520
rect 340 5396 1584 5468
rect 340 5344 378 5396
rect 430 5344 502 5396
rect 554 5344 626 5396
rect 678 5344 750 5396
rect 802 5344 874 5396
rect 926 5344 998 5396
rect 1050 5344 1122 5396
rect 1174 5344 1246 5396
rect 1298 5344 1370 5396
rect 1422 5344 1494 5396
rect 1546 5344 1584 5396
rect 340 5272 1584 5344
rect 340 5220 378 5272
rect 430 5220 502 5272
rect 554 5220 626 5272
rect 678 5220 750 5272
rect 802 5220 874 5272
rect 926 5220 998 5272
rect 1050 5220 1122 5272
rect 1174 5220 1246 5272
rect 1298 5220 1370 5272
rect 1422 5220 1494 5272
rect 1546 5220 1584 5272
rect 340 5148 1584 5220
rect 340 5096 378 5148
rect 430 5096 502 5148
rect 554 5096 626 5148
rect 678 5096 750 5148
rect 802 5096 874 5148
rect 926 5096 998 5148
rect 1050 5096 1122 5148
rect 1174 5096 1246 5148
rect 1298 5096 1370 5148
rect 1422 5096 1494 5148
rect 1546 5096 1584 5148
rect 340 5024 1584 5096
rect 340 4972 378 5024
rect 430 4972 502 5024
rect 554 4972 626 5024
rect 678 4972 750 5024
rect 802 4972 874 5024
rect 926 4972 998 5024
rect 1050 4972 1122 5024
rect 1174 4972 1246 5024
rect 1298 4972 1370 5024
rect 1422 4972 1494 5024
rect 1546 4972 1584 5024
rect 340 4900 1584 4972
rect 340 4848 378 4900
rect 430 4848 502 4900
rect 554 4848 626 4900
rect 678 4848 750 4900
rect 802 4848 874 4900
rect 926 4848 998 4900
rect 1050 4848 1122 4900
rect 1174 4848 1246 4900
rect 1298 4848 1370 4900
rect 1422 4848 1494 4900
rect 1546 4848 1584 4900
rect 340 4776 1584 4848
rect 340 4724 378 4776
rect 430 4724 502 4776
rect 554 4724 626 4776
rect 678 4724 750 4776
rect 802 4724 874 4776
rect 926 4724 998 4776
rect 1050 4724 1122 4776
rect 1174 4724 1246 4776
rect 1298 4724 1370 4776
rect 1422 4724 1494 4776
rect 1546 4724 1584 4776
rect 340 4652 1584 4724
rect 340 4600 378 4652
rect 430 4600 502 4652
rect 554 4600 626 4652
rect 678 4600 750 4652
rect 802 4600 874 4652
rect 926 4600 998 4652
rect 1050 4600 1122 4652
rect 1174 4600 1246 4652
rect 1298 4600 1370 4652
rect 1422 4600 1494 4652
rect 1546 4600 1584 4652
rect 340 4528 1584 4600
rect 340 4476 378 4528
rect 430 4476 502 4528
rect 554 4476 626 4528
rect 678 4476 750 4528
rect 802 4476 874 4528
rect 926 4476 998 4528
rect 1050 4476 1122 4528
rect 1174 4476 1246 4528
rect 1298 4476 1370 4528
rect 1422 4476 1494 4528
rect 1546 4476 1584 4528
rect 340 4404 1584 4476
rect 340 4352 378 4404
rect 430 4352 502 4404
rect 554 4352 626 4404
rect 678 4352 750 4404
rect 802 4352 874 4404
rect 926 4352 998 4404
rect 1050 4352 1122 4404
rect 1174 4352 1246 4404
rect 1298 4352 1370 4404
rect 1422 4352 1494 4404
rect 1546 4352 1584 4404
rect 340 4280 1584 4352
rect 340 4228 378 4280
rect 430 4228 502 4280
rect 554 4228 626 4280
rect 678 4228 750 4280
rect 802 4228 874 4280
rect 926 4228 998 4280
rect 1050 4228 1122 4280
rect 1174 4228 1246 4280
rect 1298 4228 1370 4280
rect 1422 4228 1494 4280
rect 1546 4228 1584 4280
rect 340 4156 1584 4228
rect 340 4104 378 4156
rect 430 4104 502 4156
rect 554 4104 626 4156
rect 678 4104 750 4156
rect 802 4104 874 4156
rect 926 4104 998 4156
rect 1050 4104 1122 4156
rect 1174 4104 1246 4156
rect 1298 4104 1370 4156
rect 1422 4104 1494 4156
rect 1546 4104 1584 4156
rect 340 4032 1584 4104
rect 340 3980 378 4032
rect 430 3980 502 4032
rect 554 3980 626 4032
rect 678 3980 750 4032
rect 802 3980 874 4032
rect 926 3980 998 4032
rect 1050 3980 1122 4032
rect 1174 3980 1246 4032
rect 1298 3980 1370 4032
rect 1422 3980 1494 4032
rect 1546 3980 1584 4032
rect 340 3908 1584 3980
rect 340 3856 378 3908
rect 430 3856 502 3908
rect 554 3856 626 3908
rect 678 3856 750 3908
rect 802 3856 874 3908
rect 926 3856 998 3908
rect 1050 3856 1122 3908
rect 1174 3856 1246 3908
rect 1298 3856 1370 3908
rect 1422 3856 1494 3908
rect 1546 3856 1584 3908
rect 340 3784 1584 3856
rect 340 3732 378 3784
rect 430 3732 502 3784
rect 554 3732 626 3784
rect 678 3732 750 3784
rect 802 3732 874 3784
rect 926 3732 998 3784
rect 1050 3732 1122 3784
rect 1174 3732 1246 3784
rect 1298 3732 1370 3784
rect 1422 3732 1494 3784
rect 1546 3732 1584 3784
rect 340 3660 1584 3732
rect 340 3608 378 3660
rect 430 3608 502 3660
rect 554 3608 626 3660
rect 678 3608 750 3660
rect 802 3608 874 3660
rect 926 3608 998 3660
rect 1050 3608 1122 3660
rect 1174 3608 1246 3660
rect 1298 3608 1370 3660
rect 1422 3608 1494 3660
rect 1546 3608 1584 3660
rect 340 3536 1584 3608
rect 340 3484 378 3536
rect 430 3484 502 3536
rect 554 3484 626 3536
rect 678 3484 750 3536
rect 802 3484 874 3536
rect 926 3484 998 3536
rect 1050 3484 1122 3536
rect 1174 3484 1246 3536
rect 1298 3484 1370 3536
rect 1422 3484 1494 3536
rect 1546 3484 1584 3536
rect 340 3412 1584 3484
rect 340 3360 378 3412
rect 430 3360 502 3412
rect 554 3360 626 3412
rect 678 3360 750 3412
rect 802 3360 874 3412
rect 926 3360 998 3412
rect 1050 3360 1122 3412
rect 1174 3360 1246 3412
rect 1298 3360 1370 3412
rect 1422 3360 1494 3412
rect 1546 3360 1584 3412
rect 340 3288 1584 3360
rect 340 3236 378 3288
rect 430 3236 502 3288
rect 554 3236 626 3288
rect 678 3236 750 3288
rect 802 3236 874 3288
rect 926 3236 998 3288
rect 1050 3236 1122 3288
rect 1174 3236 1246 3288
rect 1298 3236 1370 3288
rect 1422 3236 1494 3288
rect 1546 3236 1584 3288
rect 340 3164 1584 3236
rect 340 3112 378 3164
rect 430 3112 502 3164
rect 554 3112 626 3164
rect 678 3112 750 3164
rect 802 3112 874 3164
rect 926 3112 998 3164
rect 1050 3112 1122 3164
rect 1174 3112 1246 3164
rect 1298 3112 1370 3164
rect 1422 3112 1494 3164
rect 1546 3112 1584 3164
rect 340 3040 1584 3112
rect 340 2988 378 3040
rect 430 2988 502 3040
rect 554 2988 626 3040
rect 678 2988 750 3040
rect 802 2988 874 3040
rect 926 2988 998 3040
rect 1050 2988 1122 3040
rect 1174 2988 1246 3040
rect 1298 2988 1370 3040
rect 1422 2988 1494 3040
rect 1546 2988 1584 3040
rect 340 2916 1584 2988
rect 340 2864 378 2916
rect 430 2864 502 2916
rect 554 2864 626 2916
rect 678 2864 750 2916
rect 802 2864 874 2916
rect 926 2864 998 2916
rect 1050 2864 1122 2916
rect 1174 2864 1246 2916
rect 1298 2864 1370 2916
rect 1422 2864 1494 2916
rect 1546 2864 1584 2916
rect 340 2792 1584 2864
rect 340 2740 378 2792
rect 430 2740 502 2792
rect 554 2740 626 2792
rect 678 2740 750 2792
rect 802 2740 874 2792
rect 926 2740 998 2792
rect 1050 2740 1122 2792
rect 1174 2740 1246 2792
rect 1298 2740 1370 2792
rect 1422 2740 1494 2792
rect 1546 2740 1584 2792
rect 340 2668 1584 2740
rect 340 2616 378 2668
rect 430 2616 502 2668
rect 554 2616 626 2668
rect 678 2616 750 2668
rect 802 2616 874 2668
rect 926 2616 998 2668
rect 1050 2616 1122 2668
rect 1174 2616 1246 2668
rect 1298 2616 1370 2668
rect 1422 2616 1494 2668
rect 1546 2616 1584 2668
rect 340 2544 1584 2616
rect 340 2492 378 2544
rect 430 2492 502 2544
rect 554 2492 626 2544
rect 678 2492 750 2544
rect 802 2492 874 2544
rect 926 2492 998 2544
rect 1050 2492 1122 2544
rect 1174 2492 1246 2544
rect 1298 2492 1370 2544
rect 1422 2492 1494 2544
rect 1546 2492 1584 2544
rect 340 2420 1584 2492
rect 340 2368 378 2420
rect 430 2368 502 2420
rect 554 2368 626 2420
rect 678 2368 750 2420
rect 802 2368 874 2420
rect 926 2368 998 2420
rect 1050 2368 1122 2420
rect 1174 2368 1246 2420
rect 1298 2368 1370 2420
rect 1422 2368 1494 2420
rect 1546 2368 1584 2420
rect 340 2296 1584 2368
rect 340 2244 378 2296
rect 430 2244 502 2296
rect 554 2244 626 2296
rect 678 2244 750 2296
rect 802 2244 874 2296
rect 926 2244 998 2296
rect 1050 2244 1122 2296
rect 1174 2244 1246 2296
rect 1298 2244 1370 2296
rect 1422 2244 1494 2296
rect 1546 2244 1584 2296
rect 340 2172 1584 2244
rect 340 2120 378 2172
rect 430 2120 502 2172
rect 554 2120 626 2172
rect 678 2120 750 2172
rect 802 2120 874 2172
rect 926 2120 998 2172
rect 1050 2120 1122 2172
rect 1174 2120 1246 2172
rect 1298 2120 1370 2172
rect 1422 2120 1494 2172
rect 1546 2120 1584 2172
rect 340 2048 1584 2120
rect 340 1996 378 2048
rect 430 1996 502 2048
rect 554 1996 626 2048
rect 678 1996 750 2048
rect 802 1996 874 2048
rect 926 1996 998 2048
rect 1050 1996 1122 2048
rect 1174 1996 1246 2048
rect 1298 1996 1370 2048
rect 1422 1996 1494 2048
rect 1546 1996 1584 2048
rect 340 1924 1584 1996
rect 340 1872 378 1924
rect 430 1872 502 1924
rect 554 1872 626 1924
rect 678 1872 750 1924
rect 802 1872 874 1924
rect 926 1872 998 1924
rect 1050 1872 1122 1924
rect 1174 1872 1246 1924
rect 1298 1872 1370 1924
rect 1422 1872 1494 1924
rect 1546 1872 1584 1924
rect 340 1800 1584 1872
rect 340 1748 378 1800
rect 430 1748 502 1800
rect 554 1748 626 1800
rect 678 1748 750 1800
rect 802 1748 874 1800
rect 926 1748 998 1800
rect 1050 1748 1122 1800
rect 1174 1748 1246 1800
rect 1298 1748 1370 1800
rect 1422 1748 1494 1800
rect 1546 1748 1584 1800
rect 340 1676 1584 1748
rect 340 1624 378 1676
rect 430 1624 502 1676
rect 554 1624 626 1676
rect 678 1624 750 1676
rect 802 1624 874 1676
rect 926 1624 998 1676
rect 1050 1624 1122 1676
rect 1174 1624 1246 1676
rect 1298 1624 1370 1676
rect 1422 1624 1494 1676
rect 1546 1624 1584 1676
rect 340 1552 1584 1624
rect 340 1500 378 1552
rect 430 1500 502 1552
rect 554 1500 626 1552
rect 678 1500 750 1552
rect 802 1500 874 1552
rect 926 1500 998 1552
rect 1050 1500 1122 1552
rect 1174 1500 1246 1552
rect 1298 1500 1370 1552
rect 1422 1500 1494 1552
rect 1546 1500 1584 1552
rect 340 1428 1584 1500
rect 340 1376 378 1428
rect 430 1376 502 1428
rect 554 1376 626 1428
rect 678 1376 750 1428
rect 802 1376 874 1428
rect 926 1376 998 1428
rect 1050 1376 1122 1428
rect 1174 1376 1246 1428
rect 1298 1376 1370 1428
rect 1422 1376 1494 1428
rect 1546 1376 1584 1428
rect 340 1304 1584 1376
rect 340 1252 378 1304
rect 430 1252 502 1304
rect 554 1252 626 1304
rect 678 1252 750 1304
rect 802 1252 874 1304
rect 926 1252 998 1304
rect 1050 1252 1122 1304
rect 1174 1252 1246 1304
rect 1298 1252 1370 1304
rect 1422 1252 1494 1304
rect 1546 1252 1584 1304
rect 340 1180 1584 1252
rect 340 1128 378 1180
rect 430 1128 502 1180
rect 554 1128 626 1180
rect 678 1128 750 1180
rect 802 1128 874 1180
rect 926 1128 998 1180
rect 1050 1128 1122 1180
rect 1174 1128 1246 1180
rect 1298 1128 1370 1180
rect 1422 1128 1494 1180
rect 1546 1128 1584 1180
rect 340 1056 1584 1128
rect 340 1004 378 1056
rect 430 1004 502 1056
rect 554 1004 626 1056
rect 678 1004 750 1056
rect 802 1004 874 1056
rect 926 1004 998 1056
rect 1050 1004 1122 1056
rect 1174 1004 1246 1056
rect 1298 1004 1370 1056
rect 1422 1004 1494 1056
rect 1546 1004 1584 1056
rect 340 932 1584 1004
rect 340 880 378 932
rect 430 880 502 932
rect 554 880 626 932
rect 678 880 750 932
rect 802 880 874 932
rect 926 880 998 932
rect 1050 880 1122 932
rect 1174 880 1246 932
rect 1298 880 1370 932
rect 1422 880 1494 932
rect 1546 880 1584 932
rect 340 808 1584 880
rect 340 756 378 808
rect 430 756 502 808
rect 554 756 626 808
rect 678 756 750 808
rect 802 756 874 808
rect 926 756 998 808
rect 1050 756 1122 808
rect 1174 756 1246 808
rect 1298 756 1370 808
rect 1422 756 1494 808
rect 1546 756 1584 808
rect 340 684 1584 756
rect 340 632 378 684
rect 430 632 502 684
rect 554 632 626 684
rect 678 632 750 684
rect 802 632 874 684
rect 926 632 998 684
rect 1050 632 1122 684
rect 1174 632 1246 684
rect 1298 632 1370 684
rect 1422 632 1494 684
rect 1546 632 1584 684
rect 340 560 1584 632
rect 340 508 378 560
rect 430 508 502 560
rect 554 508 626 560
rect 678 508 750 560
rect 802 508 874 560
rect 926 508 998 560
rect 1050 508 1122 560
rect 1174 508 1246 560
rect 1298 508 1370 560
rect 1422 508 1494 560
rect 1546 508 1584 560
rect 340 436 1584 508
rect 340 384 378 436
rect 430 384 502 436
rect 554 384 626 436
rect 678 384 750 436
rect 802 384 874 436
rect 926 384 998 436
rect 1050 384 1122 436
rect 1174 384 1246 436
rect 1298 384 1370 436
rect 1422 384 1494 436
rect 1546 384 1584 436
rect 340 312 1584 384
rect 340 260 378 312
rect 430 260 502 312
rect 554 260 626 312
rect 678 260 750 312
rect 802 260 874 312
rect 926 260 998 312
rect 1050 260 1122 312
rect 1174 260 1246 312
rect 1298 260 1370 312
rect 1422 260 1494 312
rect 1546 260 1584 312
rect 340 188 1584 260
rect 340 136 378 188
rect 430 136 502 188
rect 554 136 626 188
rect 678 136 750 188
rect 802 136 874 188
rect 926 136 998 188
rect 1050 136 1122 188
rect 1174 136 1246 188
rect 1298 136 1370 188
rect 1422 136 1494 188
rect 1546 136 1584 188
rect 340 64 1584 136
rect 340 12 378 64
rect 430 12 502 64
rect 554 12 626 64
rect 678 12 750 64
rect 802 12 874 64
rect 926 12 998 64
rect 1050 12 1122 64
rect 1174 12 1246 64
rect 1298 12 1370 64
rect 1422 12 1494 64
rect 1546 12 1584 64
rect 340 0 1584 12
<< via2 >>
rect -22 11916 0 11938
rect 0 11916 34 11938
rect 120 11916 156 11938
rect 156 11916 176 11938
rect -22 11882 34 11916
rect 120 11882 176 11916
rect -22 11792 0 11796
rect 0 11792 34 11796
rect 120 11792 156 11796
rect 156 11792 176 11796
rect -22 11740 34 11792
rect 120 11740 176 11792
rect -22 11598 34 11654
rect 120 11598 176 11654
rect -22 11472 34 11512
rect 120 11472 176 11512
rect -22 11456 0 11472
rect 0 11456 34 11472
rect 120 11456 156 11472
rect 156 11456 176 11472
rect -22 11348 34 11370
rect 120 11348 176 11370
rect -22 11314 0 11348
rect 0 11314 34 11348
rect 120 11314 156 11348
rect 156 11314 176 11348
rect -22 11224 34 11228
rect 120 11224 176 11228
rect -22 11172 0 11224
rect 0 11172 34 11224
rect 120 11172 156 11224
rect 156 11172 176 11224
rect -22 11048 0 11086
rect 0 11048 34 11086
rect 120 11048 156 11086
rect 156 11048 176 11086
rect -22 11030 34 11048
rect 120 11030 176 11048
rect -22 10924 0 10944
rect 0 10924 34 10944
rect 120 10924 156 10944
rect 156 10924 176 10944
rect -22 10888 34 10924
rect 120 10888 176 10924
rect -22 10800 0 10802
rect 0 10800 34 10802
rect 120 10800 156 10802
rect 156 10800 176 10802
rect -22 10746 34 10800
rect 120 10746 176 10800
rect -22 10604 34 10660
rect 120 10604 176 10660
rect -22 10480 34 10518
rect 120 10480 176 10518
rect -22 10462 0 10480
rect 0 10462 34 10480
rect 120 10462 156 10480
rect 156 10462 176 10480
rect -22 10356 34 10376
rect 120 10356 176 10376
rect -22 10320 0 10356
rect 0 10320 34 10356
rect 120 10320 156 10356
rect 156 10320 176 10356
rect -22 10232 34 10234
rect 120 10232 176 10234
rect -22 10180 0 10232
rect 0 10180 34 10232
rect 120 10180 156 10232
rect 156 10180 176 10232
rect -22 10178 34 10180
rect 120 10178 176 10180
rect -22 10056 0 10092
rect 0 10056 34 10092
rect 120 10056 156 10092
rect 156 10056 176 10092
rect -22 10036 34 10056
rect 120 10036 176 10056
rect -22 9932 0 9950
rect 0 9932 34 9950
rect 120 9932 156 9950
rect 156 9932 176 9950
rect -22 9894 34 9932
rect 120 9894 176 9932
rect -22 9752 34 9808
rect 120 9752 176 9808
rect -22 9370 34 9426
rect 120 9370 176 9426
rect -22 9240 34 9284
rect 120 9240 176 9284
rect -22 9228 0 9240
rect 0 9228 34 9240
rect 120 9228 156 9240
rect 156 9228 176 9240
rect -22 9116 34 9142
rect 120 9116 176 9142
rect -22 9086 0 9116
rect 0 9086 34 9116
rect 120 9086 156 9116
rect 156 9086 176 9116
rect -22 8992 34 9000
rect 120 8992 176 9000
rect -22 8944 0 8992
rect 0 8944 34 8992
rect 120 8944 156 8992
rect 156 8944 176 8992
rect -22 8816 0 8858
rect 0 8816 34 8858
rect 120 8816 156 8858
rect 156 8816 176 8858
rect -22 8802 34 8816
rect 120 8802 176 8816
rect -22 8692 0 8716
rect 0 8692 34 8716
rect 120 8692 156 8716
rect 156 8692 176 8716
rect -22 8660 34 8692
rect 120 8660 176 8692
rect -22 8568 0 8574
rect 0 8568 34 8574
rect 120 8568 156 8574
rect 156 8568 176 8574
rect -22 8518 34 8568
rect 120 8518 176 8568
rect -22 8376 34 8432
rect 120 8376 176 8432
rect -22 8248 34 8290
rect 120 8248 176 8290
rect -22 8234 0 8248
rect 0 8234 34 8248
rect 120 8234 156 8248
rect 156 8234 176 8248
rect -22 8124 34 8148
rect 120 8124 176 8148
rect -22 8092 0 8124
rect 0 8092 34 8124
rect 120 8092 156 8124
rect 156 8092 176 8124
rect -22 8000 34 8006
rect 120 8000 176 8006
rect -22 7950 0 8000
rect 0 7950 34 8000
rect 120 7950 156 8000
rect 156 7950 176 8000
rect -22 7824 0 7864
rect 0 7824 34 7864
rect 120 7824 156 7864
rect 156 7824 176 7864
rect -22 7808 34 7824
rect 120 7808 176 7824
rect -22 7700 0 7722
rect 0 7700 34 7722
rect 120 7700 156 7722
rect 156 7700 176 7722
rect -22 7666 34 7700
rect 120 7666 176 7700
rect -22 7576 0 7580
rect 0 7576 34 7580
rect 120 7576 156 7580
rect 156 7576 176 7580
rect -22 7524 34 7576
rect 120 7524 176 7576
rect -22 7382 34 7438
rect 120 7382 176 7438
rect -22 7256 34 7296
rect 120 7256 176 7296
rect -22 7240 0 7256
rect 0 7240 34 7256
rect 120 7240 156 7256
rect 156 7240 176 7256
rect -22 7132 34 7154
rect 120 7132 176 7154
rect -22 7098 0 7132
rect 0 7098 34 7132
rect 120 7098 156 7132
rect 156 7098 176 7132
rect -22 7008 34 7012
rect 120 7008 176 7012
rect -22 6956 0 7008
rect 0 6956 34 7008
rect 120 6956 156 7008
rect 156 6956 176 7008
rect -22 6832 0 6870
rect 0 6832 34 6870
rect 120 6832 156 6870
rect 156 6832 176 6870
rect -22 6814 34 6832
rect 120 6814 176 6832
rect -22 6708 0 6728
rect 0 6708 34 6728
rect 120 6708 156 6728
rect 156 6708 176 6728
rect -22 6672 34 6708
rect 120 6672 176 6708
rect -22 6584 0 6586
rect 0 6584 34 6586
rect 120 6584 156 6586
rect 156 6584 176 6586
rect -22 6530 34 6584
rect 120 6530 176 6584
rect -22 6212 0 6239
rect 0 6212 34 6239
rect 120 6212 156 6239
rect 156 6212 176 6239
rect -22 6183 34 6212
rect 120 6183 176 6212
rect -22 6088 0 6097
rect 0 6088 34 6097
rect 120 6088 156 6097
rect 156 6088 176 6097
rect -22 6041 34 6088
rect 120 6041 176 6088
rect -22 5899 34 5955
rect 120 5899 176 5955
rect -22 5768 34 5813
rect 120 5768 176 5813
rect -22 5757 0 5768
rect 0 5757 34 5768
rect 120 5757 156 5768
rect 156 5757 176 5768
rect -22 5644 34 5671
rect 120 5644 176 5671
rect -22 5615 0 5644
rect 0 5615 34 5644
rect 120 5615 156 5644
rect 156 5615 176 5644
rect -22 5520 34 5529
rect 120 5520 176 5529
rect -22 5473 0 5520
rect 0 5473 34 5520
rect 120 5473 156 5520
rect 156 5473 176 5520
rect -22 5344 0 5387
rect 0 5344 34 5387
rect 120 5344 156 5387
rect 156 5344 176 5387
rect -22 5331 34 5344
rect 120 5331 176 5344
rect -22 5220 0 5245
rect 0 5220 34 5245
rect 120 5220 156 5245
rect 156 5220 176 5245
rect -22 5189 34 5220
rect 120 5189 176 5220
rect -22 5096 0 5103
rect 0 5096 34 5103
rect 120 5096 156 5103
rect 156 5096 176 5103
rect -22 5047 34 5096
rect 120 5047 176 5096
rect -22 4905 34 4961
rect 120 4905 176 4961
rect -22 4776 34 4819
rect 120 4776 176 4819
rect -22 4763 0 4776
rect 0 4763 34 4776
rect 120 4763 156 4776
rect 156 4763 176 4776
rect -22 4652 34 4677
rect 120 4652 176 4677
rect -22 4621 0 4652
rect 0 4621 34 4652
rect 120 4621 156 4652
rect 156 4621 176 4652
rect -22 4528 34 4535
rect 120 4528 176 4535
rect -22 4479 0 4528
rect 0 4479 34 4528
rect 120 4479 156 4528
rect 156 4479 176 4528
rect -22 4352 0 4393
rect 0 4352 34 4393
rect 120 4352 156 4393
rect 156 4352 176 4393
rect -22 4337 34 4352
rect 120 4337 176 4352
rect -22 4228 0 4251
rect 0 4228 34 4251
rect 120 4228 156 4251
rect 156 4228 176 4251
rect -22 4195 34 4228
rect 120 4195 176 4228
rect -22 4104 0 4109
rect 0 4104 34 4109
rect 120 4104 156 4109
rect 156 4104 176 4109
rect -22 4053 34 4104
rect 120 4053 176 4104
rect -22 3911 34 3967
rect 120 3911 176 3967
rect -22 3784 34 3825
rect 120 3784 176 3825
rect -22 3769 0 3784
rect 0 3769 34 3784
rect 120 3769 156 3784
rect 156 3769 176 3784
rect -22 3660 34 3683
rect 120 3660 176 3683
rect -22 3627 0 3660
rect 0 3627 34 3660
rect 120 3627 156 3660
rect 156 3627 176 3660
rect -22 3536 34 3541
rect 120 3536 176 3541
rect -22 3485 0 3536
rect 0 3485 34 3536
rect 120 3485 156 3536
rect 156 3485 176 3536
rect -22 3360 0 3399
rect 0 3360 34 3399
rect 120 3360 156 3399
rect 156 3360 176 3399
rect -22 3343 34 3360
rect 120 3343 176 3360
rect -22 3040 34 3051
rect 120 3040 176 3051
rect -22 2995 0 3040
rect 0 2995 34 3040
rect 120 2995 156 3040
rect 156 2995 176 3040
rect -22 2864 0 2909
rect 0 2864 34 2909
rect 120 2864 156 2909
rect 156 2864 176 2909
rect -22 2853 34 2864
rect 120 2853 176 2864
rect -22 2740 0 2767
rect 0 2740 34 2767
rect 120 2740 156 2767
rect 156 2740 176 2767
rect -22 2711 34 2740
rect 120 2711 176 2740
rect -22 2616 0 2625
rect 0 2616 34 2625
rect 120 2616 156 2625
rect 156 2616 176 2625
rect -22 2569 34 2616
rect 120 2569 176 2616
rect -22 2427 34 2483
rect 120 2427 176 2483
rect -22 2296 34 2341
rect 120 2296 176 2341
rect -22 2285 0 2296
rect 0 2285 34 2296
rect 120 2285 156 2296
rect 156 2285 176 2296
rect -22 2172 34 2199
rect 120 2172 176 2199
rect -22 2143 0 2172
rect 0 2143 34 2172
rect 120 2143 156 2172
rect 156 2143 176 2172
rect -22 2048 34 2057
rect 120 2048 176 2057
rect -22 2001 0 2048
rect 0 2001 34 2048
rect 120 2001 156 2048
rect 156 2001 176 2048
rect -22 1872 0 1915
rect 0 1872 34 1915
rect 120 1872 156 1915
rect 156 1872 176 1915
rect -22 1859 34 1872
rect 120 1859 176 1872
rect -22 1748 0 1773
rect 0 1748 34 1773
rect 120 1748 156 1773
rect 156 1748 176 1773
rect -22 1717 34 1748
rect 120 1717 176 1748
rect -22 1624 0 1631
rect 0 1624 34 1631
rect 120 1624 156 1631
rect 156 1624 176 1631
rect -22 1575 34 1624
rect 120 1575 176 1624
rect -22 1433 34 1489
rect 120 1433 176 1489
rect -22 1304 34 1347
rect 120 1304 176 1347
rect -22 1291 0 1304
rect 0 1291 34 1304
rect 120 1291 156 1304
rect 156 1291 176 1304
rect -22 1180 34 1205
rect 120 1180 176 1205
rect -22 1149 0 1180
rect 0 1149 34 1180
rect 120 1149 156 1180
rect 156 1149 176 1180
rect -22 1056 34 1063
rect 120 1056 176 1063
rect -22 1007 0 1056
rect 0 1007 34 1056
rect 120 1007 156 1056
rect 156 1007 176 1056
rect -22 880 0 921
rect 0 880 34 921
rect 120 880 156 921
rect 156 880 176 921
rect -22 865 34 880
rect 120 865 176 880
rect -22 756 0 779
rect 0 756 34 779
rect 120 756 156 779
rect 156 756 176 779
rect -22 723 34 756
rect 120 723 176 756
rect -22 632 0 637
rect 0 632 34 637
rect 120 632 156 637
rect 156 632 176 637
rect -22 581 34 632
rect 120 581 176 632
rect -22 439 34 495
rect 120 439 176 495
rect -22 312 34 353
rect 120 312 176 353
rect -22 297 0 312
rect 0 297 34 312
rect 120 297 156 312
rect 156 297 176 312
rect -22 188 34 211
rect 120 188 176 211
rect -22 155 0 188
rect 0 155 34 188
rect 120 155 156 188
rect 156 155 176 188
<< metal3 >>
rect -32 11938 186 11948
rect -32 11882 -22 11938
rect 34 11882 120 11938
rect 176 11882 186 11938
rect -32 11796 186 11882
rect -32 11740 -22 11796
rect 34 11740 120 11796
rect 176 11740 186 11796
rect -32 11654 186 11740
rect -32 11598 -22 11654
rect 34 11598 120 11654
rect 176 11598 186 11654
rect -32 11512 186 11598
rect -32 11456 -22 11512
rect 34 11456 120 11512
rect 176 11456 186 11512
rect -32 11370 186 11456
rect -32 11314 -22 11370
rect 34 11314 120 11370
rect 176 11314 186 11370
rect -32 11228 186 11314
rect -32 11172 -22 11228
rect 34 11172 120 11228
rect 176 11172 186 11228
rect -32 11086 186 11172
rect -32 11030 -22 11086
rect 34 11030 120 11086
rect 176 11030 186 11086
rect -32 10944 186 11030
rect -32 10888 -22 10944
rect 34 10888 120 10944
rect 176 10888 186 10944
rect -32 10802 186 10888
rect -32 10746 -22 10802
rect 34 10746 120 10802
rect 176 10746 186 10802
rect -32 10660 186 10746
rect -32 10604 -22 10660
rect 34 10604 120 10660
rect 176 10604 186 10660
rect -32 10518 186 10604
rect -32 10462 -22 10518
rect 34 10462 120 10518
rect 176 10462 186 10518
rect -32 10376 186 10462
rect -32 10320 -22 10376
rect 34 10320 120 10376
rect 176 10320 186 10376
rect -32 10234 186 10320
rect -32 10178 -22 10234
rect 34 10178 120 10234
rect 176 10178 186 10234
rect -32 10092 186 10178
rect -32 10036 -22 10092
rect 34 10036 120 10092
rect 176 10036 186 10092
rect -32 9950 186 10036
rect -32 9894 -22 9950
rect 34 9894 120 9950
rect 176 9894 186 9950
rect -32 9808 186 9894
rect -32 9752 -22 9808
rect 34 9752 120 9808
rect 176 9752 186 9808
rect -32 9742 186 9752
rect -32 9426 186 9436
rect -32 9370 -22 9426
rect 34 9370 120 9426
rect 176 9370 186 9426
rect -32 9284 186 9370
rect -32 9228 -22 9284
rect 34 9228 120 9284
rect 176 9228 186 9284
rect -32 9142 186 9228
rect -32 9086 -22 9142
rect 34 9086 120 9142
rect 176 9086 186 9142
rect -32 9000 186 9086
rect -32 8944 -22 9000
rect 34 8944 120 9000
rect 176 8944 186 9000
rect -32 8858 186 8944
rect -32 8802 -22 8858
rect 34 8802 120 8858
rect 176 8802 186 8858
rect -32 8716 186 8802
rect -32 8660 -22 8716
rect 34 8660 120 8716
rect 176 8660 186 8716
rect -32 8574 186 8660
rect -32 8518 -22 8574
rect 34 8518 120 8574
rect 176 8518 186 8574
rect -32 8432 186 8518
rect -32 8376 -22 8432
rect 34 8376 120 8432
rect 176 8376 186 8432
rect -32 8290 186 8376
rect -32 8234 -22 8290
rect 34 8234 120 8290
rect 176 8234 186 8290
rect -32 8148 186 8234
rect -32 8092 -22 8148
rect 34 8092 120 8148
rect 176 8092 186 8148
rect -32 8006 186 8092
rect -32 7950 -22 8006
rect 34 7950 120 8006
rect 176 7950 186 8006
rect -32 7864 186 7950
rect -32 7808 -22 7864
rect 34 7808 120 7864
rect 176 7808 186 7864
rect -32 7722 186 7808
rect -32 7666 -22 7722
rect 34 7666 120 7722
rect 176 7666 186 7722
rect -32 7580 186 7666
rect -32 7524 -22 7580
rect 34 7524 120 7580
rect 176 7524 186 7580
rect -32 7438 186 7524
rect -32 7382 -22 7438
rect 34 7382 120 7438
rect 176 7382 186 7438
rect -32 7296 186 7382
rect -32 7240 -22 7296
rect 34 7240 120 7296
rect 176 7240 186 7296
rect -32 7154 186 7240
rect -32 7098 -22 7154
rect 34 7098 120 7154
rect 176 7098 186 7154
rect -32 7012 186 7098
rect -32 6956 -22 7012
rect 34 6956 120 7012
rect 176 6956 186 7012
rect -32 6870 186 6956
rect -32 6814 -22 6870
rect 34 6814 120 6870
rect 176 6814 186 6870
rect -32 6728 186 6814
rect -32 6672 -22 6728
rect 34 6672 120 6728
rect 176 6672 186 6728
rect -32 6586 186 6672
rect -32 6530 -22 6586
rect 34 6530 120 6586
rect 176 6530 186 6586
rect -32 6520 186 6530
rect -32 6239 186 6249
rect -32 6183 -22 6239
rect 34 6183 120 6239
rect 176 6183 186 6239
rect -32 6097 186 6183
rect -32 6041 -22 6097
rect 34 6041 120 6097
rect 176 6041 186 6097
rect -32 5955 186 6041
rect -32 5899 -22 5955
rect 34 5899 120 5955
rect 176 5899 186 5955
rect -32 5813 186 5899
rect -32 5757 -22 5813
rect 34 5757 120 5813
rect 176 5757 186 5813
rect -32 5671 186 5757
rect -32 5615 -22 5671
rect 34 5615 120 5671
rect 176 5615 186 5671
rect -32 5529 186 5615
rect -32 5473 -22 5529
rect 34 5473 120 5529
rect 176 5473 186 5529
rect -32 5387 186 5473
rect -32 5331 -22 5387
rect 34 5331 120 5387
rect 176 5331 186 5387
rect -32 5245 186 5331
rect -32 5189 -22 5245
rect 34 5189 120 5245
rect 176 5189 186 5245
rect -32 5103 186 5189
rect -32 5047 -22 5103
rect 34 5047 120 5103
rect 176 5047 186 5103
rect -32 4961 186 5047
rect -32 4905 -22 4961
rect 34 4905 120 4961
rect 176 4905 186 4961
rect -32 4819 186 4905
rect -32 4763 -22 4819
rect 34 4763 120 4819
rect 176 4763 186 4819
rect -32 4677 186 4763
rect -32 4621 -22 4677
rect 34 4621 120 4677
rect 176 4621 186 4677
rect -32 4535 186 4621
rect -32 4479 -22 4535
rect 34 4479 120 4535
rect 176 4479 186 4535
rect -32 4393 186 4479
rect -32 4337 -22 4393
rect 34 4337 120 4393
rect 176 4337 186 4393
rect -32 4251 186 4337
rect -32 4195 -22 4251
rect 34 4195 120 4251
rect 176 4195 186 4251
rect -32 4109 186 4195
rect -32 4053 -22 4109
rect 34 4053 120 4109
rect 176 4053 186 4109
rect -32 3967 186 4053
rect -32 3911 -22 3967
rect 34 3911 120 3967
rect 176 3911 186 3967
rect -32 3825 186 3911
rect -32 3769 -22 3825
rect 34 3769 120 3825
rect 176 3769 186 3825
rect -32 3683 186 3769
rect -32 3627 -22 3683
rect 34 3627 120 3683
rect 176 3627 186 3683
rect -32 3541 186 3627
rect -32 3485 -22 3541
rect 34 3485 120 3541
rect 176 3485 186 3541
rect -32 3399 186 3485
rect -32 3343 -22 3399
rect 34 3343 120 3399
rect 176 3343 186 3399
rect -32 3333 186 3343
rect -32 3051 186 3061
rect -32 2995 -22 3051
rect 34 2995 120 3051
rect 176 2995 186 3051
rect -32 2909 186 2995
rect -32 2853 -22 2909
rect 34 2853 120 2909
rect 176 2853 186 2909
rect -32 2767 186 2853
rect -32 2711 -22 2767
rect 34 2711 120 2767
rect 176 2711 186 2767
rect -32 2625 186 2711
rect -32 2569 -22 2625
rect 34 2569 120 2625
rect 176 2569 186 2625
rect -32 2483 186 2569
rect -32 2427 -22 2483
rect 34 2427 120 2483
rect 176 2427 186 2483
rect -32 2341 186 2427
rect -32 2285 -22 2341
rect 34 2285 120 2341
rect 176 2285 186 2341
rect -32 2199 186 2285
rect -32 2143 -22 2199
rect 34 2143 120 2199
rect 176 2143 186 2199
rect -32 2057 186 2143
rect -32 2001 -22 2057
rect 34 2001 120 2057
rect 176 2001 186 2057
rect -32 1915 186 2001
rect -32 1859 -22 1915
rect 34 1859 120 1915
rect 176 1859 186 1915
rect -32 1773 186 1859
rect -32 1717 -22 1773
rect 34 1717 120 1773
rect 176 1717 186 1773
rect -32 1631 186 1717
rect -32 1575 -22 1631
rect 34 1575 120 1631
rect 176 1575 186 1631
rect -32 1489 186 1575
rect -32 1433 -22 1489
rect 34 1433 120 1489
rect 176 1433 186 1489
rect -32 1347 186 1433
rect -32 1291 -22 1347
rect 34 1291 120 1347
rect 176 1291 186 1347
rect -32 1205 186 1291
rect -32 1149 -22 1205
rect 34 1149 120 1205
rect 176 1149 186 1205
rect -32 1063 186 1149
rect -32 1007 -22 1063
rect 34 1007 120 1063
rect 176 1007 186 1063
rect -32 921 186 1007
rect -32 865 -22 921
rect 34 865 120 921
rect 176 865 186 921
rect -32 779 186 865
rect -32 723 -22 779
rect 34 723 120 779
rect 176 723 186 779
rect -32 637 186 723
rect -32 581 -22 637
rect 34 581 120 637
rect 176 581 186 637
rect -32 495 186 581
rect -32 439 -22 495
rect 34 439 120 495
rect 176 439 186 495
rect -32 353 186 439
rect -32 297 -22 353
rect 34 297 120 353
rect 176 297 186 353
rect -32 211 186 297
rect -32 155 -22 211
rect 34 155 120 211
rect 176 155 186 211
rect -32 145 186 155
use M2_M1_CDNS_40661953145300  M2_M1_CDNS_40661953145300_0
timestamp 1749760379
transform 1 0 962 0 1 5990
box 0 0 1 1
use M2_M1_CDNS_40661953145301  M2_M1_CDNS_40661953145301_0
timestamp 1749760379
transform 1 0 78 0 1 5990
box 0 0 1 1
use M3_M2_CDNS_40661953145208  M3_M2_CDNS_40661953145208_0
timestamp 1749760379
transform 1 0 77 0 1 1603
box 0 0 1 1
use M3_M2_CDNS_40661953145208  M3_M2_CDNS_40661953145208_1
timestamp 1749760379
transform 1 0 77 0 1 4791
box 0 0 1 1
use M3_M2_CDNS_40661953145208  M3_M2_CDNS_40661953145208_2
timestamp 1749760379
transform 1 0 77 0 1 7978
box 0 0 1 1
use M3_M2_CDNS_40661953145302  M3_M2_CDNS_40661953145302_0
timestamp 1749760379
transform 1 0 77 0 1 10845
box 0 0 1 1
<< properties >>
string GDS_END 2653018
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2652458
<< end >>
