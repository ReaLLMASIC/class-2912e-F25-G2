magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 453 982 1094
<< pwell >>
rect -86 -86 982 453
<< metal1 >>
rect 0 918 896 1098
rect 353 710 399 918
rect 49 90 95 298
rect 801 710 847 918
rect 497 90 543 298
rect 0 -90 896 90
<< obsm1 >>
rect 49 412 95 872
rect 254 494 399 540
rect 49 366 194 412
rect 353 136 399 494
rect 497 412 543 872
rect 702 494 847 540
rect 497 366 642 412
rect 801 136 847 494
<< labels >>
rlabel metal1 s 801 710 847 918 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 710 399 918 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 918 896 1098 6 VDD
port 1 nsew power bidirectional abutment
rlabel nwell s -86 453 982 1094 6 VNW
port 2 nsew power bidirectional
rlabel pwell s -86 -86 982 453 6 VPW
port 3 nsew ground bidirectional
rlabel metal1 s 0 -90 896 90 8 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 298 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 298 6 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 896 1008
string LEFclass core SPACER
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 779450
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 776048
<< end >>
