magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 355 4230 870
rect -86 352 952 355
rect 2142 352 4230 355
<< pwell >>
rect 952 352 2142 355
rect -86 -86 4230 352
<< mvnmos >>
rect 124 153 244 232
rect 348 153 468 232
rect 572 153 692 232
rect 799 153 919 232
rect 1059 156 1179 235
rect 1315 156 1435 235
rect 1683 156 1803 235
rect 1907 156 2027 235
rect 2395 93 2515 188
rect 2619 93 2739 188
rect 2843 93 2963 188
rect 3211 93 3331 219
rect 3435 93 3555 219
rect 3659 93 3779 219
rect 3883 93 4003 219
<< mvpmos >>
rect 144 475 244 660
rect 348 475 448 660
rect 588 515 688 668
rect 887 515 987 668
rect 1127 475 1227 628
rect 1335 475 1435 628
rect 1683 475 1783 628
rect 1907 475 2007 628
rect 2431 472 2531 703
rect 2635 472 2735 703
rect 2783 472 2883 703
rect 3173 472 3273 716
rect 3377 472 3477 716
rect 3581 472 3681 716
rect 3785 472 3885 716
<< mvndiff >>
rect 979 232 1059 235
rect 36 215 124 232
rect 36 169 49 215
rect 95 169 124 215
rect 36 153 124 169
rect 244 212 348 232
rect 244 166 273 212
rect 319 166 348 212
rect 244 153 348 166
rect 468 215 572 232
rect 468 169 497 215
rect 543 169 572 215
rect 468 153 572 169
rect 692 215 799 232
rect 692 169 721 215
rect 767 169 799 215
rect 692 153 799 169
rect 919 156 1059 232
rect 1179 215 1315 235
rect 1179 169 1224 215
rect 1270 169 1315 215
rect 1179 156 1315 169
rect 1435 215 1523 235
rect 1435 169 1464 215
rect 1510 169 1523 215
rect 1435 156 1523 169
rect 1595 215 1683 235
rect 1595 169 1608 215
rect 1654 169 1683 215
rect 1595 156 1683 169
rect 1803 215 1907 235
rect 1803 169 1832 215
rect 1878 169 1907 215
rect 1803 156 1907 169
rect 2027 215 2115 235
rect 2027 169 2056 215
rect 2102 169 2115 215
rect 2027 156 2115 169
rect 919 153 999 156
rect 2307 152 2395 188
rect 2307 106 2320 152
rect 2366 106 2395 152
rect 2307 93 2395 106
rect 2515 152 2619 188
rect 2515 106 2544 152
rect 2590 106 2619 152
rect 2515 93 2619 106
rect 2739 152 2843 188
rect 2739 106 2768 152
rect 2814 106 2843 152
rect 2739 93 2843 106
rect 2963 152 3051 188
rect 2963 106 2992 152
rect 3038 106 3051 152
rect 2963 93 3051 106
rect 3123 178 3211 219
rect 3123 132 3136 178
rect 3182 132 3211 178
rect 3123 93 3211 132
rect 3331 189 3435 219
rect 3331 143 3360 189
rect 3406 143 3435 189
rect 3331 93 3435 143
rect 3555 172 3659 219
rect 3555 126 3584 172
rect 3630 126 3659 172
rect 3555 93 3659 126
rect 3779 189 3883 219
rect 3779 143 3808 189
rect 3854 143 3883 189
rect 3779 93 3883 143
rect 4003 172 4091 219
rect 4003 126 4032 172
rect 4078 126 4091 172
rect 4003 93 4091 126
<< mvpdiff >>
rect 508 660 588 668
rect 56 647 144 660
rect 56 507 69 647
rect 115 507 144 647
rect 56 475 144 507
rect 244 475 348 660
rect 448 515 588 660
rect 688 614 887 668
rect 688 568 762 614
rect 808 568 887 614
rect 688 515 887 568
rect 987 628 1067 668
rect 987 515 1127 628
rect 448 475 528 515
rect 1047 475 1127 515
rect 1227 615 1335 628
rect 1227 569 1260 615
rect 1306 569 1335 615
rect 1227 475 1335 569
rect 1435 567 1523 628
rect 1435 521 1464 567
rect 1510 521 1523 567
rect 1435 475 1523 521
rect 1595 567 1683 628
rect 1595 521 1608 567
rect 1654 521 1683 567
rect 1595 475 1683 521
rect 1783 568 1907 628
rect 1783 522 1822 568
rect 1868 522 1907 568
rect 1783 475 1907 522
rect 2007 568 2095 628
rect 2007 522 2036 568
rect 2082 522 2095 568
rect 2007 475 2095 522
rect 2343 567 2431 703
rect 2343 521 2356 567
rect 2402 521 2431 567
rect 2343 472 2431 521
rect 2531 680 2635 703
rect 2531 540 2560 680
rect 2606 540 2635 680
rect 2531 472 2635 540
rect 2735 472 2783 703
rect 2883 625 2971 703
rect 2883 485 2912 625
rect 2958 485 2971 625
rect 2883 472 2971 485
rect 3085 680 3173 716
rect 3085 540 3098 680
rect 3144 540 3173 680
rect 3085 472 3173 540
rect 3273 625 3377 716
rect 3273 485 3302 625
rect 3348 485 3377 625
rect 3273 472 3377 485
rect 3477 661 3581 716
rect 3477 615 3506 661
rect 3552 615 3581 661
rect 3477 472 3581 615
rect 3681 625 3785 716
rect 3681 485 3710 625
rect 3756 485 3785 625
rect 3681 472 3785 485
rect 3885 661 3973 716
rect 3885 615 3914 661
rect 3960 615 3973 661
rect 3885 472 3973 615
<< mvndiffc >>
rect 49 169 95 215
rect 273 166 319 212
rect 497 169 543 215
rect 721 169 767 215
rect 1224 169 1270 215
rect 1464 169 1510 215
rect 1608 169 1654 215
rect 1832 169 1878 215
rect 2056 169 2102 215
rect 2320 106 2366 152
rect 2544 106 2590 152
rect 2768 106 2814 152
rect 2992 106 3038 152
rect 3136 132 3182 178
rect 3360 143 3406 189
rect 3584 126 3630 172
rect 3808 143 3854 189
rect 4032 126 4078 172
<< mvpdiffc >>
rect 69 507 115 647
rect 762 568 808 614
rect 1260 569 1306 615
rect 1464 521 1510 567
rect 1608 521 1654 567
rect 1822 522 1868 568
rect 2036 522 2082 568
rect 2356 521 2402 567
rect 2560 540 2606 680
rect 2912 485 2958 625
rect 3098 540 3144 680
rect 3302 485 3348 625
rect 3506 615 3552 661
rect 3710 485 3756 625
rect 3914 615 3960 661
<< polysilicon >>
rect 1127 720 2007 760
rect 144 660 244 704
rect 348 660 448 704
rect 588 668 688 712
rect 887 668 987 712
rect 1127 628 1227 720
rect 1335 628 1435 672
rect 1683 628 1783 672
rect 1907 628 2007 720
rect 2431 703 2531 747
rect 2635 703 2735 747
rect 2783 703 2883 747
rect 3173 716 3273 760
rect 3377 716 3477 760
rect 3581 716 3681 760
rect 3785 716 3885 760
rect 144 415 244 475
rect 144 369 159 415
rect 205 369 244 415
rect 144 279 244 369
rect 124 232 244 279
rect 348 415 448 475
rect 588 455 688 515
rect 588 415 839 455
rect 348 369 387 415
rect 433 369 448 415
rect 348 279 448 369
rect 572 354 751 367
rect 572 308 692 354
rect 738 308 751 354
rect 572 295 751 308
rect 348 232 468 279
rect 572 232 692 295
rect 799 279 839 415
rect 887 420 987 515
rect 887 374 913 420
rect 959 374 987 420
rect 887 361 987 374
rect 1127 335 1227 475
rect 1059 295 1227 335
rect 799 232 919 279
rect 1059 235 1179 295
rect 1335 279 1435 475
rect 1315 235 1435 279
rect 1683 426 1783 475
rect 1683 380 1712 426
rect 1758 380 1783 426
rect 1683 279 1783 380
rect 1907 314 2007 475
rect 1683 235 1803 279
rect 1907 268 1925 314
rect 1971 279 2007 314
rect 2431 428 2531 472
rect 2635 428 2735 472
rect 2431 304 2515 428
rect 1971 268 2027 279
rect 1907 235 2027 268
rect 2431 258 2451 304
rect 2497 258 2515 304
rect 2431 232 2515 258
rect 2635 382 2659 428
rect 2705 382 2735 428
rect 2635 232 2735 382
rect 2783 428 2883 472
rect 2783 382 2805 428
rect 2851 382 2883 428
rect 2783 369 2883 382
rect 2843 232 2883 369
rect 3173 417 3273 472
rect 3173 371 3201 417
rect 3247 398 3273 417
rect 3377 417 3477 472
rect 3377 398 3395 417
rect 3247 371 3395 398
rect 3441 398 3477 417
rect 3581 417 3681 472
rect 3581 398 3608 417
rect 3441 371 3608 398
rect 3654 398 3681 417
rect 3785 417 3885 472
rect 3785 398 3810 417
rect 3654 371 3810 398
rect 3856 398 3885 417
rect 3856 371 3923 398
rect 3173 358 3923 371
rect 3211 263 3273 358
rect 3435 263 3477 358
rect 3659 263 3717 358
rect 3883 263 3923 358
rect 2395 188 2515 232
rect 2619 188 2739 232
rect 2843 188 2963 232
rect 3211 219 3331 263
rect 3435 219 3555 263
rect 3659 219 3779 263
rect 3883 219 4003 263
rect 124 109 244 153
rect 348 109 468 153
rect 572 109 692 153
rect 799 64 919 153
rect 1059 112 1179 156
rect 1315 64 1435 156
rect 1683 112 1803 156
rect 1907 112 2027 156
rect 2175 152 2247 165
rect 2175 106 2188 152
rect 2234 106 2247 152
rect 2175 64 2247 106
rect 799 24 2247 64
rect 2395 49 2515 93
rect 2619 49 2739 93
rect 2843 49 2963 93
rect 3211 49 3331 93
rect 3435 49 3555 93
rect 3659 49 3779 93
rect 3883 49 4003 93
<< polycontact >>
rect 159 369 205 415
rect 387 369 433 415
rect 692 308 738 354
rect 913 374 959 420
rect 1712 380 1758 426
rect 1925 268 1971 314
rect 2451 258 2497 304
rect 2659 382 2705 428
rect 2805 382 2851 428
rect 3201 371 3247 417
rect 3395 371 3441 417
rect 3608 371 3654 417
rect 3810 371 3856 417
rect 2188 106 2234 152
<< metal1 >>
rect 0 724 4144 844
rect 69 647 115 724
rect 69 496 115 507
rect 468 424 550 674
rect 762 614 808 653
rect 762 512 808 568
rect 1260 615 1306 724
rect 1260 558 1306 569
rect 1362 632 1758 678
rect 1362 512 1408 632
rect 58 415 318 424
rect 58 369 159 415
rect 205 369 318 415
rect 58 360 318 369
rect 373 415 550 424
rect 373 369 387 415
rect 433 369 550 415
rect 373 360 550 369
rect 600 466 1408 512
rect 1464 567 1510 580
rect 38 261 423 308
rect 38 215 106 261
rect 38 169 49 215
rect 95 169 106 215
rect 377 215 423 261
rect 600 215 646 466
rect 1464 420 1510 521
rect 692 374 913 420
rect 959 374 1510 420
rect 692 354 738 374
rect 692 284 738 308
rect 1464 215 1510 374
rect 262 166 273 212
rect 319 166 330 212
rect 377 169 497 215
rect 543 169 554 215
rect 600 169 721 215
rect 767 169 778 215
rect 1213 169 1224 215
rect 1270 169 1281 215
rect 262 60 330 166
rect 1213 60 1281 169
rect 1464 156 1510 169
rect 1608 567 1654 580
rect 1608 315 1654 521
rect 1712 426 1758 632
rect 1822 568 1868 724
rect 2560 680 2606 724
rect 1822 494 1868 522
rect 2036 632 2514 678
rect 2036 568 2102 632
rect 2082 522 2102 568
rect 1712 364 1758 380
rect 1608 314 1982 315
rect 1608 268 1925 314
rect 1971 268 1982 314
rect 1608 215 1654 268
rect 2036 215 2102 522
rect 2356 567 2402 586
rect 2356 499 2402 521
rect 1608 156 1654 169
rect 1821 169 1832 215
rect 1878 169 1889 215
rect 1821 60 1889 169
rect 2036 169 2056 215
rect 2036 156 2102 169
rect 2172 452 2402 499
rect 2172 152 2218 452
rect 2468 428 2514 632
rect 3098 680 3144 724
rect 2560 529 2606 540
rect 2912 625 2958 636
rect 3506 661 3552 724
rect 3098 529 3144 540
rect 3302 625 3348 636
rect 2805 428 2851 439
rect 2468 382 2659 428
rect 2705 382 2726 428
rect 2805 336 2851 382
rect 2714 318 2851 336
rect 2362 304 2851 318
rect 2362 258 2451 304
rect 2497 290 2851 304
rect 2912 428 2958 485
rect 3914 661 3960 724
rect 3506 604 3552 615
rect 3710 625 3756 636
rect 3348 485 3710 542
rect 3914 604 3960 615
rect 3756 485 4014 542
rect 3302 474 4014 485
rect 2912 417 3856 428
rect 2912 371 3201 417
rect 3247 371 3395 417
rect 3441 371 3608 417
rect 3654 371 3810 417
rect 2912 358 3856 371
rect 2497 258 2773 290
rect 2362 242 2773 258
rect 2912 244 2958 358
rect 3938 307 4014 474
rect 2868 198 2958 244
rect 3350 253 4014 307
rect 2868 152 2914 198
rect 3136 178 3182 218
rect 2172 106 2188 152
rect 2234 106 2320 152
rect 2366 106 2395 152
rect 2533 106 2544 152
rect 2590 106 2601 152
rect 2757 106 2768 152
rect 2814 106 2914 152
rect 2981 106 2992 152
rect 3038 106 3049 152
rect 2533 60 2601 106
rect 2981 60 3049 106
rect 3136 60 3182 132
rect 3350 189 3444 253
rect 3350 143 3360 189
rect 3406 143 3444 189
rect 3350 120 3444 143
rect 3584 172 3630 195
rect 3584 60 3630 126
rect 3808 189 3894 253
rect 3854 143 3894 189
rect 3808 120 3894 143
rect 4032 172 4078 195
rect 4032 60 4078 126
rect 0 -60 4144 60
<< labels >>
flabel metal1 s 3710 542 3756 636 0 FreeSans 400 0 0 0 Q
port 4 nsew default output
flabel metal1 s 58 360 318 424 0 FreeSans 400 0 0 0 TE
port 3 nsew default input
flabel metal1 s 0 724 4144 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 3136 215 3182 218 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 2805 336 2851 439 0 FreeSans 400 0 0 0 CLKN
port 1 nsew clock input
flabel metal1 s 468 424 550 674 0 FreeSans 400 0 0 0 E
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 2714 318 2851 336 1 CLKN
port 1 nsew clock input
rlabel metal1 s 2362 290 2851 318 1 CLKN
port 1 nsew clock input
rlabel metal1 s 2362 242 2773 290 1 CLKN
port 1 nsew clock input
rlabel metal1 s 373 360 550 424 1 E
port 2 nsew default input
rlabel metal1 s 3302 542 3348 636 1 Q
port 4 nsew default output
rlabel metal1 s 3302 474 4014 542 1 Q
port 4 nsew default output
rlabel metal1 s 3938 307 4014 474 1 Q
port 4 nsew default output
rlabel metal1 s 3350 253 4014 307 1 Q
port 4 nsew default output
rlabel metal1 s 3808 120 3894 253 1 Q
port 4 nsew default output
rlabel metal1 s 3350 120 3444 253 1 Q
port 4 nsew default output
rlabel metal1 s 3914 604 3960 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3506 604 3552 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3098 604 3144 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2560 604 2606 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1822 604 1868 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1260 604 1306 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 604 115 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3098 558 3144 604 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2560 558 2606 604 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1822 558 1868 604 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1260 558 1306 604 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 558 115 604 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3098 529 3144 558 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2560 529 2606 558 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1822 529 1868 558 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 529 115 558 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1822 496 1868 529 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 496 115 529 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1822 494 1868 496 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3136 212 3182 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1821 212 1889 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1213 212 1281 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3136 195 3182 212 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1821 195 1889 212 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1213 195 1281 212 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 195 330 212 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4032 152 4078 195 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3584 152 3630 195 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3136 152 3182 195 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1821 152 1889 195 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1213 152 1281 195 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 152 330 195 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4032 60 4078 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3584 60 3630 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3136 60 3182 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2981 60 3049 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2533 60 2601 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1821 60 1889 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1213 60 1281 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4144 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4144 784
string GDS_END 450676
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 441986
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
