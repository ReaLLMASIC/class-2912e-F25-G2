magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect 29138 66274 56005 66790
rect 29138 65155 32850 66274
rect 29138 35918 33473 65155
rect 35260 65135 39818 66274
rect 42526 65785 43793 66075
rect 42526 65708 44118 65785
rect 42527 65135 44118 65708
rect 45169 65154 49764 66274
rect 35260 65105 39464 65135
rect 35124 65033 39464 65105
rect 35124 35949 37639 65033
rect 30658 35917 33473 35918
rect 31003 35899 33473 35917
rect 38864 35899 39464 65033
rect 44662 65104 49764 65154
rect 52285 65136 56005 66274
rect 44662 35950 50000 65104
rect 51652 65033 56005 65136
rect 44662 35900 48709 35950
rect 51652 35918 55985 65033
rect 54025 35917 54467 35918
<< pwell >>
rect 1774 65882 24710 65914
rect 1774 35138 24710 35170
<< mvnmos >>
rect 33001 65399 35023 65519
rect 40062 65399 40590 65519
rect 40963 65400 42281 65520
rect 44432 65399 44960 65519
rect 50001 65399 52023 65519
rect 33671 64755 34671 64875
rect 39727 64755 40167 64875
rect 43695 64744 44325 64864
rect 33671 64531 34671 64651
rect 50454 64755 51454 64875
rect 33671 64275 34671 64395
rect 37896 64444 38556 64564
rect 43695 64531 44325 64651
rect 37896 64220 38556 64340
rect 39598 64220 39730 64340
rect 43695 64307 44325 64427
rect 50454 64531 51454 64651
rect 50454 64275 51454 64395
rect 33671 63659 34671 63779
rect 33671 63403 34671 63523
rect 37896 63714 38556 63834
rect 37896 63490 38556 63610
rect 39598 63714 39730 63834
rect 43695 63627 44325 63747
rect 50454 63659 51454 63779
rect 43695 63403 44325 63523
rect 50454 63403 51454 63523
rect 33671 63179 34671 63299
rect 33671 62955 34671 63075
rect 39727 63179 40167 63299
rect 43695 63190 44325 63310
rect 39727 62955 40167 63075
rect 50454 63179 51454 63299
rect 43695 62944 44325 63064
rect 33671 62731 34671 62851
rect 50454 62955 51454 63075
rect 33671 62475 34671 62595
rect 37896 62644 38556 62764
rect 43695 62731 44325 62851
rect 37896 62420 38556 62540
rect 39598 62420 39730 62540
rect 43695 62507 44325 62627
rect 50454 62731 51454 62851
rect 50454 62475 51454 62595
rect 33671 61859 34671 61979
rect 33671 61603 34671 61723
rect 37896 61914 38556 62034
rect 37896 61690 38556 61810
rect 39598 61914 39730 62034
rect 43695 61827 44325 61947
rect 50454 61859 51454 61979
rect 43695 61603 44325 61723
rect 50454 61603 51454 61723
rect 33671 61379 34671 61499
rect 33671 61155 34671 61275
rect 39727 61379 40167 61499
rect 43695 61390 44325 61510
rect 39727 61155 40167 61275
rect 50454 61379 51454 61499
rect 43695 61144 44325 61264
rect 33671 60931 34671 61051
rect 50454 61155 51454 61275
rect 33671 60675 34671 60795
rect 37896 60844 38556 60964
rect 43695 60931 44325 61051
rect 37896 60620 38556 60740
rect 39598 60620 39730 60740
rect 43695 60707 44325 60827
rect 50454 60931 51454 61051
rect 50454 60675 51454 60795
rect 33671 60059 34671 60179
rect 33671 59803 34671 59923
rect 37896 60114 38556 60234
rect 37896 59890 38556 60010
rect 39598 60114 39730 60234
rect 43695 60027 44325 60147
rect 50454 60059 51454 60179
rect 43695 59803 44325 59923
rect 50454 59803 51454 59923
rect 33671 59579 34671 59699
rect 33671 59355 34671 59475
rect 39727 59579 40167 59699
rect 43695 59590 44325 59710
rect 39727 59355 40167 59475
rect 50454 59579 51454 59699
rect 43695 59344 44325 59464
rect 33671 59131 34671 59251
rect 50454 59355 51454 59475
rect 33671 58875 34671 58995
rect 37896 59044 38556 59164
rect 43695 59131 44325 59251
rect 37896 58820 38556 58940
rect 39598 58820 39730 58940
rect 43695 58907 44325 59027
rect 50454 59131 51454 59251
rect 50454 58875 51454 58995
rect 33671 58259 34671 58379
rect 33671 58003 34671 58123
rect 37896 58314 38556 58434
rect 37896 58090 38556 58210
rect 39598 58314 39730 58434
rect 43695 58227 44325 58347
rect 50454 58259 51454 58379
rect 43695 58003 44325 58123
rect 50454 58003 51454 58123
rect 33671 57779 34671 57899
rect 33671 57555 34671 57675
rect 39727 57779 40167 57899
rect 43695 57790 44325 57910
rect 39727 57555 40167 57675
rect 50454 57779 51454 57899
rect 43695 57544 44325 57664
rect 33671 57331 34671 57451
rect 50454 57555 51454 57675
rect 33671 57075 34671 57195
rect 37896 57244 38556 57364
rect 43695 57331 44325 57451
rect 37896 57020 38556 57140
rect 39598 57020 39730 57140
rect 43695 57107 44325 57227
rect 50454 57331 51454 57451
rect 50454 57075 51454 57195
rect 33671 56459 34671 56579
rect 33671 56203 34671 56323
rect 37896 56514 38556 56634
rect 37896 56290 38556 56410
rect 39598 56514 39730 56634
rect 43695 56427 44325 56547
rect 50454 56459 51454 56579
rect 43695 56203 44325 56323
rect 50454 56203 51454 56323
rect 33671 55979 34671 56099
rect 33671 55755 34671 55875
rect 39727 55979 40167 56099
rect 43695 55990 44325 56110
rect 39727 55755 40167 55875
rect 50454 55979 51454 56099
rect 43695 55744 44325 55864
rect 33671 55531 34671 55651
rect 50454 55755 51454 55875
rect 33671 55275 34671 55395
rect 37896 55444 38556 55564
rect 43695 55531 44325 55651
rect 37896 55220 38556 55340
rect 39598 55220 39730 55340
rect 43695 55307 44325 55427
rect 50454 55531 51454 55651
rect 50454 55275 51454 55395
rect 33671 54659 34671 54779
rect 33671 54403 34671 54523
rect 37896 54714 38556 54834
rect 37896 54490 38556 54610
rect 39598 54714 39730 54834
rect 43695 54627 44325 54747
rect 50454 54659 51454 54779
rect 43695 54403 44325 54523
rect 50454 54403 51454 54523
rect 33671 54179 34671 54299
rect 33671 53955 34671 54075
rect 39727 54179 40167 54299
rect 43695 54190 44325 54310
rect 39727 53955 40167 54075
rect 50454 54179 51454 54299
rect 43695 53944 44325 54064
rect 33671 53731 34671 53851
rect 50454 53955 51454 54075
rect 33671 53475 34671 53595
rect 37896 53644 38556 53764
rect 43695 53731 44325 53851
rect 37896 53420 38556 53540
rect 39598 53420 39730 53540
rect 43695 53507 44325 53627
rect 50454 53731 51454 53851
rect 50454 53475 51454 53595
rect 33671 52859 34671 52979
rect 33671 52603 34671 52723
rect 37896 52914 38556 53034
rect 37896 52690 38556 52810
rect 39598 52914 39730 53034
rect 43695 52827 44325 52947
rect 50454 52859 51454 52979
rect 43695 52603 44325 52723
rect 50454 52603 51454 52723
rect 33671 52379 34671 52499
rect 33671 52155 34671 52275
rect 39727 52379 40167 52499
rect 43695 52390 44325 52510
rect 39727 52155 40167 52275
rect 50454 52379 51454 52499
rect 43695 52144 44325 52264
rect 33671 51931 34671 52051
rect 50454 52155 51454 52275
rect 33671 51675 34671 51795
rect 37896 51844 38556 51964
rect 43695 51931 44325 52051
rect 37896 51620 38556 51740
rect 39598 51620 39730 51740
rect 43695 51707 44325 51827
rect 50454 51931 51454 52051
rect 50454 51675 51454 51795
rect 33671 51059 34671 51179
rect 33671 50803 34671 50923
rect 37896 51114 38556 51234
rect 37896 50890 38556 51010
rect 39598 51114 39730 51234
rect 43695 51027 44325 51147
rect 50454 51059 51454 51179
rect 43695 50803 44325 50923
rect 50454 50803 51454 50923
rect 33671 50579 34671 50699
rect 33671 50355 34671 50475
rect 39727 50579 40167 50699
rect 43695 50590 44325 50710
rect 39727 50355 40167 50475
rect 50454 50579 51454 50699
rect 43695 50344 44325 50464
rect 33671 50131 34671 50251
rect 50454 50355 51454 50475
rect 33671 49875 34671 49995
rect 37896 50044 38556 50164
rect 43695 50131 44325 50251
rect 37896 49820 38556 49940
rect 39598 49820 39730 49940
rect 43695 49907 44325 50027
rect 50454 50131 51454 50251
rect 50454 49875 51454 49995
rect 33671 49259 34671 49379
rect 33671 49003 34671 49123
rect 37896 49314 38556 49434
rect 37896 49090 38556 49210
rect 39598 49314 39730 49434
rect 43695 49227 44325 49347
rect 50454 49259 51454 49379
rect 43695 49003 44325 49123
rect 50454 49003 51454 49123
rect 33671 48779 34671 48899
rect 33671 48555 34671 48675
rect 39727 48779 40167 48899
rect 43695 48790 44325 48910
rect 39727 48555 40167 48675
rect 50454 48779 51454 48899
rect 43695 48544 44325 48664
rect 33671 48331 34671 48451
rect 50454 48555 51454 48675
rect 33671 48075 34671 48195
rect 37896 48244 38556 48364
rect 43695 48331 44325 48451
rect 37896 48020 38556 48140
rect 39598 48020 39730 48140
rect 43695 48107 44325 48227
rect 50454 48331 51454 48451
rect 50454 48075 51454 48195
rect 33671 47459 34671 47579
rect 33671 47203 34671 47323
rect 37896 47514 38556 47634
rect 37896 47290 38556 47410
rect 39598 47514 39730 47634
rect 43695 47427 44325 47547
rect 50454 47459 51454 47579
rect 43695 47203 44325 47323
rect 50454 47203 51454 47323
rect 33671 46979 34671 47099
rect 33671 46755 34671 46875
rect 39727 46979 40167 47099
rect 43695 46990 44325 47110
rect 39727 46755 40167 46875
rect 50454 46979 51454 47099
rect 43695 46744 44325 46864
rect 33671 46531 34671 46651
rect 50454 46755 51454 46875
rect 33671 46275 34671 46395
rect 37896 46444 38556 46564
rect 43695 46531 44325 46651
rect 37896 46220 38556 46340
rect 39598 46220 39730 46340
rect 43695 46307 44325 46427
rect 50454 46531 51454 46651
rect 50454 46275 51454 46395
rect 33671 45659 34671 45779
rect 33671 45403 34671 45523
rect 37896 45714 38556 45834
rect 37896 45490 38556 45610
rect 39598 45714 39730 45834
rect 43695 45627 44325 45747
rect 50454 45659 51454 45779
rect 43695 45403 44325 45523
rect 50454 45403 51454 45523
rect 33671 45179 34671 45299
rect 33671 44955 34671 45075
rect 39727 45179 40167 45299
rect 43695 45190 44325 45310
rect 39727 44955 40167 45075
rect 50454 45179 51454 45299
rect 43695 44944 44325 45064
rect 33671 44731 34671 44851
rect 50454 44955 51454 45075
rect 33671 44475 34671 44595
rect 37896 44644 38556 44764
rect 43695 44731 44325 44851
rect 37896 44420 38556 44540
rect 39598 44420 39730 44540
rect 43695 44507 44325 44627
rect 50454 44731 51454 44851
rect 50454 44475 51454 44595
rect 33671 43859 34671 43979
rect 33671 43603 34671 43723
rect 37896 43914 38556 44034
rect 37896 43690 38556 43810
rect 39598 43914 39730 44034
rect 43695 43827 44325 43947
rect 50454 43859 51454 43979
rect 43695 43603 44325 43723
rect 50454 43603 51454 43723
rect 33671 43379 34671 43499
rect 33671 43155 34671 43275
rect 39727 43379 40167 43499
rect 43695 43390 44325 43510
rect 39727 43155 40167 43275
rect 50454 43379 51454 43499
rect 43695 43144 44325 43264
rect 33671 42931 34671 43051
rect 50454 43155 51454 43275
rect 33671 42675 34671 42795
rect 37896 42844 38556 42964
rect 43695 42931 44325 43051
rect 37896 42620 38556 42740
rect 39598 42620 39730 42740
rect 43695 42707 44325 42827
rect 50454 42931 51454 43051
rect 50454 42675 51454 42795
rect 33671 42059 34671 42179
rect 33671 41803 34671 41923
rect 37896 42114 38556 42234
rect 37896 41890 38556 42010
rect 39598 42114 39730 42234
rect 43695 42027 44325 42147
rect 50454 42059 51454 42179
rect 43695 41803 44325 41923
rect 50454 41803 51454 41923
rect 33671 41579 34671 41699
rect 33671 41355 34671 41475
rect 39727 41579 40167 41699
rect 43695 41590 44325 41710
rect 39727 41355 40167 41475
rect 50454 41579 51454 41699
rect 43695 41344 44325 41464
rect 33671 41131 34671 41251
rect 50454 41355 51454 41475
rect 33671 40875 34671 40995
rect 37896 41044 38556 41164
rect 43695 41131 44325 41251
rect 37896 40820 38556 40940
rect 39598 40820 39730 40940
rect 43695 40907 44325 41027
rect 50454 41131 51454 41251
rect 50454 40875 51454 40995
rect 33671 40259 34671 40379
rect 33671 40003 34671 40123
rect 37896 40314 38556 40434
rect 37896 40090 38556 40210
rect 39598 40314 39730 40434
rect 43695 40227 44325 40347
rect 50454 40259 51454 40379
rect 43695 40003 44325 40123
rect 50454 40003 51454 40123
rect 33671 39779 34671 39899
rect 33671 39555 34671 39675
rect 39727 39779 40167 39899
rect 43695 39790 44325 39910
rect 39727 39555 40167 39675
rect 50454 39779 51454 39899
rect 43695 39544 44325 39664
rect 33671 39331 34671 39451
rect 50454 39555 51454 39675
rect 33671 39075 34671 39195
rect 37896 39244 38556 39364
rect 43695 39331 44325 39451
rect 37896 39020 38556 39140
rect 39598 39020 39730 39140
rect 43695 39107 44325 39227
rect 50454 39331 51454 39451
rect 50454 39075 51454 39195
rect 33671 38459 34671 38579
rect 33671 38203 34671 38323
rect 37896 38514 38556 38634
rect 37896 38290 38556 38410
rect 39598 38514 39730 38634
rect 43695 38427 44325 38547
rect 50454 38459 51454 38579
rect 43695 38203 44325 38323
rect 50454 38203 51454 38323
rect 33671 37979 34671 38099
rect 33671 37755 34671 37875
rect 39727 37979 40167 38099
rect 43695 37990 44325 38110
rect 39727 37755 40167 37875
rect 50454 37979 51454 38099
rect 43695 37744 44325 37864
rect 33671 37531 34671 37651
rect 50454 37755 51454 37875
rect 33671 37275 34671 37395
rect 37896 37444 38556 37564
rect 43695 37531 44325 37651
rect 37896 37220 38556 37340
rect 39598 37220 39730 37340
rect 43695 37307 44325 37427
rect 50454 37531 51454 37651
rect 50454 37275 51454 37395
rect 33671 36659 34671 36779
rect 33671 36403 34671 36523
rect 37896 36714 38556 36834
rect 37896 36490 38556 36610
rect 39598 36714 39730 36834
rect 43695 36627 44325 36747
rect 50454 36659 51454 36779
rect 43695 36403 44325 36523
rect 50454 36403 51454 36523
rect 33671 36179 34671 36299
rect 39727 36179 40167 36299
rect 43695 36190 44325 36310
rect 50454 36179 51454 36299
<< mvpmos >>
rect 29274 64983 30373 65771
rect 35396 65623 37922 65743
rect 35396 65399 37922 65519
rect 38363 65399 39681 65519
rect 42663 65399 43981 65519
rect 45333 65399 46651 65519
rect 47101 65623 49627 65743
rect 47101 65399 49627 65519
rect 29274 64083 30373 64871
rect 31336 64755 33336 64875
rect 31336 64531 33336 64651
rect 31336 64307 33336 64427
rect 44799 64755 45323 64875
rect 51789 64755 53789 64875
rect 54750 64983 55849 65771
rect 35260 64444 36360 64564
rect 35260 64220 36360 64340
rect 36841 64444 37501 64564
rect 44799 64531 45323 64651
rect 36841 64220 37501 64340
rect 39008 64220 39326 64340
rect 44799 64307 45323 64427
rect 48765 64444 49865 64564
rect 48765 64220 49865 64340
rect 51789 64531 53789 64651
rect 51789 64307 53789 64427
rect 29274 63183 30373 63971
rect 54750 64083 55849 64871
rect 31336 63627 33336 63747
rect 31336 63403 33336 63523
rect 29274 62283 30373 63071
rect 31336 63179 33336 63299
rect 35260 63714 36360 63834
rect 35260 63490 36360 63610
rect 36841 63714 37501 63834
rect 36841 63490 37501 63610
rect 39008 63714 39326 63834
rect 44799 63627 45323 63747
rect 48765 63714 49865 63834
rect 44799 63403 45323 63523
rect 48765 63490 49865 63610
rect 31336 62955 33336 63075
rect 31336 62731 33336 62851
rect 31336 62507 33336 62627
rect 44799 63179 45323 63299
rect 51789 63627 53789 63747
rect 51789 63403 53789 63523
rect 51789 63179 53789 63299
rect 44799 62955 45323 63075
rect 51789 62955 53789 63075
rect 54750 63183 55849 63971
rect 35260 62644 36360 62764
rect 35260 62420 36360 62540
rect 36841 62644 37501 62764
rect 44799 62731 45323 62851
rect 36841 62420 37501 62540
rect 39008 62420 39326 62540
rect 44799 62507 45323 62627
rect 48765 62644 49865 62764
rect 48765 62420 49865 62540
rect 51789 62731 53789 62851
rect 51789 62507 53789 62627
rect 29274 61383 30373 62171
rect 54750 62283 55849 63071
rect 31336 61827 33336 61947
rect 31336 61603 33336 61723
rect 29274 60483 30373 61271
rect 31336 61379 33336 61499
rect 35260 61914 36360 62034
rect 35260 61690 36360 61810
rect 36841 61914 37501 62034
rect 36841 61690 37501 61810
rect 39008 61914 39326 62034
rect 44799 61827 45323 61947
rect 48765 61914 49865 62034
rect 44799 61603 45323 61723
rect 48765 61690 49865 61810
rect 31336 61155 33336 61275
rect 31336 60931 33336 61051
rect 31336 60707 33336 60827
rect 44799 61379 45323 61499
rect 51789 61827 53789 61947
rect 51789 61603 53789 61723
rect 51789 61379 53789 61499
rect 44799 61155 45323 61275
rect 51789 61155 53789 61275
rect 54750 61383 55849 62171
rect 35260 60844 36360 60964
rect 35260 60620 36360 60740
rect 36841 60844 37501 60964
rect 44799 60931 45323 61051
rect 36841 60620 37501 60740
rect 39008 60620 39326 60740
rect 44799 60707 45323 60827
rect 48765 60844 49865 60964
rect 48765 60620 49865 60740
rect 51789 60931 53789 61051
rect 51789 60707 53789 60827
rect 29274 59583 30373 60371
rect 54750 60483 55849 61271
rect 31336 60027 33336 60147
rect 31336 59803 33336 59923
rect 29274 58683 30373 59471
rect 31336 59579 33336 59699
rect 35260 60114 36360 60234
rect 35260 59890 36360 60010
rect 36841 60114 37501 60234
rect 36841 59890 37501 60010
rect 39008 60114 39326 60234
rect 44799 60027 45323 60147
rect 48765 60114 49865 60234
rect 44799 59803 45323 59923
rect 48765 59890 49865 60010
rect 31336 59355 33336 59475
rect 31336 59131 33336 59251
rect 31336 58907 33336 59027
rect 44799 59579 45323 59699
rect 51789 60027 53789 60147
rect 51789 59803 53789 59923
rect 51789 59579 53789 59699
rect 44799 59355 45323 59475
rect 51789 59355 53789 59475
rect 54750 59583 55849 60371
rect 35260 59044 36360 59164
rect 35260 58820 36360 58940
rect 36841 59044 37501 59164
rect 44799 59131 45323 59251
rect 36841 58820 37501 58940
rect 39008 58820 39326 58940
rect 44799 58907 45323 59027
rect 48765 59044 49865 59164
rect 48765 58820 49865 58940
rect 51789 59131 53789 59251
rect 51789 58907 53789 59027
rect 29274 57783 30373 58571
rect 54750 58683 55849 59471
rect 31336 58227 33336 58347
rect 31336 58003 33336 58123
rect 29274 56883 30373 57671
rect 31336 57779 33336 57899
rect 35260 58314 36360 58434
rect 35260 58090 36360 58210
rect 36841 58314 37501 58434
rect 36841 58090 37501 58210
rect 39008 58314 39326 58434
rect 44799 58227 45323 58347
rect 48765 58314 49865 58434
rect 44799 58003 45323 58123
rect 48765 58090 49865 58210
rect 31336 57555 33336 57675
rect 31336 57331 33336 57451
rect 31336 57107 33336 57227
rect 44799 57779 45323 57899
rect 51789 58227 53789 58347
rect 51789 58003 53789 58123
rect 51789 57779 53789 57899
rect 44799 57555 45323 57675
rect 51789 57555 53789 57675
rect 54750 57783 55849 58571
rect 35260 57244 36360 57364
rect 35260 57020 36360 57140
rect 36841 57244 37501 57364
rect 44799 57331 45323 57451
rect 36841 57020 37501 57140
rect 39008 57020 39326 57140
rect 44799 57107 45323 57227
rect 48765 57244 49865 57364
rect 48765 57020 49865 57140
rect 51789 57331 53789 57451
rect 51789 57107 53789 57227
rect 29274 55983 30373 56771
rect 54750 56883 55849 57671
rect 31336 56427 33336 56547
rect 31336 56203 33336 56323
rect 29274 55083 30373 55871
rect 31336 55979 33336 56099
rect 35260 56514 36360 56634
rect 35260 56290 36360 56410
rect 36841 56514 37501 56634
rect 36841 56290 37501 56410
rect 39008 56514 39326 56634
rect 44799 56427 45323 56547
rect 48765 56514 49865 56634
rect 44799 56203 45323 56323
rect 48765 56290 49865 56410
rect 31336 55755 33336 55875
rect 31336 55531 33336 55651
rect 31336 55307 33336 55427
rect 44799 55979 45323 56099
rect 51789 56427 53789 56547
rect 51789 56203 53789 56323
rect 51789 55979 53789 56099
rect 44799 55755 45323 55875
rect 51789 55755 53789 55875
rect 54750 55983 55849 56771
rect 35260 55444 36360 55564
rect 35260 55220 36360 55340
rect 36841 55444 37501 55564
rect 44799 55531 45323 55651
rect 36841 55220 37501 55340
rect 39008 55220 39326 55340
rect 44799 55307 45323 55427
rect 48765 55444 49865 55564
rect 48765 55220 49865 55340
rect 51789 55531 53789 55651
rect 51789 55307 53789 55427
rect 29274 54183 30373 54971
rect 54750 55083 55849 55871
rect 31336 54627 33336 54747
rect 31336 54403 33336 54523
rect 29274 53283 30373 54071
rect 31336 54179 33336 54299
rect 35260 54714 36360 54834
rect 35260 54490 36360 54610
rect 36841 54714 37501 54834
rect 36841 54490 37501 54610
rect 39008 54714 39326 54834
rect 44799 54627 45323 54747
rect 48765 54714 49865 54834
rect 44799 54403 45323 54523
rect 48765 54490 49865 54610
rect 31336 53955 33336 54075
rect 31336 53731 33336 53851
rect 31336 53507 33336 53627
rect 44799 54179 45323 54299
rect 51789 54627 53789 54747
rect 51789 54403 53789 54523
rect 51789 54179 53789 54299
rect 44799 53955 45323 54075
rect 51789 53955 53789 54075
rect 54750 54183 55849 54971
rect 35260 53644 36360 53764
rect 35260 53420 36360 53540
rect 36841 53644 37501 53764
rect 44799 53731 45323 53851
rect 36841 53420 37501 53540
rect 39008 53420 39326 53540
rect 44799 53507 45323 53627
rect 48765 53644 49865 53764
rect 48765 53420 49865 53540
rect 51789 53731 53789 53851
rect 51789 53507 53789 53627
rect 29274 52383 30373 53171
rect 54750 53283 55849 54071
rect 31336 52827 33336 52947
rect 31336 52603 33336 52723
rect 29274 51483 30373 52271
rect 31336 52379 33336 52499
rect 35260 52914 36360 53034
rect 35260 52690 36360 52810
rect 36841 52914 37501 53034
rect 36841 52690 37501 52810
rect 39008 52914 39326 53034
rect 44799 52827 45323 52947
rect 48765 52914 49865 53034
rect 44799 52603 45323 52723
rect 48765 52690 49865 52810
rect 31336 52155 33336 52275
rect 31336 51931 33336 52051
rect 31336 51707 33336 51827
rect 44799 52379 45323 52499
rect 51789 52827 53789 52947
rect 51789 52603 53789 52723
rect 51789 52379 53789 52499
rect 44799 52155 45323 52275
rect 51789 52155 53789 52275
rect 54750 52383 55849 53171
rect 35260 51844 36360 51964
rect 35260 51620 36360 51740
rect 36841 51844 37501 51964
rect 44799 51931 45323 52051
rect 36841 51620 37501 51740
rect 39008 51620 39326 51740
rect 44799 51707 45323 51827
rect 48765 51844 49865 51964
rect 48765 51620 49865 51740
rect 51789 51931 53789 52051
rect 51789 51707 53789 51827
rect 29274 50583 30373 51371
rect 54750 51483 55849 52271
rect 31336 51027 33336 51147
rect 31336 50803 33336 50923
rect 29274 49683 30373 50471
rect 31336 50579 33336 50699
rect 35260 51114 36360 51234
rect 35260 50890 36360 51010
rect 36841 51114 37501 51234
rect 36841 50890 37501 51010
rect 39008 51114 39326 51234
rect 44799 51027 45323 51147
rect 48765 51114 49865 51234
rect 44799 50803 45323 50923
rect 48765 50890 49865 51010
rect 31336 50355 33336 50475
rect 31336 50131 33336 50251
rect 31336 49907 33336 50027
rect 44799 50579 45323 50699
rect 51789 51027 53789 51147
rect 51789 50803 53789 50923
rect 51789 50579 53789 50699
rect 44799 50355 45323 50475
rect 51789 50355 53789 50475
rect 54750 50583 55849 51371
rect 35260 50044 36360 50164
rect 35260 49820 36360 49940
rect 36841 50044 37501 50164
rect 44799 50131 45323 50251
rect 36841 49820 37501 49940
rect 39008 49820 39326 49940
rect 44799 49907 45323 50027
rect 48765 50044 49865 50164
rect 48765 49820 49865 49940
rect 51789 50131 53789 50251
rect 51789 49907 53789 50027
rect 29274 48783 30373 49571
rect 54750 49683 55849 50471
rect 31336 49227 33336 49347
rect 31336 49003 33336 49123
rect 29274 47883 30373 48671
rect 31336 48779 33336 48899
rect 35260 49314 36360 49434
rect 35260 49090 36360 49210
rect 36841 49314 37501 49434
rect 36841 49090 37501 49210
rect 39008 49314 39326 49434
rect 44799 49227 45323 49347
rect 48765 49314 49865 49434
rect 44799 49003 45323 49123
rect 48765 49090 49865 49210
rect 31336 48555 33336 48675
rect 31336 48331 33336 48451
rect 31336 48107 33336 48227
rect 44799 48779 45323 48899
rect 51789 49227 53789 49347
rect 51789 49003 53789 49123
rect 51789 48779 53789 48899
rect 44799 48555 45323 48675
rect 51789 48555 53789 48675
rect 54750 48783 55849 49571
rect 35260 48244 36360 48364
rect 35260 48020 36360 48140
rect 36841 48244 37501 48364
rect 44799 48331 45323 48451
rect 36841 48020 37501 48140
rect 39008 48020 39326 48140
rect 44799 48107 45323 48227
rect 48765 48244 49865 48364
rect 48765 48020 49865 48140
rect 51789 48331 53789 48451
rect 51789 48107 53789 48227
rect 29274 46983 30373 47771
rect 54750 47883 55849 48671
rect 31336 47427 33336 47547
rect 31336 47203 33336 47323
rect 29274 46083 30373 46871
rect 31336 46979 33336 47099
rect 35260 47514 36360 47634
rect 35260 47290 36360 47410
rect 36841 47514 37501 47634
rect 36841 47290 37501 47410
rect 39008 47514 39326 47634
rect 44799 47427 45323 47547
rect 48765 47514 49865 47634
rect 44799 47203 45323 47323
rect 48765 47290 49865 47410
rect 31336 46755 33336 46875
rect 31336 46531 33336 46651
rect 31336 46307 33336 46427
rect 44799 46979 45323 47099
rect 51789 47427 53789 47547
rect 51789 47203 53789 47323
rect 51789 46979 53789 47099
rect 44799 46755 45323 46875
rect 51789 46755 53789 46875
rect 54750 46983 55849 47771
rect 35260 46444 36360 46564
rect 35260 46220 36360 46340
rect 36841 46444 37501 46564
rect 44799 46531 45323 46651
rect 36841 46220 37501 46340
rect 39008 46220 39326 46340
rect 44799 46307 45323 46427
rect 48765 46444 49865 46564
rect 48765 46220 49865 46340
rect 51789 46531 53789 46651
rect 51789 46307 53789 46427
rect 29274 45183 30373 45971
rect 54750 46083 55849 46871
rect 31336 45627 33336 45747
rect 31336 45403 33336 45523
rect 29274 44283 30373 45071
rect 31336 45179 33336 45299
rect 35260 45714 36360 45834
rect 35260 45490 36360 45610
rect 36841 45714 37501 45834
rect 36841 45490 37501 45610
rect 39008 45714 39326 45834
rect 44799 45627 45323 45747
rect 48765 45714 49865 45834
rect 44799 45403 45323 45523
rect 48765 45490 49865 45610
rect 31336 44955 33336 45075
rect 31336 44731 33336 44851
rect 31336 44507 33336 44627
rect 44799 45179 45323 45299
rect 51789 45627 53789 45747
rect 51789 45403 53789 45523
rect 51789 45179 53789 45299
rect 44799 44955 45323 45075
rect 51789 44955 53789 45075
rect 54750 45183 55849 45971
rect 35260 44644 36360 44764
rect 35260 44420 36360 44540
rect 36841 44644 37501 44764
rect 44799 44731 45323 44851
rect 36841 44420 37501 44540
rect 39008 44420 39326 44540
rect 44799 44507 45323 44627
rect 48765 44644 49865 44764
rect 48765 44420 49865 44540
rect 51789 44731 53789 44851
rect 51789 44507 53789 44627
rect 29274 43383 30373 44171
rect 54750 44283 55849 45071
rect 31336 43827 33336 43947
rect 31336 43603 33336 43723
rect 29274 42483 30373 43271
rect 31336 43379 33336 43499
rect 35260 43914 36360 44034
rect 35260 43690 36360 43810
rect 36841 43914 37501 44034
rect 36841 43690 37501 43810
rect 39008 43914 39326 44034
rect 44799 43827 45323 43947
rect 48765 43914 49865 44034
rect 44799 43603 45323 43723
rect 48765 43690 49865 43810
rect 31336 43155 33336 43275
rect 31336 42931 33336 43051
rect 31336 42707 33336 42827
rect 44799 43379 45323 43499
rect 51789 43827 53789 43947
rect 51789 43603 53789 43723
rect 51789 43379 53789 43499
rect 44799 43155 45323 43275
rect 51789 43155 53789 43275
rect 54750 43383 55849 44171
rect 35260 42844 36360 42964
rect 35260 42620 36360 42740
rect 36841 42844 37501 42964
rect 44799 42931 45323 43051
rect 36841 42620 37501 42740
rect 39008 42620 39326 42740
rect 44799 42707 45323 42827
rect 48765 42844 49865 42964
rect 48765 42620 49865 42740
rect 51789 42931 53789 43051
rect 51789 42707 53789 42827
rect 29274 41583 30373 42371
rect 54750 42483 55849 43271
rect 31336 42027 33336 42147
rect 31336 41803 33336 41923
rect 29274 40683 30373 41471
rect 31336 41579 33336 41699
rect 35260 42114 36360 42234
rect 35260 41890 36360 42010
rect 36841 42114 37501 42234
rect 36841 41890 37501 42010
rect 39008 42114 39326 42234
rect 44799 42027 45323 42147
rect 48765 42114 49865 42234
rect 44799 41803 45323 41923
rect 48765 41890 49865 42010
rect 31336 41355 33336 41475
rect 31336 41131 33336 41251
rect 31336 40907 33336 41027
rect 44799 41579 45323 41699
rect 51789 42027 53789 42147
rect 51789 41803 53789 41923
rect 51789 41579 53789 41699
rect 44799 41355 45323 41475
rect 51789 41355 53789 41475
rect 54750 41583 55849 42371
rect 35260 41044 36360 41164
rect 35260 40820 36360 40940
rect 36841 41044 37501 41164
rect 44799 41131 45323 41251
rect 36841 40820 37501 40940
rect 39008 40820 39326 40940
rect 44799 40907 45323 41027
rect 48765 41044 49865 41164
rect 48765 40820 49865 40940
rect 51789 41131 53789 41251
rect 51789 40907 53789 41027
rect 29274 39783 30373 40571
rect 54750 40683 55849 41471
rect 31336 40227 33336 40347
rect 31336 40003 33336 40123
rect 29274 38883 30373 39671
rect 31336 39779 33336 39899
rect 35260 40314 36360 40434
rect 35260 40090 36360 40210
rect 36841 40314 37501 40434
rect 36841 40090 37501 40210
rect 39008 40314 39326 40434
rect 44799 40227 45323 40347
rect 48765 40314 49865 40434
rect 44799 40003 45323 40123
rect 48765 40090 49865 40210
rect 31336 39555 33336 39675
rect 31336 39331 33336 39451
rect 31336 39107 33336 39227
rect 44799 39779 45323 39899
rect 51789 40227 53789 40347
rect 51789 40003 53789 40123
rect 51789 39779 53789 39899
rect 44799 39555 45323 39675
rect 51789 39555 53789 39675
rect 54750 39783 55849 40571
rect 35260 39244 36360 39364
rect 35260 39020 36360 39140
rect 36841 39244 37501 39364
rect 44799 39331 45323 39451
rect 36841 39020 37501 39140
rect 39008 39020 39326 39140
rect 44799 39107 45323 39227
rect 48765 39244 49865 39364
rect 48765 39020 49865 39140
rect 51789 39331 53789 39451
rect 51789 39107 53789 39227
rect 29274 37983 30373 38771
rect 54750 38883 55849 39671
rect 31336 38427 33336 38547
rect 31336 38203 33336 38323
rect 29274 37083 30373 37871
rect 31336 37979 33336 38099
rect 35260 38514 36360 38634
rect 35260 38290 36360 38410
rect 36841 38514 37501 38634
rect 36841 38290 37501 38410
rect 39008 38514 39326 38634
rect 44799 38427 45323 38547
rect 48765 38514 49865 38634
rect 44799 38203 45323 38323
rect 48765 38290 49865 38410
rect 31336 37755 33336 37875
rect 31336 37531 33336 37651
rect 31336 37307 33336 37427
rect 44799 37979 45323 38099
rect 51789 38427 53789 38547
rect 51789 38203 53789 38323
rect 51789 37979 53789 38099
rect 44799 37755 45323 37875
rect 51789 37755 53789 37875
rect 54750 37983 55849 38771
rect 35260 37444 36360 37564
rect 35260 37220 36360 37340
rect 36841 37444 37501 37564
rect 44799 37531 45323 37651
rect 36841 37220 37501 37340
rect 39008 37220 39326 37340
rect 44799 37307 45323 37427
rect 48765 37444 49865 37564
rect 48765 37220 49865 37340
rect 51789 37531 53789 37651
rect 51789 37307 53789 37427
rect 29274 36183 30373 36971
rect 54750 37083 55849 37871
rect 31336 36627 33336 36747
rect 31336 36403 33336 36523
rect 31336 36179 33336 36299
rect 35260 36714 36360 36834
rect 35260 36490 36360 36610
rect 36841 36714 37501 36834
rect 36841 36490 37501 36610
rect 39008 36714 39326 36834
rect 44799 36627 45323 36747
rect 48765 36714 49865 36834
rect 44799 36403 45323 36523
rect 48765 36490 49865 36610
rect 44799 36179 45323 36299
rect 51789 36627 53789 36747
rect 51789 36403 53789 36523
rect 51789 36179 53789 36299
rect 54750 36183 55849 36971
<< mvndiff >>
rect 33001 65594 35023 65607
rect 33001 65548 33014 65594
rect 33774 65548 33831 65594
rect 33877 65548 33934 65594
rect 33980 65548 34037 65594
rect 34083 65548 34140 65594
rect 34186 65548 34243 65594
rect 34289 65548 34346 65594
rect 34392 65548 34449 65594
rect 34495 65548 34552 65594
rect 34598 65548 34655 65594
rect 34701 65548 34758 65594
rect 34804 65548 34861 65594
rect 34907 65548 34964 65594
rect 35010 65548 35023 65594
rect 33001 65519 35023 65548
rect 40062 65594 40590 65607
rect 40062 65548 40075 65594
rect 40121 65548 40189 65594
rect 40235 65548 40303 65594
rect 40349 65548 40417 65594
rect 40463 65548 40531 65594
rect 40577 65548 40590 65594
rect 40963 65595 42281 65608
rect 40062 65519 40590 65548
rect 40963 65549 40976 65595
rect 41022 65549 41079 65595
rect 41125 65549 41182 65595
rect 41228 65549 41286 65595
rect 41332 65549 41390 65595
rect 41436 65549 41494 65595
rect 41540 65549 41598 65595
rect 41644 65549 41702 65595
rect 41748 65549 41806 65595
rect 41852 65549 41910 65595
rect 41956 65549 42014 65595
rect 42060 65549 42118 65595
rect 42164 65549 42222 65595
rect 42268 65549 42281 65595
rect 40963 65520 42281 65549
rect 33001 65370 35023 65399
rect 33001 65324 33014 65370
rect 33774 65324 33831 65370
rect 33877 65324 33934 65370
rect 33980 65324 34037 65370
rect 34083 65324 34140 65370
rect 34186 65324 34243 65370
rect 34289 65324 34346 65370
rect 34392 65324 34449 65370
rect 34495 65324 34552 65370
rect 34598 65324 34655 65370
rect 34701 65324 34758 65370
rect 34804 65324 34861 65370
rect 34907 65324 34964 65370
rect 35010 65324 35023 65370
rect 33001 65311 35023 65324
rect 40062 65370 40590 65399
rect 40062 65324 40075 65370
rect 40121 65324 40189 65370
rect 40235 65324 40303 65370
rect 40349 65324 40417 65370
rect 40463 65324 40531 65370
rect 40577 65324 40590 65370
rect 40062 65311 40590 65324
rect 40963 65371 42281 65400
rect 44432 65594 44960 65607
rect 44432 65548 44445 65594
rect 44491 65548 44559 65594
rect 44605 65548 44673 65594
rect 44719 65548 44787 65594
rect 44833 65548 44901 65594
rect 44947 65548 44960 65594
rect 44432 65519 44960 65548
rect 50001 65594 52023 65607
rect 50001 65548 50014 65594
rect 50774 65548 50831 65594
rect 50877 65548 50934 65594
rect 50980 65548 51037 65594
rect 51083 65548 51140 65594
rect 51186 65548 51243 65594
rect 51289 65548 51346 65594
rect 51392 65548 51449 65594
rect 51495 65548 51552 65594
rect 51598 65548 51655 65594
rect 51701 65548 51758 65594
rect 51804 65548 51861 65594
rect 51907 65548 51964 65594
rect 52010 65548 52023 65594
rect 50001 65519 52023 65548
rect 40963 65325 40976 65371
rect 41022 65325 41079 65371
rect 41125 65325 41182 65371
rect 41228 65325 41286 65371
rect 41332 65325 41390 65371
rect 41436 65325 41494 65371
rect 41540 65325 41598 65371
rect 41644 65325 41702 65371
rect 41748 65325 41806 65371
rect 41852 65325 41910 65371
rect 41956 65325 42014 65371
rect 42060 65325 42118 65371
rect 42164 65325 42222 65371
rect 42268 65325 42281 65371
rect 40963 65312 42281 65325
rect 44432 65370 44960 65399
rect 44432 65324 44445 65370
rect 44491 65324 44559 65370
rect 44605 65324 44673 65370
rect 44719 65324 44787 65370
rect 44833 65324 44901 65370
rect 44947 65324 44960 65370
rect 44432 65311 44960 65324
rect 50001 65370 52023 65399
rect 50001 65324 50014 65370
rect 50774 65324 50831 65370
rect 50877 65324 50934 65370
rect 50980 65324 51037 65370
rect 51083 65324 51140 65370
rect 51186 65324 51243 65370
rect 51289 65324 51346 65370
rect 51392 65324 51449 65370
rect 51495 65324 51552 65370
rect 51598 65324 51655 65370
rect 51701 65324 51758 65370
rect 51804 65324 51861 65370
rect 51907 65324 51964 65370
rect 52010 65324 52023 65370
rect 50001 65311 52023 65324
rect 33671 64950 34671 64963
rect 33671 64904 33684 64950
rect 33730 64904 33787 64950
rect 33833 64904 33890 64950
rect 33936 64904 33993 64950
rect 34039 64904 34096 64950
rect 34142 64904 34199 64950
rect 34245 64904 34302 64950
rect 34348 64904 34405 64950
rect 34451 64904 34508 64950
rect 34554 64904 34612 64950
rect 34658 64904 34671 64950
rect 33671 64875 34671 64904
rect 39727 64950 40167 64963
rect 39727 64904 39740 64950
rect 39786 64904 39862 64950
rect 39908 64904 39985 64950
rect 40031 64904 40108 64950
rect 40154 64904 40167 64950
rect 39727 64875 40167 64904
rect 43695 64950 44325 64996
rect 43695 64904 43739 64950
rect 43785 64904 43906 64950
rect 43952 64904 44071 64950
rect 44117 64904 44236 64950
rect 44282 64904 44325 64950
rect 43695 64864 44325 64904
rect 33671 64726 34671 64755
rect 33671 64680 33684 64726
rect 33730 64680 33787 64726
rect 33833 64680 33890 64726
rect 33936 64680 33993 64726
rect 34039 64680 34096 64726
rect 34142 64680 34199 64726
rect 34245 64680 34302 64726
rect 34348 64680 34405 64726
rect 34451 64680 34508 64726
rect 34554 64680 34612 64726
rect 34658 64680 34671 64726
rect 33671 64651 34671 64680
rect 39727 64726 40167 64755
rect 39727 64680 39740 64726
rect 39786 64680 39862 64726
rect 39908 64680 39985 64726
rect 40031 64680 40108 64726
rect 40154 64680 40167 64726
rect 39727 64667 40167 64680
rect 50454 64950 51454 64963
rect 50454 64904 50467 64950
rect 50513 64904 50571 64950
rect 50617 64904 50674 64950
rect 50720 64904 50777 64950
rect 50823 64904 50880 64950
rect 50926 64904 50983 64950
rect 51029 64904 51086 64950
rect 51132 64904 51189 64950
rect 51235 64904 51292 64950
rect 51338 64904 51395 64950
rect 51441 64904 51454 64950
rect 50454 64875 51454 64904
rect 37896 64639 38556 64652
rect 43695 64651 44325 64744
rect 50454 64726 51454 64755
rect 50454 64680 50467 64726
rect 50513 64680 50571 64726
rect 50617 64680 50674 64726
rect 50720 64680 50777 64726
rect 50823 64680 50880 64726
rect 50926 64680 50983 64726
rect 51029 64680 51086 64726
rect 51132 64680 51189 64726
rect 51235 64680 51292 64726
rect 51338 64680 51395 64726
rect 51441 64680 51454 64726
rect 37896 64593 37909 64639
rect 37955 64593 38026 64639
rect 38072 64593 38143 64639
rect 38189 64593 38261 64639
rect 38307 64593 38379 64639
rect 38425 64593 38497 64639
rect 38543 64593 38556 64639
rect 37896 64564 38556 64593
rect 33671 64502 34671 64531
rect 33671 64456 33684 64502
rect 33730 64456 33787 64502
rect 33833 64456 33890 64502
rect 33936 64456 33993 64502
rect 34039 64456 34096 64502
rect 34142 64456 34199 64502
rect 34245 64456 34302 64502
rect 34348 64456 34405 64502
rect 34451 64456 34508 64502
rect 34554 64456 34612 64502
rect 34658 64456 34671 64502
rect 33671 64395 34671 64456
rect 33671 64243 34671 64275
rect 33671 64197 33816 64243
rect 33862 64197 34002 64243
rect 34048 64197 34189 64243
rect 34235 64197 34376 64243
rect 34422 64197 34562 64243
rect 34608 64197 34671 64243
rect 50454 64651 51454 64680
rect 37896 64415 38556 64444
rect 37896 64369 37909 64415
rect 37955 64369 38026 64415
rect 38072 64369 38143 64415
rect 38189 64369 38261 64415
rect 38307 64369 38379 64415
rect 38425 64369 38497 64415
rect 38543 64369 38556 64415
rect 37896 64340 38556 64369
rect 39598 64415 39730 64428
rect 43695 64427 44325 64531
rect 39598 64369 39641 64415
rect 39687 64369 39730 64415
rect 39598 64340 39730 64369
rect 50454 64502 51454 64531
rect 50454 64456 50467 64502
rect 50513 64456 50571 64502
rect 50617 64456 50674 64502
rect 50720 64456 50777 64502
rect 50823 64456 50880 64502
rect 50926 64456 50983 64502
rect 51029 64456 51086 64502
rect 51132 64456 51189 64502
rect 51235 64456 51292 64502
rect 51338 64456 51395 64502
rect 51441 64456 51454 64502
rect 50454 64395 51454 64456
rect 43695 64257 44325 64307
rect 33671 64151 34671 64197
rect 37896 64191 38556 64220
rect 37896 64145 37909 64191
rect 37955 64145 38026 64191
rect 38072 64145 38143 64191
rect 38189 64145 38261 64191
rect 38307 64145 38379 64191
rect 38425 64145 38497 64191
rect 38543 64145 38556 64191
rect 37896 64132 38556 64145
rect 39598 64191 39730 64220
rect 39598 64145 39641 64191
rect 39687 64145 39730 64191
rect 43695 64211 43739 64257
rect 43785 64211 43906 64257
rect 43952 64211 44071 64257
rect 44117 64211 44236 64257
rect 44282 64211 44325 64257
rect 50454 64243 51454 64275
rect 43695 64164 44325 64211
rect 39598 64132 39730 64145
rect 50454 64197 50516 64243
rect 50562 64197 50703 64243
rect 50749 64197 50890 64243
rect 50936 64197 51076 64243
rect 51122 64197 51263 64243
rect 51309 64197 51454 64243
rect 50454 64151 51454 64197
rect 33671 63857 34671 63903
rect 33671 63811 33816 63857
rect 33862 63811 34002 63857
rect 34048 63811 34189 63857
rect 34235 63811 34376 63857
rect 34422 63811 34562 63857
rect 34608 63811 34671 63857
rect 37896 63909 38556 63922
rect 37896 63863 37909 63909
rect 37955 63863 38026 63909
rect 38072 63863 38143 63909
rect 38189 63863 38261 63909
rect 38307 63863 38379 63909
rect 38425 63863 38497 63909
rect 38543 63863 38556 63909
rect 37896 63834 38556 63863
rect 39598 63909 39730 63922
rect 39598 63863 39641 63909
rect 39687 63863 39730 63909
rect 39598 63834 39730 63863
rect 43695 63843 44325 63890
rect 33671 63779 34671 63811
rect 33671 63598 34671 63659
rect 33671 63552 33684 63598
rect 33730 63552 33787 63598
rect 33833 63552 33890 63598
rect 33936 63552 33993 63598
rect 34039 63552 34096 63598
rect 34142 63552 34199 63598
rect 34245 63552 34302 63598
rect 34348 63552 34405 63598
rect 34451 63552 34508 63598
rect 34554 63552 34612 63598
rect 34658 63552 34671 63598
rect 33671 63523 34671 63552
rect 37896 63685 38556 63714
rect 37896 63639 37909 63685
rect 37955 63639 38026 63685
rect 38072 63639 38143 63685
rect 38189 63639 38261 63685
rect 38307 63639 38379 63685
rect 38425 63639 38497 63685
rect 38543 63639 38556 63685
rect 37896 63610 38556 63639
rect 43695 63797 43739 63843
rect 43785 63797 43906 63843
rect 43952 63797 44071 63843
rect 44117 63797 44236 63843
rect 44282 63797 44325 63843
rect 43695 63747 44325 63797
rect 50454 63857 51454 63903
rect 39598 63685 39730 63714
rect 39598 63639 39641 63685
rect 39687 63639 39730 63685
rect 39598 63626 39730 63639
rect 50454 63811 50516 63857
rect 50562 63811 50703 63857
rect 50749 63811 50890 63857
rect 50936 63811 51076 63857
rect 51122 63811 51263 63857
rect 51309 63811 51454 63857
rect 50454 63779 51454 63811
rect 43695 63523 44325 63627
rect 33671 63374 34671 63403
rect 37896 63461 38556 63490
rect 37896 63415 37909 63461
rect 37955 63415 38026 63461
rect 38072 63415 38143 63461
rect 38189 63415 38261 63461
rect 38307 63415 38379 63461
rect 38425 63415 38497 63461
rect 38543 63415 38556 63461
rect 37896 63402 38556 63415
rect 50454 63598 51454 63659
rect 50454 63552 50467 63598
rect 50513 63552 50571 63598
rect 50617 63552 50674 63598
rect 50720 63552 50777 63598
rect 50823 63552 50880 63598
rect 50926 63552 50983 63598
rect 51029 63552 51086 63598
rect 51132 63552 51189 63598
rect 51235 63552 51292 63598
rect 51338 63552 51395 63598
rect 51441 63552 51454 63598
rect 50454 63523 51454 63552
rect 33671 63328 33684 63374
rect 33730 63328 33787 63374
rect 33833 63328 33890 63374
rect 33936 63328 33993 63374
rect 34039 63328 34096 63374
rect 34142 63328 34199 63374
rect 34245 63328 34302 63374
rect 34348 63328 34405 63374
rect 34451 63328 34508 63374
rect 34554 63328 34612 63374
rect 34658 63328 34671 63374
rect 33671 63299 34671 63328
rect 39727 63374 40167 63387
rect 39727 63328 39740 63374
rect 39786 63328 39862 63374
rect 39908 63328 39985 63374
rect 40031 63328 40108 63374
rect 40154 63328 40167 63374
rect 39727 63299 40167 63328
rect 43695 63310 44325 63403
rect 50454 63374 51454 63403
rect 33671 63150 34671 63179
rect 33671 63104 33684 63150
rect 33730 63104 33787 63150
rect 33833 63104 33890 63150
rect 33936 63104 33993 63150
rect 34039 63104 34096 63150
rect 34142 63104 34199 63150
rect 34245 63104 34302 63150
rect 34348 63104 34405 63150
rect 34451 63104 34508 63150
rect 34554 63104 34612 63150
rect 34658 63104 34671 63150
rect 33671 63075 34671 63104
rect 39727 63150 40167 63179
rect 39727 63104 39740 63150
rect 39786 63104 39862 63150
rect 39908 63104 39985 63150
rect 40031 63104 40108 63150
rect 40154 63104 40167 63150
rect 39727 63075 40167 63104
rect 43695 63150 44325 63190
rect 50454 63328 50467 63374
rect 50513 63328 50571 63374
rect 50617 63328 50674 63374
rect 50720 63328 50777 63374
rect 50823 63328 50880 63374
rect 50926 63328 50983 63374
rect 51029 63328 51086 63374
rect 51132 63328 51189 63374
rect 51235 63328 51292 63374
rect 51338 63328 51395 63374
rect 51441 63328 51454 63374
rect 50454 63299 51454 63328
rect 43695 63104 43739 63150
rect 43785 63104 43906 63150
rect 43952 63104 44071 63150
rect 44117 63104 44236 63150
rect 44282 63104 44325 63150
rect 43695 63064 44325 63104
rect 33671 62926 34671 62955
rect 33671 62880 33684 62926
rect 33730 62880 33787 62926
rect 33833 62880 33890 62926
rect 33936 62880 33993 62926
rect 34039 62880 34096 62926
rect 34142 62880 34199 62926
rect 34245 62880 34302 62926
rect 34348 62880 34405 62926
rect 34451 62880 34508 62926
rect 34554 62880 34612 62926
rect 34658 62880 34671 62926
rect 33671 62851 34671 62880
rect 39727 62926 40167 62955
rect 39727 62880 39740 62926
rect 39786 62880 39862 62926
rect 39908 62880 39985 62926
rect 40031 62880 40108 62926
rect 40154 62880 40167 62926
rect 39727 62867 40167 62880
rect 50454 63150 51454 63179
rect 50454 63104 50467 63150
rect 50513 63104 50571 63150
rect 50617 63104 50674 63150
rect 50720 63104 50777 63150
rect 50823 63104 50880 63150
rect 50926 63104 50983 63150
rect 51029 63104 51086 63150
rect 51132 63104 51189 63150
rect 51235 63104 51292 63150
rect 51338 63104 51395 63150
rect 51441 63104 51454 63150
rect 50454 63075 51454 63104
rect 37896 62839 38556 62852
rect 43695 62851 44325 62944
rect 50454 62926 51454 62955
rect 50454 62880 50467 62926
rect 50513 62880 50571 62926
rect 50617 62880 50674 62926
rect 50720 62880 50777 62926
rect 50823 62880 50880 62926
rect 50926 62880 50983 62926
rect 51029 62880 51086 62926
rect 51132 62880 51189 62926
rect 51235 62880 51292 62926
rect 51338 62880 51395 62926
rect 51441 62880 51454 62926
rect 37896 62793 37909 62839
rect 37955 62793 38026 62839
rect 38072 62793 38143 62839
rect 38189 62793 38261 62839
rect 38307 62793 38379 62839
rect 38425 62793 38497 62839
rect 38543 62793 38556 62839
rect 37896 62764 38556 62793
rect 33671 62702 34671 62731
rect 33671 62656 33684 62702
rect 33730 62656 33787 62702
rect 33833 62656 33890 62702
rect 33936 62656 33993 62702
rect 34039 62656 34096 62702
rect 34142 62656 34199 62702
rect 34245 62656 34302 62702
rect 34348 62656 34405 62702
rect 34451 62656 34508 62702
rect 34554 62656 34612 62702
rect 34658 62656 34671 62702
rect 33671 62595 34671 62656
rect 33671 62443 34671 62475
rect 33671 62397 33816 62443
rect 33862 62397 34002 62443
rect 34048 62397 34189 62443
rect 34235 62397 34376 62443
rect 34422 62397 34562 62443
rect 34608 62397 34671 62443
rect 50454 62851 51454 62880
rect 37896 62615 38556 62644
rect 37896 62569 37909 62615
rect 37955 62569 38026 62615
rect 38072 62569 38143 62615
rect 38189 62569 38261 62615
rect 38307 62569 38379 62615
rect 38425 62569 38497 62615
rect 38543 62569 38556 62615
rect 37896 62540 38556 62569
rect 39598 62615 39730 62628
rect 43695 62627 44325 62731
rect 39598 62569 39641 62615
rect 39687 62569 39730 62615
rect 39598 62540 39730 62569
rect 50454 62702 51454 62731
rect 50454 62656 50467 62702
rect 50513 62656 50571 62702
rect 50617 62656 50674 62702
rect 50720 62656 50777 62702
rect 50823 62656 50880 62702
rect 50926 62656 50983 62702
rect 51029 62656 51086 62702
rect 51132 62656 51189 62702
rect 51235 62656 51292 62702
rect 51338 62656 51395 62702
rect 51441 62656 51454 62702
rect 50454 62595 51454 62656
rect 43695 62457 44325 62507
rect 33671 62351 34671 62397
rect 37896 62391 38556 62420
rect 37896 62345 37909 62391
rect 37955 62345 38026 62391
rect 38072 62345 38143 62391
rect 38189 62345 38261 62391
rect 38307 62345 38379 62391
rect 38425 62345 38497 62391
rect 38543 62345 38556 62391
rect 37896 62332 38556 62345
rect 39598 62391 39730 62420
rect 39598 62345 39641 62391
rect 39687 62345 39730 62391
rect 43695 62411 43739 62457
rect 43785 62411 43906 62457
rect 43952 62411 44071 62457
rect 44117 62411 44236 62457
rect 44282 62411 44325 62457
rect 50454 62443 51454 62475
rect 43695 62364 44325 62411
rect 39598 62332 39730 62345
rect 50454 62397 50516 62443
rect 50562 62397 50703 62443
rect 50749 62397 50890 62443
rect 50936 62397 51076 62443
rect 51122 62397 51263 62443
rect 51309 62397 51454 62443
rect 50454 62351 51454 62397
rect 33671 62057 34671 62103
rect 33671 62011 33816 62057
rect 33862 62011 34002 62057
rect 34048 62011 34189 62057
rect 34235 62011 34376 62057
rect 34422 62011 34562 62057
rect 34608 62011 34671 62057
rect 37896 62109 38556 62122
rect 37896 62063 37909 62109
rect 37955 62063 38026 62109
rect 38072 62063 38143 62109
rect 38189 62063 38261 62109
rect 38307 62063 38379 62109
rect 38425 62063 38497 62109
rect 38543 62063 38556 62109
rect 37896 62034 38556 62063
rect 39598 62109 39730 62122
rect 39598 62063 39641 62109
rect 39687 62063 39730 62109
rect 39598 62034 39730 62063
rect 43695 62043 44325 62090
rect 33671 61979 34671 62011
rect 33671 61798 34671 61859
rect 33671 61752 33684 61798
rect 33730 61752 33787 61798
rect 33833 61752 33890 61798
rect 33936 61752 33993 61798
rect 34039 61752 34096 61798
rect 34142 61752 34199 61798
rect 34245 61752 34302 61798
rect 34348 61752 34405 61798
rect 34451 61752 34508 61798
rect 34554 61752 34612 61798
rect 34658 61752 34671 61798
rect 33671 61723 34671 61752
rect 37896 61885 38556 61914
rect 37896 61839 37909 61885
rect 37955 61839 38026 61885
rect 38072 61839 38143 61885
rect 38189 61839 38261 61885
rect 38307 61839 38379 61885
rect 38425 61839 38497 61885
rect 38543 61839 38556 61885
rect 37896 61810 38556 61839
rect 43695 61997 43739 62043
rect 43785 61997 43906 62043
rect 43952 61997 44071 62043
rect 44117 61997 44236 62043
rect 44282 61997 44325 62043
rect 43695 61947 44325 61997
rect 50454 62057 51454 62103
rect 39598 61885 39730 61914
rect 39598 61839 39641 61885
rect 39687 61839 39730 61885
rect 39598 61826 39730 61839
rect 50454 62011 50516 62057
rect 50562 62011 50703 62057
rect 50749 62011 50890 62057
rect 50936 62011 51076 62057
rect 51122 62011 51263 62057
rect 51309 62011 51454 62057
rect 50454 61979 51454 62011
rect 43695 61723 44325 61827
rect 33671 61574 34671 61603
rect 37896 61661 38556 61690
rect 37896 61615 37909 61661
rect 37955 61615 38026 61661
rect 38072 61615 38143 61661
rect 38189 61615 38261 61661
rect 38307 61615 38379 61661
rect 38425 61615 38497 61661
rect 38543 61615 38556 61661
rect 37896 61602 38556 61615
rect 50454 61798 51454 61859
rect 50454 61752 50467 61798
rect 50513 61752 50571 61798
rect 50617 61752 50674 61798
rect 50720 61752 50777 61798
rect 50823 61752 50880 61798
rect 50926 61752 50983 61798
rect 51029 61752 51086 61798
rect 51132 61752 51189 61798
rect 51235 61752 51292 61798
rect 51338 61752 51395 61798
rect 51441 61752 51454 61798
rect 50454 61723 51454 61752
rect 33671 61528 33684 61574
rect 33730 61528 33787 61574
rect 33833 61528 33890 61574
rect 33936 61528 33993 61574
rect 34039 61528 34096 61574
rect 34142 61528 34199 61574
rect 34245 61528 34302 61574
rect 34348 61528 34405 61574
rect 34451 61528 34508 61574
rect 34554 61528 34612 61574
rect 34658 61528 34671 61574
rect 33671 61499 34671 61528
rect 39727 61574 40167 61587
rect 39727 61528 39740 61574
rect 39786 61528 39862 61574
rect 39908 61528 39985 61574
rect 40031 61528 40108 61574
rect 40154 61528 40167 61574
rect 39727 61499 40167 61528
rect 43695 61510 44325 61603
rect 50454 61574 51454 61603
rect 33671 61350 34671 61379
rect 33671 61304 33684 61350
rect 33730 61304 33787 61350
rect 33833 61304 33890 61350
rect 33936 61304 33993 61350
rect 34039 61304 34096 61350
rect 34142 61304 34199 61350
rect 34245 61304 34302 61350
rect 34348 61304 34405 61350
rect 34451 61304 34508 61350
rect 34554 61304 34612 61350
rect 34658 61304 34671 61350
rect 33671 61275 34671 61304
rect 39727 61350 40167 61379
rect 39727 61304 39740 61350
rect 39786 61304 39862 61350
rect 39908 61304 39985 61350
rect 40031 61304 40108 61350
rect 40154 61304 40167 61350
rect 39727 61275 40167 61304
rect 43695 61350 44325 61390
rect 50454 61528 50467 61574
rect 50513 61528 50571 61574
rect 50617 61528 50674 61574
rect 50720 61528 50777 61574
rect 50823 61528 50880 61574
rect 50926 61528 50983 61574
rect 51029 61528 51086 61574
rect 51132 61528 51189 61574
rect 51235 61528 51292 61574
rect 51338 61528 51395 61574
rect 51441 61528 51454 61574
rect 50454 61499 51454 61528
rect 43695 61304 43739 61350
rect 43785 61304 43906 61350
rect 43952 61304 44071 61350
rect 44117 61304 44236 61350
rect 44282 61304 44325 61350
rect 43695 61264 44325 61304
rect 33671 61126 34671 61155
rect 33671 61080 33684 61126
rect 33730 61080 33787 61126
rect 33833 61080 33890 61126
rect 33936 61080 33993 61126
rect 34039 61080 34096 61126
rect 34142 61080 34199 61126
rect 34245 61080 34302 61126
rect 34348 61080 34405 61126
rect 34451 61080 34508 61126
rect 34554 61080 34612 61126
rect 34658 61080 34671 61126
rect 33671 61051 34671 61080
rect 39727 61126 40167 61155
rect 39727 61080 39740 61126
rect 39786 61080 39862 61126
rect 39908 61080 39985 61126
rect 40031 61080 40108 61126
rect 40154 61080 40167 61126
rect 39727 61067 40167 61080
rect 50454 61350 51454 61379
rect 50454 61304 50467 61350
rect 50513 61304 50571 61350
rect 50617 61304 50674 61350
rect 50720 61304 50777 61350
rect 50823 61304 50880 61350
rect 50926 61304 50983 61350
rect 51029 61304 51086 61350
rect 51132 61304 51189 61350
rect 51235 61304 51292 61350
rect 51338 61304 51395 61350
rect 51441 61304 51454 61350
rect 50454 61275 51454 61304
rect 37896 61039 38556 61052
rect 43695 61051 44325 61144
rect 50454 61126 51454 61155
rect 50454 61080 50467 61126
rect 50513 61080 50571 61126
rect 50617 61080 50674 61126
rect 50720 61080 50777 61126
rect 50823 61080 50880 61126
rect 50926 61080 50983 61126
rect 51029 61080 51086 61126
rect 51132 61080 51189 61126
rect 51235 61080 51292 61126
rect 51338 61080 51395 61126
rect 51441 61080 51454 61126
rect 37896 60993 37909 61039
rect 37955 60993 38026 61039
rect 38072 60993 38143 61039
rect 38189 60993 38261 61039
rect 38307 60993 38379 61039
rect 38425 60993 38497 61039
rect 38543 60993 38556 61039
rect 37896 60964 38556 60993
rect 33671 60902 34671 60931
rect 33671 60856 33684 60902
rect 33730 60856 33787 60902
rect 33833 60856 33890 60902
rect 33936 60856 33993 60902
rect 34039 60856 34096 60902
rect 34142 60856 34199 60902
rect 34245 60856 34302 60902
rect 34348 60856 34405 60902
rect 34451 60856 34508 60902
rect 34554 60856 34612 60902
rect 34658 60856 34671 60902
rect 33671 60795 34671 60856
rect 33671 60643 34671 60675
rect 33671 60597 33816 60643
rect 33862 60597 34002 60643
rect 34048 60597 34189 60643
rect 34235 60597 34376 60643
rect 34422 60597 34562 60643
rect 34608 60597 34671 60643
rect 50454 61051 51454 61080
rect 37896 60815 38556 60844
rect 37896 60769 37909 60815
rect 37955 60769 38026 60815
rect 38072 60769 38143 60815
rect 38189 60769 38261 60815
rect 38307 60769 38379 60815
rect 38425 60769 38497 60815
rect 38543 60769 38556 60815
rect 37896 60740 38556 60769
rect 39598 60815 39730 60828
rect 43695 60827 44325 60931
rect 39598 60769 39641 60815
rect 39687 60769 39730 60815
rect 39598 60740 39730 60769
rect 50454 60902 51454 60931
rect 50454 60856 50467 60902
rect 50513 60856 50571 60902
rect 50617 60856 50674 60902
rect 50720 60856 50777 60902
rect 50823 60856 50880 60902
rect 50926 60856 50983 60902
rect 51029 60856 51086 60902
rect 51132 60856 51189 60902
rect 51235 60856 51292 60902
rect 51338 60856 51395 60902
rect 51441 60856 51454 60902
rect 50454 60795 51454 60856
rect 43695 60657 44325 60707
rect 33671 60551 34671 60597
rect 37896 60591 38556 60620
rect 37896 60545 37909 60591
rect 37955 60545 38026 60591
rect 38072 60545 38143 60591
rect 38189 60545 38261 60591
rect 38307 60545 38379 60591
rect 38425 60545 38497 60591
rect 38543 60545 38556 60591
rect 37896 60532 38556 60545
rect 39598 60591 39730 60620
rect 39598 60545 39641 60591
rect 39687 60545 39730 60591
rect 43695 60611 43739 60657
rect 43785 60611 43906 60657
rect 43952 60611 44071 60657
rect 44117 60611 44236 60657
rect 44282 60611 44325 60657
rect 50454 60643 51454 60675
rect 43695 60564 44325 60611
rect 39598 60532 39730 60545
rect 50454 60597 50516 60643
rect 50562 60597 50703 60643
rect 50749 60597 50890 60643
rect 50936 60597 51076 60643
rect 51122 60597 51263 60643
rect 51309 60597 51454 60643
rect 50454 60551 51454 60597
rect 33671 60257 34671 60303
rect 33671 60211 33816 60257
rect 33862 60211 34002 60257
rect 34048 60211 34189 60257
rect 34235 60211 34376 60257
rect 34422 60211 34562 60257
rect 34608 60211 34671 60257
rect 37896 60309 38556 60322
rect 37896 60263 37909 60309
rect 37955 60263 38026 60309
rect 38072 60263 38143 60309
rect 38189 60263 38261 60309
rect 38307 60263 38379 60309
rect 38425 60263 38497 60309
rect 38543 60263 38556 60309
rect 37896 60234 38556 60263
rect 39598 60309 39730 60322
rect 39598 60263 39641 60309
rect 39687 60263 39730 60309
rect 39598 60234 39730 60263
rect 43695 60243 44325 60290
rect 33671 60179 34671 60211
rect 33671 59998 34671 60059
rect 33671 59952 33684 59998
rect 33730 59952 33787 59998
rect 33833 59952 33890 59998
rect 33936 59952 33993 59998
rect 34039 59952 34096 59998
rect 34142 59952 34199 59998
rect 34245 59952 34302 59998
rect 34348 59952 34405 59998
rect 34451 59952 34508 59998
rect 34554 59952 34612 59998
rect 34658 59952 34671 59998
rect 33671 59923 34671 59952
rect 37896 60085 38556 60114
rect 37896 60039 37909 60085
rect 37955 60039 38026 60085
rect 38072 60039 38143 60085
rect 38189 60039 38261 60085
rect 38307 60039 38379 60085
rect 38425 60039 38497 60085
rect 38543 60039 38556 60085
rect 37896 60010 38556 60039
rect 43695 60197 43739 60243
rect 43785 60197 43906 60243
rect 43952 60197 44071 60243
rect 44117 60197 44236 60243
rect 44282 60197 44325 60243
rect 43695 60147 44325 60197
rect 50454 60257 51454 60303
rect 39598 60085 39730 60114
rect 39598 60039 39641 60085
rect 39687 60039 39730 60085
rect 39598 60026 39730 60039
rect 50454 60211 50516 60257
rect 50562 60211 50703 60257
rect 50749 60211 50890 60257
rect 50936 60211 51076 60257
rect 51122 60211 51263 60257
rect 51309 60211 51454 60257
rect 50454 60179 51454 60211
rect 43695 59923 44325 60027
rect 33671 59774 34671 59803
rect 37896 59861 38556 59890
rect 37896 59815 37909 59861
rect 37955 59815 38026 59861
rect 38072 59815 38143 59861
rect 38189 59815 38261 59861
rect 38307 59815 38379 59861
rect 38425 59815 38497 59861
rect 38543 59815 38556 59861
rect 37896 59802 38556 59815
rect 50454 59998 51454 60059
rect 50454 59952 50467 59998
rect 50513 59952 50571 59998
rect 50617 59952 50674 59998
rect 50720 59952 50777 59998
rect 50823 59952 50880 59998
rect 50926 59952 50983 59998
rect 51029 59952 51086 59998
rect 51132 59952 51189 59998
rect 51235 59952 51292 59998
rect 51338 59952 51395 59998
rect 51441 59952 51454 59998
rect 50454 59923 51454 59952
rect 33671 59728 33684 59774
rect 33730 59728 33787 59774
rect 33833 59728 33890 59774
rect 33936 59728 33993 59774
rect 34039 59728 34096 59774
rect 34142 59728 34199 59774
rect 34245 59728 34302 59774
rect 34348 59728 34405 59774
rect 34451 59728 34508 59774
rect 34554 59728 34612 59774
rect 34658 59728 34671 59774
rect 33671 59699 34671 59728
rect 39727 59774 40167 59787
rect 39727 59728 39740 59774
rect 39786 59728 39862 59774
rect 39908 59728 39985 59774
rect 40031 59728 40108 59774
rect 40154 59728 40167 59774
rect 39727 59699 40167 59728
rect 43695 59710 44325 59803
rect 50454 59774 51454 59803
rect 33671 59550 34671 59579
rect 33671 59504 33684 59550
rect 33730 59504 33787 59550
rect 33833 59504 33890 59550
rect 33936 59504 33993 59550
rect 34039 59504 34096 59550
rect 34142 59504 34199 59550
rect 34245 59504 34302 59550
rect 34348 59504 34405 59550
rect 34451 59504 34508 59550
rect 34554 59504 34612 59550
rect 34658 59504 34671 59550
rect 33671 59475 34671 59504
rect 39727 59550 40167 59579
rect 39727 59504 39740 59550
rect 39786 59504 39862 59550
rect 39908 59504 39985 59550
rect 40031 59504 40108 59550
rect 40154 59504 40167 59550
rect 39727 59475 40167 59504
rect 43695 59550 44325 59590
rect 50454 59728 50467 59774
rect 50513 59728 50571 59774
rect 50617 59728 50674 59774
rect 50720 59728 50777 59774
rect 50823 59728 50880 59774
rect 50926 59728 50983 59774
rect 51029 59728 51086 59774
rect 51132 59728 51189 59774
rect 51235 59728 51292 59774
rect 51338 59728 51395 59774
rect 51441 59728 51454 59774
rect 50454 59699 51454 59728
rect 43695 59504 43739 59550
rect 43785 59504 43906 59550
rect 43952 59504 44071 59550
rect 44117 59504 44236 59550
rect 44282 59504 44325 59550
rect 43695 59464 44325 59504
rect 33671 59326 34671 59355
rect 33671 59280 33684 59326
rect 33730 59280 33787 59326
rect 33833 59280 33890 59326
rect 33936 59280 33993 59326
rect 34039 59280 34096 59326
rect 34142 59280 34199 59326
rect 34245 59280 34302 59326
rect 34348 59280 34405 59326
rect 34451 59280 34508 59326
rect 34554 59280 34612 59326
rect 34658 59280 34671 59326
rect 33671 59251 34671 59280
rect 39727 59326 40167 59355
rect 39727 59280 39740 59326
rect 39786 59280 39862 59326
rect 39908 59280 39985 59326
rect 40031 59280 40108 59326
rect 40154 59280 40167 59326
rect 39727 59267 40167 59280
rect 50454 59550 51454 59579
rect 50454 59504 50467 59550
rect 50513 59504 50571 59550
rect 50617 59504 50674 59550
rect 50720 59504 50777 59550
rect 50823 59504 50880 59550
rect 50926 59504 50983 59550
rect 51029 59504 51086 59550
rect 51132 59504 51189 59550
rect 51235 59504 51292 59550
rect 51338 59504 51395 59550
rect 51441 59504 51454 59550
rect 50454 59475 51454 59504
rect 37896 59239 38556 59252
rect 43695 59251 44325 59344
rect 50454 59326 51454 59355
rect 50454 59280 50467 59326
rect 50513 59280 50571 59326
rect 50617 59280 50674 59326
rect 50720 59280 50777 59326
rect 50823 59280 50880 59326
rect 50926 59280 50983 59326
rect 51029 59280 51086 59326
rect 51132 59280 51189 59326
rect 51235 59280 51292 59326
rect 51338 59280 51395 59326
rect 51441 59280 51454 59326
rect 37896 59193 37909 59239
rect 37955 59193 38026 59239
rect 38072 59193 38143 59239
rect 38189 59193 38261 59239
rect 38307 59193 38379 59239
rect 38425 59193 38497 59239
rect 38543 59193 38556 59239
rect 37896 59164 38556 59193
rect 33671 59102 34671 59131
rect 33671 59056 33684 59102
rect 33730 59056 33787 59102
rect 33833 59056 33890 59102
rect 33936 59056 33993 59102
rect 34039 59056 34096 59102
rect 34142 59056 34199 59102
rect 34245 59056 34302 59102
rect 34348 59056 34405 59102
rect 34451 59056 34508 59102
rect 34554 59056 34612 59102
rect 34658 59056 34671 59102
rect 33671 58995 34671 59056
rect 33671 58843 34671 58875
rect 33671 58797 33816 58843
rect 33862 58797 34002 58843
rect 34048 58797 34189 58843
rect 34235 58797 34376 58843
rect 34422 58797 34562 58843
rect 34608 58797 34671 58843
rect 50454 59251 51454 59280
rect 37896 59015 38556 59044
rect 37896 58969 37909 59015
rect 37955 58969 38026 59015
rect 38072 58969 38143 59015
rect 38189 58969 38261 59015
rect 38307 58969 38379 59015
rect 38425 58969 38497 59015
rect 38543 58969 38556 59015
rect 37896 58940 38556 58969
rect 39598 59015 39730 59028
rect 43695 59027 44325 59131
rect 39598 58969 39641 59015
rect 39687 58969 39730 59015
rect 39598 58940 39730 58969
rect 50454 59102 51454 59131
rect 50454 59056 50467 59102
rect 50513 59056 50571 59102
rect 50617 59056 50674 59102
rect 50720 59056 50777 59102
rect 50823 59056 50880 59102
rect 50926 59056 50983 59102
rect 51029 59056 51086 59102
rect 51132 59056 51189 59102
rect 51235 59056 51292 59102
rect 51338 59056 51395 59102
rect 51441 59056 51454 59102
rect 50454 58995 51454 59056
rect 43695 58857 44325 58907
rect 33671 58751 34671 58797
rect 37896 58791 38556 58820
rect 37896 58745 37909 58791
rect 37955 58745 38026 58791
rect 38072 58745 38143 58791
rect 38189 58745 38261 58791
rect 38307 58745 38379 58791
rect 38425 58745 38497 58791
rect 38543 58745 38556 58791
rect 37896 58732 38556 58745
rect 39598 58791 39730 58820
rect 39598 58745 39641 58791
rect 39687 58745 39730 58791
rect 43695 58811 43739 58857
rect 43785 58811 43906 58857
rect 43952 58811 44071 58857
rect 44117 58811 44236 58857
rect 44282 58811 44325 58857
rect 50454 58843 51454 58875
rect 43695 58764 44325 58811
rect 39598 58732 39730 58745
rect 50454 58797 50516 58843
rect 50562 58797 50703 58843
rect 50749 58797 50890 58843
rect 50936 58797 51076 58843
rect 51122 58797 51263 58843
rect 51309 58797 51454 58843
rect 50454 58751 51454 58797
rect 33671 58457 34671 58503
rect 33671 58411 33816 58457
rect 33862 58411 34002 58457
rect 34048 58411 34189 58457
rect 34235 58411 34376 58457
rect 34422 58411 34562 58457
rect 34608 58411 34671 58457
rect 37896 58509 38556 58522
rect 37896 58463 37909 58509
rect 37955 58463 38026 58509
rect 38072 58463 38143 58509
rect 38189 58463 38261 58509
rect 38307 58463 38379 58509
rect 38425 58463 38497 58509
rect 38543 58463 38556 58509
rect 37896 58434 38556 58463
rect 39598 58509 39730 58522
rect 39598 58463 39641 58509
rect 39687 58463 39730 58509
rect 39598 58434 39730 58463
rect 43695 58443 44325 58490
rect 33671 58379 34671 58411
rect 33671 58198 34671 58259
rect 33671 58152 33684 58198
rect 33730 58152 33787 58198
rect 33833 58152 33890 58198
rect 33936 58152 33993 58198
rect 34039 58152 34096 58198
rect 34142 58152 34199 58198
rect 34245 58152 34302 58198
rect 34348 58152 34405 58198
rect 34451 58152 34508 58198
rect 34554 58152 34612 58198
rect 34658 58152 34671 58198
rect 33671 58123 34671 58152
rect 37896 58285 38556 58314
rect 37896 58239 37909 58285
rect 37955 58239 38026 58285
rect 38072 58239 38143 58285
rect 38189 58239 38261 58285
rect 38307 58239 38379 58285
rect 38425 58239 38497 58285
rect 38543 58239 38556 58285
rect 37896 58210 38556 58239
rect 43695 58397 43739 58443
rect 43785 58397 43906 58443
rect 43952 58397 44071 58443
rect 44117 58397 44236 58443
rect 44282 58397 44325 58443
rect 43695 58347 44325 58397
rect 50454 58457 51454 58503
rect 39598 58285 39730 58314
rect 39598 58239 39641 58285
rect 39687 58239 39730 58285
rect 39598 58226 39730 58239
rect 50454 58411 50516 58457
rect 50562 58411 50703 58457
rect 50749 58411 50890 58457
rect 50936 58411 51076 58457
rect 51122 58411 51263 58457
rect 51309 58411 51454 58457
rect 50454 58379 51454 58411
rect 43695 58123 44325 58227
rect 33671 57974 34671 58003
rect 37896 58061 38556 58090
rect 37896 58015 37909 58061
rect 37955 58015 38026 58061
rect 38072 58015 38143 58061
rect 38189 58015 38261 58061
rect 38307 58015 38379 58061
rect 38425 58015 38497 58061
rect 38543 58015 38556 58061
rect 37896 58002 38556 58015
rect 50454 58198 51454 58259
rect 50454 58152 50467 58198
rect 50513 58152 50571 58198
rect 50617 58152 50674 58198
rect 50720 58152 50777 58198
rect 50823 58152 50880 58198
rect 50926 58152 50983 58198
rect 51029 58152 51086 58198
rect 51132 58152 51189 58198
rect 51235 58152 51292 58198
rect 51338 58152 51395 58198
rect 51441 58152 51454 58198
rect 50454 58123 51454 58152
rect 33671 57928 33684 57974
rect 33730 57928 33787 57974
rect 33833 57928 33890 57974
rect 33936 57928 33993 57974
rect 34039 57928 34096 57974
rect 34142 57928 34199 57974
rect 34245 57928 34302 57974
rect 34348 57928 34405 57974
rect 34451 57928 34508 57974
rect 34554 57928 34612 57974
rect 34658 57928 34671 57974
rect 33671 57899 34671 57928
rect 39727 57974 40167 57987
rect 39727 57928 39740 57974
rect 39786 57928 39862 57974
rect 39908 57928 39985 57974
rect 40031 57928 40108 57974
rect 40154 57928 40167 57974
rect 39727 57899 40167 57928
rect 43695 57910 44325 58003
rect 50454 57974 51454 58003
rect 33671 57750 34671 57779
rect 33671 57704 33684 57750
rect 33730 57704 33787 57750
rect 33833 57704 33890 57750
rect 33936 57704 33993 57750
rect 34039 57704 34096 57750
rect 34142 57704 34199 57750
rect 34245 57704 34302 57750
rect 34348 57704 34405 57750
rect 34451 57704 34508 57750
rect 34554 57704 34612 57750
rect 34658 57704 34671 57750
rect 33671 57675 34671 57704
rect 39727 57750 40167 57779
rect 39727 57704 39740 57750
rect 39786 57704 39862 57750
rect 39908 57704 39985 57750
rect 40031 57704 40108 57750
rect 40154 57704 40167 57750
rect 39727 57675 40167 57704
rect 43695 57750 44325 57790
rect 50454 57928 50467 57974
rect 50513 57928 50571 57974
rect 50617 57928 50674 57974
rect 50720 57928 50777 57974
rect 50823 57928 50880 57974
rect 50926 57928 50983 57974
rect 51029 57928 51086 57974
rect 51132 57928 51189 57974
rect 51235 57928 51292 57974
rect 51338 57928 51395 57974
rect 51441 57928 51454 57974
rect 50454 57899 51454 57928
rect 43695 57704 43739 57750
rect 43785 57704 43906 57750
rect 43952 57704 44071 57750
rect 44117 57704 44236 57750
rect 44282 57704 44325 57750
rect 43695 57664 44325 57704
rect 33671 57526 34671 57555
rect 33671 57480 33684 57526
rect 33730 57480 33787 57526
rect 33833 57480 33890 57526
rect 33936 57480 33993 57526
rect 34039 57480 34096 57526
rect 34142 57480 34199 57526
rect 34245 57480 34302 57526
rect 34348 57480 34405 57526
rect 34451 57480 34508 57526
rect 34554 57480 34612 57526
rect 34658 57480 34671 57526
rect 33671 57451 34671 57480
rect 39727 57526 40167 57555
rect 39727 57480 39740 57526
rect 39786 57480 39862 57526
rect 39908 57480 39985 57526
rect 40031 57480 40108 57526
rect 40154 57480 40167 57526
rect 39727 57467 40167 57480
rect 50454 57750 51454 57779
rect 50454 57704 50467 57750
rect 50513 57704 50571 57750
rect 50617 57704 50674 57750
rect 50720 57704 50777 57750
rect 50823 57704 50880 57750
rect 50926 57704 50983 57750
rect 51029 57704 51086 57750
rect 51132 57704 51189 57750
rect 51235 57704 51292 57750
rect 51338 57704 51395 57750
rect 51441 57704 51454 57750
rect 50454 57675 51454 57704
rect 37896 57439 38556 57452
rect 43695 57451 44325 57544
rect 50454 57526 51454 57555
rect 50454 57480 50467 57526
rect 50513 57480 50571 57526
rect 50617 57480 50674 57526
rect 50720 57480 50777 57526
rect 50823 57480 50880 57526
rect 50926 57480 50983 57526
rect 51029 57480 51086 57526
rect 51132 57480 51189 57526
rect 51235 57480 51292 57526
rect 51338 57480 51395 57526
rect 51441 57480 51454 57526
rect 37896 57393 37909 57439
rect 37955 57393 38026 57439
rect 38072 57393 38143 57439
rect 38189 57393 38261 57439
rect 38307 57393 38379 57439
rect 38425 57393 38497 57439
rect 38543 57393 38556 57439
rect 37896 57364 38556 57393
rect 33671 57302 34671 57331
rect 33671 57256 33684 57302
rect 33730 57256 33787 57302
rect 33833 57256 33890 57302
rect 33936 57256 33993 57302
rect 34039 57256 34096 57302
rect 34142 57256 34199 57302
rect 34245 57256 34302 57302
rect 34348 57256 34405 57302
rect 34451 57256 34508 57302
rect 34554 57256 34612 57302
rect 34658 57256 34671 57302
rect 33671 57195 34671 57256
rect 33671 57043 34671 57075
rect 33671 56997 33816 57043
rect 33862 56997 34002 57043
rect 34048 56997 34189 57043
rect 34235 56997 34376 57043
rect 34422 56997 34562 57043
rect 34608 56997 34671 57043
rect 50454 57451 51454 57480
rect 37896 57215 38556 57244
rect 37896 57169 37909 57215
rect 37955 57169 38026 57215
rect 38072 57169 38143 57215
rect 38189 57169 38261 57215
rect 38307 57169 38379 57215
rect 38425 57169 38497 57215
rect 38543 57169 38556 57215
rect 37896 57140 38556 57169
rect 39598 57215 39730 57228
rect 43695 57227 44325 57331
rect 39598 57169 39641 57215
rect 39687 57169 39730 57215
rect 39598 57140 39730 57169
rect 50454 57302 51454 57331
rect 50454 57256 50467 57302
rect 50513 57256 50571 57302
rect 50617 57256 50674 57302
rect 50720 57256 50777 57302
rect 50823 57256 50880 57302
rect 50926 57256 50983 57302
rect 51029 57256 51086 57302
rect 51132 57256 51189 57302
rect 51235 57256 51292 57302
rect 51338 57256 51395 57302
rect 51441 57256 51454 57302
rect 50454 57195 51454 57256
rect 43695 57057 44325 57107
rect 33671 56951 34671 56997
rect 37896 56991 38556 57020
rect 37896 56945 37909 56991
rect 37955 56945 38026 56991
rect 38072 56945 38143 56991
rect 38189 56945 38261 56991
rect 38307 56945 38379 56991
rect 38425 56945 38497 56991
rect 38543 56945 38556 56991
rect 37896 56932 38556 56945
rect 39598 56991 39730 57020
rect 39598 56945 39641 56991
rect 39687 56945 39730 56991
rect 43695 57011 43739 57057
rect 43785 57011 43906 57057
rect 43952 57011 44071 57057
rect 44117 57011 44236 57057
rect 44282 57011 44325 57057
rect 50454 57043 51454 57075
rect 43695 56964 44325 57011
rect 39598 56932 39730 56945
rect 50454 56997 50516 57043
rect 50562 56997 50703 57043
rect 50749 56997 50890 57043
rect 50936 56997 51076 57043
rect 51122 56997 51263 57043
rect 51309 56997 51454 57043
rect 50454 56951 51454 56997
rect 33671 56657 34671 56703
rect 33671 56611 33816 56657
rect 33862 56611 34002 56657
rect 34048 56611 34189 56657
rect 34235 56611 34376 56657
rect 34422 56611 34562 56657
rect 34608 56611 34671 56657
rect 37896 56709 38556 56722
rect 37896 56663 37909 56709
rect 37955 56663 38026 56709
rect 38072 56663 38143 56709
rect 38189 56663 38261 56709
rect 38307 56663 38379 56709
rect 38425 56663 38497 56709
rect 38543 56663 38556 56709
rect 37896 56634 38556 56663
rect 39598 56709 39730 56722
rect 39598 56663 39641 56709
rect 39687 56663 39730 56709
rect 39598 56634 39730 56663
rect 43695 56643 44325 56690
rect 33671 56579 34671 56611
rect 33671 56398 34671 56459
rect 33671 56352 33684 56398
rect 33730 56352 33787 56398
rect 33833 56352 33890 56398
rect 33936 56352 33993 56398
rect 34039 56352 34096 56398
rect 34142 56352 34199 56398
rect 34245 56352 34302 56398
rect 34348 56352 34405 56398
rect 34451 56352 34508 56398
rect 34554 56352 34612 56398
rect 34658 56352 34671 56398
rect 33671 56323 34671 56352
rect 37896 56485 38556 56514
rect 37896 56439 37909 56485
rect 37955 56439 38026 56485
rect 38072 56439 38143 56485
rect 38189 56439 38261 56485
rect 38307 56439 38379 56485
rect 38425 56439 38497 56485
rect 38543 56439 38556 56485
rect 37896 56410 38556 56439
rect 43695 56597 43739 56643
rect 43785 56597 43906 56643
rect 43952 56597 44071 56643
rect 44117 56597 44236 56643
rect 44282 56597 44325 56643
rect 43695 56547 44325 56597
rect 50454 56657 51454 56703
rect 39598 56485 39730 56514
rect 39598 56439 39641 56485
rect 39687 56439 39730 56485
rect 39598 56426 39730 56439
rect 50454 56611 50516 56657
rect 50562 56611 50703 56657
rect 50749 56611 50890 56657
rect 50936 56611 51076 56657
rect 51122 56611 51263 56657
rect 51309 56611 51454 56657
rect 50454 56579 51454 56611
rect 43695 56323 44325 56427
rect 33671 56174 34671 56203
rect 37896 56261 38556 56290
rect 37896 56215 37909 56261
rect 37955 56215 38026 56261
rect 38072 56215 38143 56261
rect 38189 56215 38261 56261
rect 38307 56215 38379 56261
rect 38425 56215 38497 56261
rect 38543 56215 38556 56261
rect 37896 56202 38556 56215
rect 50454 56398 51454 56459
rect 50454 56352 50467 56398
rect 50513 56352 50571 56398
rect 50617 56352 50674 56398
rect 50720 56352 50777 56398
rect 50823 56352 50880 56398
rect 50926 56352 50983 56398
rect 51029 56352 51086 56398
rect 51132 56352 51189 56398
rect 51235 56352 51292 56398
rect 51338 56352 51395 56398
rect 51441 56352 51454 56398
rect 50454 56323 51454 56352
rect 33671 56128 33684 56174
rect 33730 56128 33787 56174
rect 33833 56128 33890 56174
rect 33936 56128 33993 56174
rect 34039 56128 34096 56174
rect 34142 56128 34199 56174
rect 34245 56128 34302 56174
rect 34348 56128 34405 56174
rect 34451 56128 34508 56174
rect 34554 56128 34612 56174
rect 34658 56128 34671 56174
rect 33671 56099 34671 56128
rect 39727 56174 40167 56187
rect 39727 56128 39740 56174
rect 39786 56128 39862 56174
rect 39908 56128 39985 56174
rect 40031 56128 40108 56174
rect 40154 56128 40167 56174
rect 39727 56099 40167 56128
rect 43695 56110 44325 56203
rect 50454 56174 51454 56203
rect 33671 55950 34671 55979
rect 33671 55904 33684 55950
rect 33730 55904 33787 55950
rect 33833 55904 33890 55950
rect 33936 55904 33993 55950
rect 34039 55904 34096 55950
rect 34142 55904 34199 55950
rect 34245 55904 34302 55950
rect 34348 55904 34405 55950
rect 34451 55904 34508 55950
rect 34554 55904 34612 55950
rect 34658 55904 34671 55950
rect 33671 55875 34671 55904
rect 39727 55950 40167 55979
rect 39727 55904 39740 55950
rect 39786 55904 39862 55950
rect 39908 55904 39985 55950
rect 40031 55904 40108 55950
rect 40154 55904 40167 55950
rect 39727 55875 40167 55904
rect 43695 55950 44325 55990
rect 50454 56128 50467 56174
rect 50513 56128 50571 56174
rect 50617 56128 50674 56174
rect 50720 56128 50777 56174
rect 50823 56128 50880 56174
rect 50926 56128 50983 56174
rect 51029 56128 51086 56174
rect 51132 56128 51189 56174
rect 51235 56128 51292 56174
rect 51338 56128 51395 56174
rect 51441 56128 51454 56174
rect 50454 56099 51454 56128
rect 43695 55904 43739 55950
rect 43785 55904 43906 55950
rect 43952 55904 44071 55950
rect 44117 55904 44236 55950
rect 44282 55904 44325 55950
rect 43695 55864 44325 55904
rect 33671 55726 34671 55755
rect 33671 55680 33684 55726
rect 33730 55680 33787 55726
rect 33833 55680 33890 55726
rect 33936 55680 33993 55726
rect 34039 55680 34096 55726
rect 34142 55680 34199 55726
rect 34245 55680 34302 55726
rect 34348 55680 34405 55726
rect 34451 55680 34508 55726
rect 34554 55680 34612 55726
rect 34658 55680 34671 55726
rect 33671 55651 34671 55680
rect 39727 55726 40167 55755
rect 39727 55680 39740 55726
rect 39786 55680 39862 55726
rect 39908 55680 39985 55726
rect 40031 55680 40108 55726
rect 40154 55680 40167 55726
rect 39727 55667 40167 55680
rect 50454 55950 51454 55979
rect 50454 55904 50467 55950
rect 50513 55904 50571 55950
rect 50617 55904 50674 55950
rect 50720 55904 50777 55950
rect 50823 55904 50880 55950
rect 50926 55904 50983 55950
rect 51029 55904 51086 55950
rect 51132 55904 51189 55950
rect 51235 55904 51292 55950
rect 51338 55904 51395 55950
rect 51441 55904 51454 55950
rect 50454 55875 51454 55904
rect 37896 55639 38556 55652
rect 43695 55651 44325 55744
rect 50454 55726 51454 55755
rect 50454 55680 50467 55726
rect 50513 55680 50571 55726
rect 50617 55680 50674 55726
rect 50720 55680 50777 55726
rect 50823 55680 50880 55726
rect 50926 55680 50983 55726
rect 51029 55680 51086 55726
rect 51132 55680 51189 55726
rect 51235 55680 51292 55726
rect 51338 55680 51395 55726
rect 51441 55680 51454 55726
rect 37896 55593 37909 55639
rect 37955 55593 38026 55639
rect 38072 55593 38143 55639
rect 38189 55593 38261 55639
rect 38307 55593 38379 55639
rect 38425 55593 38497 55639
rect 38543 55593 38556 55639
rect 37896 55564 38556 55593
rect 33671 55502 34671 55531
rect 33671 55456 33684 55502
rect 33730 55456 33787 55502
rect 33833 55456 33890 55502
rect 33936 55456 33993 55502
rect 34039 55456 34096 55502
rect 34142 55456 34199 55502
rect 34245 55456 34302 55502
rect 34348 55456 34405 55502
rect 34451 55456 34508 55502
rect 34554 55456 34612 55502
rect 34658 55456 34671 55502
rect 33671 55395 34671 55456
rect 33671 55243 34671 55275
rect 33671 55197 33816 55243
rect 33862 55197 34002 55243
rect 34048 55197 34189 55243
rect 34235 55197 34376 55243
rect 34422 55197 34562 55243
rect 34608 55197 34671 55243
rect 50454 55651 51454 55680
rect 37896 55415 38556 55444
rect 37896 55369 37909 55415
rect 37955 55369 38026 55415
rect 38072 55369 38143 55415
rect 38189 55369 38261 55415
rect 38307 55369 38379 55415
rect 38425 55369 38497 55415
rect 38543 55369 38556 55415
rect 37896 55340 38556 55369
rect 39598 55415 39730 55428
rect 43695 55427 44325 55531
rect 39598 55369 39641 55415
rect 39687 55369 39730 55415
rect 39598 55340 39730 55369
rect 50454 55502 51454 55531
rect 50454 55456 50467 55502
rect 50513 55456 50571 55502
rect 50617 55456 50674 55502
rect 50720 55456 50777 55502
rect 50823 55456 50880 55502
rect 50926 55456 50983 55502
rect 51029 55456 51086 55502
rect 51132 55456 51189 55502
rect 51235 55456 51292 55502
rect 51338 55456 51395 55502
rect 51441 55456 51454 55502
rect 50454 55395 51454 55456
rect 43695 55257 44325 55307
rect 33671 55151 34671 55197
rect 37896 55191 38556 55220
rect 37896 55145 37909 55191
rect 37955 55145 38026 55191
rect 38072 55145 38143 55191
rect 38189 55145 38261 55191
rect 38307 55145 38379 55191
rect 38425 55145 38497 55191
rect 38543 55145 38556 55191
rect 37896 55132 38556 55145
rect 39598 55191 39730 55220
rect 39598 55145 39641 55191
rect 39687 55145 39730 55191
rect 43695 55211 43739 55257
rect 43785 55211 43906 55257
rect 43952 55211 44071 55257
rect 44117 55211 44236 55257
rect 44282 55211 44325 55257
rect 50454 55243 51454 55275
rect 43695 55164 44325 55211
rect 39598 55132 39730 55145
rect 50454 55197 50516 55243
rect 50562 55197 50703 55243
rect 50749 55197 50890 55243
rect 50936 55197 51076 55243
rect 51122 55197 51263 55243
rect 51309 55197 51454 55243
rect 50454 55151 51454 55197
rect 33671 54857 34671 54903
rect 33671 54811 33816 54857
rect 33862 54811 34002 54857
rect 34048 54811 34189 54857
rect 34235 54811 34376 54857
rect 34422 54811 34562 54857
rect 34608 54811 34671 54857
rect 37896 54909 38556 54922
rect 37896 54863 37909 54909
rect 37955 54863 38026 54909
rect 38072 54863 38143 54909
rect 38189 54863 38261 54909
rect 38307 54863 38379 54909
rect 38425 54863 38497 54909
rect 38543 54863 38556 54909
rect 37896 54834 38556 54863
rect 39598 54909 39730 54922
rect 39598 54863 39641 54909
rect 39687 54863 39730 54909
rect 39598 54834 39730 54863
rect 43695 54843 44325 54890
rect 33671 54779 34671 54811
rect 33671 54598 34671 54659
rect 33671 54552 33684 54598
rect 33730 54552 33787 54598
rect 33833 54552 33890 54598
rect 33936 54552 33993 54598
rect 34039 54552 34096 54598
rect 34142 54552 34199 54598
rect 34245 54552 34302 54598
rect 34348 54552 34405 54598
rect 34451 54552 34508 54598
rect 34554 54552 34612 54598
rect 34658 54552 34671 54598
rect 33671 54523 34671 54552
rect 37896 54685 38556 54714
rect 37896 54639 37909 54685
rect 37955 54639 38026 54685
rect 38072 54639 38143 54685
rect 38189 54639 38261 54685
rect 38307 54639 38379 54685
rect 38425 54639 38497 54685
rect 38543 54639 38556 54685
rect 37896 54610 38556 54639
rect 43695 54797 43739 54843
rect 43785 54797 43906 54843
rect 43952 54797 44071 54843
rect 44117 54797 44236 54843
rect 44282 54797 44325 54843
rect 43695 54747 44325 54797
rect 50454 54857 51454 54903
rect 39598 54685 39730 54714
rect 39598 54639 39641 54685
rect 39687 54639 39730 54685
rect 39598 54626 39730 54639
rect 50454 54811 50516 54857
rect 50562 54811 50703 54857
rect 50749 54811 50890 54857
rect 50936 54811 51076 54857
rect 51122 54811 51263 54857
rect 51309 54811 51454 54857
rect 50454 54779 51454 54811
rect 43695 54523 44325 54627
rect 33671 54374 34671 54403
rect 37896 54461 38556 54490
rect 37896 54415 37909 54461
rect 37955 54415 38026 54461
rect 38072 54415 38143 54461
rect 38189 54415 38261 54461
rect 38307 54415 38379 54461
rect 38425 54415 38497 54461
rect 38543 54415 38556 54461
rect 37896 54402 38556 54415
rect 50454 54598 51454 54659
rect 50454 54552 50467 54598
rect 50513 54552 50571 54598
rect 50617 54552 50674 54598
rect 50720 54552 50777 54598
rect 50823 54552 50880 54598
rect 50926 54552 50983 54598
rect 51029 54552 51086 54598
rect 51132 54552 51189 54598
rect 51235 54552 51292 54598
rect 51338 54552 51395 54598
rect 51441 54552 51454 54598
rect 50454 54523 51454 54552
rect 33671 54328 33684 54374
rect 33730 54328 33787 54374
rect 33833 54328 33890 54374
rect 33936 54328 33993 54374
rect 34039 54328 34096 54374
rect 34142 54328 34199 54374
rect 34245 54328 34302 54374
rect 34348 54328 34405 54374
rect 34451 54328 34508 54374
rect 34554 54328 34612 54374
rect 34658 54328 34671 54374
rect 33671 54299 34671 54328
rect 39727 54374 40167 54387
rect 39727 54328 39740 54374
rect 39786 54328 39862 54374
rect 39908 54328 39985 54374
rect 40031 54328 40108 54374
rect 40154 54328 40167 54374
rect 39727 54299 40167 54328
rect 43695 54310 44325 54403
rect 50454 54374 51454 54403
rect 33671 54150 34671 54179
rect 33671 54104 33684 54150
rect 33730 54104 33787 54150
rect 33833 54104 33890 54150
rect 33936 54104 33993 54150
rect 34039 54104 34096 54150
rect 34142 54104 34199 54150
rect 34245 54104 34302 54150
rect 34348 54104 34405 54150
rect 34451 54104 34508 54150
rect 34554 54104 34612 54150
rect 34658 54104 34671 54150
rect 33671 54075 34671 54104
rect 39727 54150 40167 54179
rect 39727 54104 39740 54150
rect 39786 54104 39862 54150
rect 39908 54104 39985 54150
rect 40031 54104 40108 54150
rect 40154 54104 40167 54150
rect 39727 54075 40167 54104
rect 43695 54150 44325 54190
rect 50454 54328 50467 54374
rect 50513 54328 50571 54374
rect 50617 54328 50674 54374
rect 50720 54328 50777 54374
rect 50823 54328 50880 54374
rect 50926 54328 50983 54374
rect 51029 54328 51086 54374
rect 51132 54328 51189 54374
rect 51235 54328 51292 54374
rect 51338 54328 51395 54374
rect 51441 54328 51454 54374
rect 50454 54299 51454 54328
rect 43695 54104 43739 54150
rect 43785 54104 43906 54150
rect 43952 54104 44071 54150
rect 44117 54104 44236 54150
rect 44282 54104 44325 54150
rect 43695 54064 44325 54104
rect 33671 53926 34671 53955
rect 33671 53880 33684 53926
rect 33730 53880 33787 53926
rect 33833 53880 33890 53926
rect 33936 53880 33993 53926
rect 34039 53880 34096 53926
rect 34142 53880 34199 53926
rect 34245 53880 34302 53926
rect 34348 53880 34405 53926
rect 34451 53880 34508 53926
rect 34554 53880 34612 53926
rect 34658 53880 34671 53926
rect 33671 53851 34671 53880
rect 39727 53926 40167 53955
rect 39727 53880 39740 53926
rect 39786 53880 39862 53926
rect 39908 53880 39985 53926
rect 40031 53880 40108 53926
rect 40154 53880 40167 53926
rect 39727 53867 40167 53880
rect 50454 54150 51454 54179
rect 50454 54104 50467 54150
rect 50513 54104 50571 54150
rect 50617 54104 50674 54150
rect 50720 54104 50777 54150
rect 50823 54104 50880 54150
rect 50926 54104 50983 54150
rect 51029 54104 51086 54150
rect 51132 54104 51189 54150
rect 51235 54104 51292 54150
rect 51338 54104 51395 54150
rect 51441 54104 51454 54150
rect 50454 54075 51454 54104
rect 37896 53839 38556 53852
rect 43695 53851 44325 53944
rect 50454 53926 51454 53955
rect 50454 53880 50467 53926
rect 50513 53880 50571 53926
rect 50617 53880 50674 53926
rect 50720 53880 50777 53926
rect 50823 53880 50880 53926
rect 50926 53880 50983 53926
rect 51029 53880 51086 53926
rect 51132 53880 51189 53926
rect 51235 53880 51292 53926
rect 51338 53880 51395 53926
rect 51441 53880 51454 53926
rect 37896 53793 37909 53839
rect 37955 53793 38026 53839
rect 38072 53793 38143 53839
rect 38189 53793 38261 53839
rect 38307 53793 38379 53839
rect 38425 53793 38497 53839
rect 38543 53793 38556 53839
rect 37896 53764 38556 53793
rect 33671 53702 34671 53731
rect 33671 53656 33684 53702
rect 33730 53656 33787 53702
rect 33833 53656 33890 53702
rect 33936 53656 33993 53702
rect 34039 53656 34096 53702
rect 34142 53656 34199 53702
rect 34245 53656 34302 53702
rect 34348 53656 34405 53702
rect 34451 53656 34508 53702
rect 34554 53656 34612 53702
rect 34658 53656 34671 53702
rect 33671 53595 34671 53656
rect 33671 53443 34671 53475
rect 33671 53397 33816 53443
rect 33862 53397 34002 53443
rect 34048 53397 34189 53443
rect 34235 53397 34376 53443
rect 34422 53397 34562 53443
rect 34608 53397 34671 53443
rect 50454 53851 51454 53880
rect 37896 53615 38556 53644
rect 37896 53569 37909 53615
rect 37955 53569 38026 53615
rect 38072 53569 38143 53615
rect 38189 53569 38261 53615
rect 38307 53569 38379 53615
rect 38425 53569 38497 53615
rect 38543 53569 38556 53615
rect 37896 53540 38556 53569
rect 39598 53615 39730 53628
rect 43695 53627 44325 53731
rect 39598 53569 39641 53615
rect 39687 53569 39730 53615
rect 39598 53540 39730 53569
rect 50454 53702 51454 53731
rect 50454 53656 50467 53702
rect 50513 53656 50571 53702
rect 50617 53656 50674 53702
rect 50720 53656 50777 53702
rect 50823 53656 50880 53702
rect 50926 53656 50983 53702
rect 51029 53656 51086 53702
rect 51132 53656 51189 53702
rect 51235 53656 51292 53702
rect 51338 53656 51395 53702
rect 51441 53656 51454 53702
rect 50454 53595 51454 53656
rect 43695 53457 44325 53507
rect 33671 53351 34671 53397
rect 37896 53391 38556 53420
rect 37896 53345 37909 53391
rect 37955 53345 38026 53391
rect 38072 53345 38143 53391
rect 38189 53345 38261 53391
rect 38307 53345 38379 53391
rect 38425 53345 38497 53391
rect 38543 53345 38556 53391
rect 37896 53332 38556 53345
rect 39598 53391 39730 53420
rect 39598 53345 39641 53391
rect 39687 53345 39730 53391
rect 43695 53411 43739 53457
rect 43785 53411 43906 53457
rect 43952 53411 44071 53457
rect 44117 53411 44236 53457
rect 44282 53411 44325 53457
rect 50454 53443 51454 53475
rect 43695 53364 44325 53411
rect 39598 53332 39730 53345
rect 50454 53397 50516 53443
rect 50562 53397 50703 53443
rect 50749 53397 50890 53443
rect 50936 53397 51076 53443
rect 51122 53397 51263 53443
rect 51309 53397 51454 53443
rect 50454 53351 51454 53397
rect 33671 53057 34671 53103
rect 33671 53011 33816 53057
rect 33862 53011 34002 53057
rect 34048 53011 34189 53057
rect 34235 53011 34376 53057
rect 34422 53011 34562 53057
rect 34608 53011 34671 53057
rect 37896 53109 38556 53122
rect 37896 53063 37909 53109
rect 37955 53063 38026 53109
rect 38072 53063 38143 53109
rect 38189 53063 38261 53109
rect 38307 53063 38379 53109
rect 38425 53063 38497 53109
rect 38543 53063 38556 53109
rect 37896 53034 38556 53063
rect 39598 53109 39730 53122
rect 39598 53063 39641 53109
rect 39687 53063 39730 53109
rect 39598 53034 39730 53063
rect 43695 53043 44325 53090
rect 33671 52979 34671 53011
rect 33671 52798 34671 52859
rect 33671 52752 33684 52798
rect 33730 52752 33787 52798
rect 33833 52752 33890 52798
rect 33936 52752 33993 52798
rect 34039 52752 34096 52798
rect 34142 52752 34199 52798
rect 34245 52752 34302 52798
rect 34348 52752 34405 52798
rect 34451 52752 34508 52798
rect 34554 52752 34612 52798
rect 34658 52752 34671 52798
rect 33671 52723 34671 52752
rect 37896 52885 38556 52914
rect 37896 52839 37909 52885
rect 37955 52839 38026 52885
rect 38072 52839 38143 52885
rect 38189 52839 38261 52885
rect 38307 52839 38379 52885
rect 38425 52839 38497 52885
rect 38543 52839 38556 52885
rect 37896 52810 38556 52839
rect 43695 52997 43739 53043
rect 43785 52997 43906 53043
rect 43952 52997 44071 53043
rect 44117 52997 44236 53043
rect 44282 52997 44325 53043
rect 43695 52947 44325 52997
rect 50454 53057 51454 53103
rect 39598 52885 39730 52914
rect 39598 52839 39641 52885
rect 39687 52839 39730 52885
rect 39598 52826 39730 52839
rect 50454 53011 50516 53057
rect 50562 53011 50703 53057
rect 50749 53011 50890 53057
rect 50936 53011 51076 53057
rect 51122 53011 51263 53057
rect 51309 53011 51454 53057
rect 50454 52979 51454 53011
rect 43695 52723 44325 52827
rect 33671 52574 34671 52603
rect 37896 52661 38556 52690
rect 37896 52615 37909 52661
rect 37955 52615 38026 52661
rect 38072 52615 38143 52661
rect 38189 52615 38261 52661
rect 38307 52615 38379 52661
rect 38425 52615 38497 52661
rect 38543 52615 38556 52661
rect 37896 52602 38556 52615
rect 50454 52798 51454 52859
rect 50454 52752 50467 52798
rect 50513 52752 50571 52798
rect 50617 52752 50674 52798
rect 50720 52752 50777 52798
rect 50823 52752 50880 52798
rect 50926 52752 50983 52798
rect 51029 52752 51086 52798
rect 51132 52752 51189 52798
rect 51235 52752 51292 52798
rect 51338 52752 51395 52798
rect 51441 52752 51454 52798
rect 50454 52723 51454 52752
rect 33671 52528 33684 52574
rect 33730 52528 33787 52574
rect 33833 52528 33890 52574
rect 33936 52528 33993 52574
rect 34039 52528 34096 52574
rect 34142 52528 34199 52574
rect 34245 52528 34302 52574
rect 34348 52528 34405 52574
rect 34451 52528 34508 52574
rect 34554 52528 34612 52574
rect 34658 52528 34671 52574
rect 33671 52499 34671 52528
rect 39727 52574 40167 52587
rect 39727 52528 39740 52574
rect 39786 52528 39862 52574
rect 39908 52528 39985 52574
rect 40031 52528 40108 52574
rect 40154 52528 40167 52574
rect 39727 52499 40167 52528
rect 43695 52510 44325 52603
rect 50454 52574 51454 52603
rect 33671 52350 34671 52379
rect 33671 52304 33684 52350
rect 33730 52304 33787 52350
rect 33833 52304 33890 52350
rect 33936 52304 33993 52350
rect 34039 52304 34096 52350
rect 34142 52304 34199 52350
rect 34245 52304 34302 52350
rect 34348 52304 34405 52350
rect 34451 52304 34508 52350
rect 34554 52304 34612 52350
rect 34658 52304 34671 52350
rect 33671 52275 34671 52304
rect 39727 52350 40167 52379
rect 39727 52304 39740 52350
rect 39786 52304 39862 52350
rect 39908 52304 39985 52350
rect 40031 52304 40108 52350
rect 40154 52304 40167 52350
rect 39727 52275 40167 52304
rect 43695 52350 44325 52390
rect 50454 52528 50467 52574
rect 50513 52528 50571 52574
rect 50617 52528 50674 52574
rect 50720 52528 50777 52574
rect 50823 52528 50880 52574
rect 50926 52528 50983 52574
rect 51029 52528 51086 52574
rect 51132 52528 51189 52574
rect 51235 52528 51292 52574
rect 51338 52528 51395 52574
rect 51441 52528 51454 52574
rect 50454 52499 51454 52528
rect 43695 52304 43739 52350
rect 43785 52304 43906 52350
rect 43952 52304 44071 52350
rect 44117 52304 44236 52350
rect 44282 52304 44325 52350
rect 43695 52264 44325 52304
rect 33671 52126 34671 52155
rect 33671 52080 33684 52126
rect 33730 52080 33787 52126
rect 33833 52080 33890 52126
rect 33936 52080 33993 52126
rect 34039 52080 34096 52126
rect 34142 52080 34199 52126
rect 34245 52080 34302 52126
rect 34348 52080 34405 52126
rect 34451 52080 34508 52126
rect 34554 52080 34612 52126
rect 34658 52080 34671 52126
rect 33671 52051 34671 52080
rect 39727 52126 40167 52155
rect 39727 52080 39740 52126
rect 39786 52080 39862 52126
rect 39908 52080 39985 52126
rect 40031 52080 40108 52126
rect 40154 52080 40167 52126
rect 39727 52067 40167 52080
rect 50454 52350 51454 52379
rect 50454 52304 50467 52350
rect 50513 52304 50571 52350
rect 50617 52304 50674 52350
rect 50720 52304 50777 52350
rect 50823 52304 50880 52350
rect 50926 52304 50983 52350
rect 51029 52304 51086 52350
rect 51132 52304 51189 52350
rect 51235 52304 51292 52350
rect 51338 52304 51395 52350
rect 51441 52304 51454 52350
rect 50454 52275 51454 52304
rect 37896 52039 38556 52052
rect 43695 52051 44325 52144
rect 50454 52126 51454 52155
rect 50454 52080 50467 52126
rect 50513 52080 50571 52126
rect 50617 52080 50674 52126
rect 50720 52080 50777 52126
rect 50823 52080 50880 52126
rect 50926 52080 50983 52126
rect 51029 52080 51086 52126
rect 51132 52080 51189 52126
rect 51235 52080 51292 52126
rect 51338 52080 51395 52126
rect 51441 52080 51454 52126
rect 37896 51993 37909 52039
rect 37955 51993 38026 52039
rect 38072 51993 38143 52039
rect 38189 51993 38261 52039
rect 38307 51993 38379 52039
rect 38425 51993 38497 52039
rect 38543 51993 38556 52039
rect 37896 51964 38556 51993
rect 33671 51902 34671 51931
rect 33671 51856 33684 51902
rect 33730 51856 33787 51902
rect 33833 51856 33890 51902
rect 33936 51856 33993 51902
rect 34039 51856 34096 51902
rect 34142 51856 34199 51902
rect 34245 51856 34302 51902
rect 34348 51856 34405 51902
rect 34451 51856 34508 51902
rect 34554 51856 34612 51902
rect 34658 51856 34671 51902
rect 33671 51795 34671 51856
rect 33671 51643 34671 51675
rect 33671 51597 33816 51643
rect 33862 51597 34002 51643
rect 34048 51597 34189 51643
rect 34235 51597 34376 51643
rect 34422 51597 34562 51643
rect 34608 51597 34671 51643
rect 50454 52051 51454 52080
rect 37896 51815 38556 51844
rect 37896 51769 37909 51815
rect 37955 51769 38026 51815
rect 38072 51769 38143 51815
rect 38189 51769 38261 51815
rect 38307 51769 38379 51815
rect 38425 51769 38497 51815
rect 38543 51769 38556 51815
rect 37896 51740 38556 51769
rect 39598 51815 39730 51828
rect 43695 51827 44325 51931
rect 39598 51769 39641 51815
rect 39687 51769 39730 51815
rect 39598 51740 39730 51769
rect 50454 51902 51454 51931
rect 50454 51856 50467 51902
rect 50513 51856 50571 51902
rect 50617 51856 50674 51902
rect 50720 51856 50777 51902
rect 50823 51856 50880 51902
rect 50926 51856 50983 51902
rect 51029 51856 51086 51902
rect 51132 51856 51189 51902
rect 51235 51856 51292 51902
rect 51338 51856 51395 51902
rect 51441 51856 51454 51902
rect 50454 51795 51454 51856
rect 43695 51657 44325 51707
rect 33671 51551 34671 51597
rect 37896 51591 38556 51620
rect 37896 51545 37909 51591
rect 37955 51545 38026 51591
rect 38072 51545 38143 51591
rect 38189 51545 38261 51591
rect 38307 51545 38379 51591
rect 38425 51545 38497 51591
rect 38543 51545 38556 51591
rect 37896 51532 38556 51545
rect 39598 51591 39730 51620
rect 39598 51545 39641 51591
rect 39687 51545 39730 51591
rect 43695 51611 43739 51657
rect 43785 51611 43906 51657
rect 43952 51611 44071 51657
rect 44117 51611 44236 51657
rect 44282 51611 44325 51657
rect 50454 51643 51454 51675
rect 43695 51564 44325 51611
rect 39598 51532 39730 51545
rect 50454 51597 50516 51643
rect 50562 51597 50703 51643
rect 50749 51597 50890 51643
rect 50936 51597 51076 51643
rect 51122 51597 51263 51643
rect 51309 51597 51454 51643
rect 50454 51551 51454 51597
rect 33671 51257 34671 51303
rect 33671 51211 33816 51257
rect 33862 51211 34002 51257
rect 34048 51211 34189 51257
rect 34235 51211 34376 51257
rect 34422 51211 34562 51257
rect 34608 51211 34671 51257
rect 37896 51309 38556 51322
rect 37896 51263 37909 51309
rect 37955 51263 38026 51309
rect 38072 51263 38143 51309
rect 38189 51263 38261 51309
rect 38307 51263 38379 51309
rect 38425 51263 38497 51309
rect 38543 51263 38556 51309
rect 37896 51234 38556 51263
rect 39598 51309 39730 51322
rect 39598 51263 39641 51309
rect 39687 51263 39730 51309
rect 39598 51234 39730 51263
rect 43695 51243 44325 51290
rect 33671 51179 34671 51211
rect 33671 50998 34671 51059
rect 33671 50952 33684 50998
rect 33730 50952 33787 50998
rect 33833 50952 33890 50998
rect 33936 50952 33993 50998
rect 34039 50952 34096 50998
rect 34142 50952 34199 50998
rect 34245 50952 34302 50998
rect 34348 50952 34405 50998
rect 34451 50952 34508 50998
rect 34554 50952 34612 50998
rect 34658 50952 34671 50998
rect 33671 50923 34671 50952
rect 37896 51085 38556 51114
rect 37896 51039 37909 51085
rect 37955 51039 38026 51085
rect 38072 51039 38143 51085
rect 38189 51039 38261 51085
rect 38307 51039 38379 51085
rect 38425 51039 38497 51085
rect 38543 51039 38556 51085
rect 37896 51010 38556 51039
rect 43695 51197 43739 51243
rect 43785 51197 43906 51243
rect 43952 51197 44071 51243
rect 44117 51197 44236 51243
rect 44282 51197 44325 51243
rect 43695 51147 44325 51197
rect 50454 51257 51454 51303
rect 39598 51085 39730 51114
rect 39598 51039 39641 51085
rect 39687 51039 39730 51085
rect 39598 51026 39730 51039
rect 50454 51211 50516 51257
rect 50562 51211 50703 51257
rect 50749 51211 50890 51257
rect 50936 51211 51076 51257
rect 51122 51211 51263 51257
rect 51309 51211 51454 51257
rect 50454 51179 51454 51211
rect 43695 50923 44325 51027
rect 33671 50774 34671 50803
rect 37896 50861 38556 50890
rect 37896 50815 37909 50861
rect 37955 50815 38026 50861
rect 38072 50815 38143 50861
rect 38189 50815 38261 50861
rect 38307 50815 38379 50861
rect 38425 50815 38497 50861
rect 38543 50815 38556 50861
rect 37896 50802 38556 50815
rect 50454 50998 51454 51059
rect 50454 50952 50467 50998
rect 50513 50952 50571 50998
rect 50617 50952 50674 50998
rect 50720 50952 50777 50998
rect 50823 50952 50880 50998
rect 50926 50952 50983 50998
rect 51029 50952 51086 50998
rect 51132 50952 51189 50998
rect 51235 50952 51292 50998
rect 51338 50952 51395 50998
rect 51441 50952 51454 50998
rect 50454 50923 51454 50952
rect 33671 50728 33684 50774
rect 33730 50728 33787 50774
rect 33833 50728 33890 50774
rect 33936 50728 33993 50774
rect 34039 50728 34096 50774
rect 34142 50728 34199 50774
rect 34245 50728 34302 50774
rect 34348 50728 34405 50774
rect 34451 50728 34508 50774
rect 34554 50728 34612 50774
rect 34658 50728 34671 50774
rect 33671 50699 34671 50728
rect 39727 50774 40167 50787
rect 39727 50728 39740 50774
rect 39786 50728 39862 50774
rect 39908 50728 39985 50774
rect 40031 50728 40108 50774
rect 40154 50728 40167 50774
rect 39727 50699 40167 50728
rect 43695 50710 44325 50803
rect 50454 50774 51454 50803
rect 33671 50550 34671 50579
rect 33671 50504 33684 50550
rect 33730 50504 33787 50550
rect 33833 50504 33890 50550
rect 33936 50504 33993 50550
rect 34039 50504 34096 50550
rect 34142 50504 34199 50550
rect 34245 50504 34302 50550
rect 34348 50504 34405 50550
rect 34451 50504 34508 50550
rect 34554 50504 34612 50550
rect 34658 50504 34671 50550
rect 33671 50475 34671 50504
rect 39727 50550 40167 50579
rect 39727 50504 39740 50550
rect 39786 50504 39862 50550
rect 39908 50504 39985 50550
rect 40031 50504 40108 50550
rect 40154 50504 40167 50550
rect 39727 50475 40167 50504
rect 43695 50550 44325 50590
rect 50454 50728 50467 50774
rect 50513 50728 50571 50774
rect 50617 50728 50674 50774
rect 50720 50728 50777 50774
rect 50823 50728 50880 50774
rect 50926 50728 50983 50774
rect 51029 50728 51086 50774
rect 51132 50728 51189 50774
rect 51235 50728 51292 50774
rect 51338 50728 51395 50774
rect 51441 50728 51454 50774
rect 50454 50699 51454 50728
rect 43695 50504 43739 50550
rect 43785 50504 43906 50550
rect 43952 50504 44071 50550
rect 44117 50504 44236 50550
rect 44282 50504 44325 50550
rect 43695 50464 44325 50504
rect 33671 50326 34671 50355
rect 33671 50280 33684 50326
rect 33730 50280 33787 50326
rect 33833 50280 33890 50326
rect 33936 50280 33993 50326
rect 34039 50280 34096 50326
rect 34142 50280 34199 50326
rect 34245 50280 34302 50326
rect 34348 50280 34405 50326
rect 34451 50280 34508 50326
rect 34554 50280 34612 50326
rect 34658 50280 34671 50326
rect 33671 50251 34671 50280
rect 39727 50326 40167 50355
rect 39727 50280 39740 50326
rect 39786 50280 39862 50326
rect 39908 50280 39985 50326
rect 40031 50280 40108 50326
rect 40154 50280 40167 50326
rect 39727 50267 40167 50280
rect 50454 50550 51454 50579
rect 50454 50504 50467 50550
rect 50513 50504 50571 50550
rect 50617 50504 50674 50550
rect 50720 50504 50777 50550
rect 50823 50504 50880 50550
rect 50926 50504 50983 50550
rect 51029 50504 51086 50550
rect 51132 50504 51189 50550
rect 51235 50504 51292 50550
rect 51338 50504 51395 50550
rect 51441 50504 51454 50550
rect 50454 50475 51454 50504
rect 37896 50239 38556 50252
rect 43695 50251 44325 50344
rect 50454 50326 51454 50355
rect 50454 50280 50467 50326
rect 50513 50280 50571 50326
rect 50617 50280 50674 50326
rect 50720 50280 50777 50326
rect 50823 50280 50880 50326
rect 50926 50280 50983 50326
rect 51029 50280 51086 50326
rect 51132 50280 51189 50326
rect 51235 50280 51292 50326
rect 51338 50280 51395 50326
rect 51441 50280 51454 50326
rect 37896 50193 37909 50239
rect 37955 50193 38026 50239
rect 38072 50193 38143 50239
rect 38189 50193 38261 50239
rect 38307 50193 38379 50239
rect 38425 50193 38497 50239
rect 38543 50193 38556 50239
rect 37896 50164 38556 50193
rect 33671 50102 34671 50131
rect 33671 50056 33684 50102
rect 33730 50056 33787 50102
rect 33833 50056 33890 50102
rect 33936 50056 33993 50102
rect 34039 50056 34096 50102
rect 34142 50056 34199 50102
rect 34245 50056 34302 50102
rect 34348 50056 34405 50102
rect 34451 50056 34508 50102
rect 34554 50056 34612 50102
rect 34658 50056 34671 50102
rect 33671 49995 34671 50056
rect 33671 49843 34671 49875
rect 33671 49797 33816 49843
rect 33862 49797 34002 49843
rect 34048 49797 34189 49843
rect 34235 49797 34376 49843
rect 34422 49797 34562 49843
rect 34608 49797 34671 49843
rect 50454 50251 51454 50280
rect 37896 50015 38556 50044
rect 37896 49969 37909 50015
rect 37955 49969 38026 50015
rect 38072 49969 38143 50015
rect 38189 49969 38261 50015
rect 38307 49969 38379 50015
rect 38425 49969 38497 50015
rect 38543 49969 38556 50015
rect 37896 49940 38556 49969
rect 39598 50015 39730 50028
rect 43695 50027 44325 50131
rect 39598 49969 39641 50015
rect 39687 49969 39730 50015
rect 39598 49940 39730 49969
rect 50454 50102 51454 50131
rect 50454 50056 50467 50102
rect 50513 50056 50571 50102
rect 50617 50056 50674 50102
rect 50720 50056 50777 50102
rect 50823 50056 50880 50102
rect 50926 50056 50983 50102
rect 51029 50056 51086 50102
rect 51132 50056 51189 50102
rect 51235 50056 51292 50102
rect 51338 50056 51395 50102
rect 51441 50056 51454 50102
rect 50454 49995 51454 50056
rect 43695 49857 44325 49907
rect 33671 49751 34671 49797
rect 37896 49791 38556 49820
rect 37896 49745 37909 49791
rect 37955 49745 38026 49791
rect 38072 49745 38143 49791
rect 38189 49745 38261 49791
rect 38307 49745 38379 49791
rect 38425 49745 38497 49791
rect 38543 49745 38556 49791
rect 37896 49732 38556 49745
rect 39598 49791 39730 49820
rect 39598 49745 39641 49791
rect 39687 49745 39730 49791
rect 43695 49811 43739 49857
rect 43785 49811 43906 49857
rect 43952 49811 44071 49857
rect 44117 49811 44236 49857
rect 44282 49811 44325 49857
rect 50454 49843 51454 49875
rect 43695 49764 44325 49811
rect 39598 49732 39730 49745
rect 50454 49797 50516 49843
rect 50562 49797 50703 49843
rect 50749 49797 50890 49843
rect 50936 49797 51076 49843
rect 51122 49797 51263 49843
rect 51309 49797 51454 49843
rect 50454 49751 51454 49797
rect 33671 49457 34671 49503
rect 33671 49411 33816 49457
rect 33862 49411 34002 49457
rect 34048 49411 34189 49457
rect 34235 49411 34376 49457
rect 34422 49411 34562 49457
rect 34608 49411 34671 49457
rect 37896 49509 38556 49522
rect 37896 49463 37909 49509
rect 37955 49463 38026 49509
rect 38072 49463 38143 49509
rect 38189 49463 38261 49509
rect 38307 49463 38379 49509
rect 38425 49463 38497 49509
rect 38543 49463 38556 49509
rect 37896 49434 38556 49463
rect 39598 49509 39730 49522
rect 39598 49463 39641 49509
rect 39687 49463 39730 49509
rect 39598 49434 39730 49463
rect 43695 49443 44325 49490
rect 33671 49379 34671 49411
rect 33671 49198 34671 49259
rect 33671 49152 33684 49198
rect 33730 49152 33787 49198
rect 33833 49152 33890 49198
rect 33936 49152 33993 49198
rect 34039 49152 34096 49198
rect 34142 49152 34199 49198
rect 34245 49152 34302 49198
rect 34348 49152 34405 49198
rect 34451 49152 34508 49198
rect 34554 49152 34612 49198
rect 34658 49152 34671 49198
rect 33671 49123 34671 49152
rect 37896 49285 38556 49314
rect 37896 49239 37909 49285
rect 37955 49239 38026 49285
rect 38072 49239 38143 49285
rect 38189 49239 38261 49285
rect 38307 49239 38379 49285
rect 38425 49239 38497 49285
rect 38543 49239 38556 49285
rect 37896 49210 38556 49239
rect 43695 49397 43739 49443
rect 43785 49397 43906 49443
rect 43952 49397 44071 49443
rect 44117 49397 44236 49443
rect 44282 49397 44325 49443
rect 43695 49347 44325 49397
rect 50454 49457 51454 49503
rect 39598 49285 39730 49314
rect 39598 49239 39641 49285
rect 39687 49239 39730 49285
rect 39598 49226 39730 49239
rect 50454 49411 50516 49457
rect 50562 49411 50703 49457
rect 50749 49411 50890 49457
rect 50936 49411 51076 49457
rect 51122 49411 51263 49457
rect 51309 49411 51454 49457
rect 50454 49379 51454 49411
rect 43695 49123 44325 49227
rect 33671 48974 34671 49003
rect 37896 49061 38556 49090
rect 37896 49015 37909 49061
rect 37955 49015 38026 49061
rect 38072 49015 38143 49061
rect 38189 49015 38261 49061
rect 38307 49015 38379 49061
rect 38425 49015 38497 49061
rect 38543 49015 38556 49061
rect 37896 49002 38556 49015
rect 50454 49198 51454 49259
rect 50454 49152 50467 49198
rect 50513 49152 50571 49198
rect 50617 49152 50674 49198
rect 50720 49152 50777 49198
rect 50823 49152 50880 49198
rect 50926 49152 50983 49198
rect 51029 49152 51086 49198
rect 51132 49152 51189 49198
rect 51235 49152 51292 49198
rect 51338 49152 51395 49198
rect 51441 49152 51454 49198
rect 50454 49123 51454 49152
rect 33671 48928 33684 48974
rect 33730 48928 33787 48974
rect 33833 48928 33890 48974
rect 33936 48928 33993 48974
rect 34039 48928 34096 48974
rect 34142 48928 34199 48974
rect 34245 48928 34302 48974
rect 34348 48928 34405 48974
rect 34451 48928 34508 48974
rect 34554 48928 34612 48974
rect 34658 48928 34671 48974
rect 33671 48899 34671 48928
rect 39727 48974 40167 48987
rect 39727 48928 39740 48974
rect 39786 48928 39862 48974
rect 39908 48928 39985 48974
rect 40031 48928 40108 48974
rect 40154 48928 40167 48974
rect 39727 48899 40167 48928
rect 43695 48910 44325 49003
rect 50454 48974 51454 49003
rect 33671 48750 34671 48779
rect 33671 48704 33684 48750
rect 33730 48704 33787 48750
rect 33833 48704 33890 48750
rect 33936 48704 33993 48750
rect 34039 48704 34096 48750
rect 34142 48704 34199 48750
rect 34245 48704 34302 48750
rect 34348 48704 34405 48750
rect 34451 48704 34508 48750
rect 34554 48704 34612 48750
rect 34658 48704 34671 48750
rect 33671 48675 34671 48704
rect 39727 48750 40167 48779
rect 39727 48704 39740 48750
rect 39786 48704 39862 48750
rect 39908 48704 39985 48750
rect 40031 48704 40108 48750
rect 40154 48704 40167 48750
rect 39727 48675 40167 48704
rect 43695 48750 44325 48790
rect 50454 48928 50467 48974
rect 50513 48928 50571 48974
rect 50617 48928 50674 48974
rect 50720 48928 50777 48974
rect 50823 48928 50880 48974
rect 50926 48928 50983 48974
rect 51029 48928 51086 48974
rect 51132 48928 51189 48974
rect 51235 48928 51292 48974
rect 51338 48928 51395 48974
rect 51441 48928 51454 48974
rect 50454 48899 51454 48928
rect 43695 48704 43739 48750
rect 43785 48704 43906 48750
rect 43952 48704 44071 48750
rect 44117 48704 44236 48750
rect 44282 48704 44325 48750
rect 43695 48664 44325 48704
rect 33671 48526 34671 48555
rect 33671 48480 33684 48526
rect 33730 48480 33787 48526
rect 33833 48480 33890 48526
rect 33936 48480 33993 48526
rect 34039 48480 34096 48526
rect 34142 48480 34199 48526
rect 34245 48480 34302 48526
rect 34348 48480 34405 48526
rect 34451 48480 34508 48526
rect 34554 48480 34612 48526
rect 34658 48480 34671 48526
rect 33671 48451 34671 48480
rect 39727 48526 40167 48555
rect 39727 48480 39740 48526
rect 39786 48480 39862 48526
rect 39908 48480 39985 48526
rect 40031 48480 40108 48526
rect 40154 48480 40167 48526
rect 39727 48467 40167 48480
rect 50454 48750 51454 48779
rect 50454 48704 50467 48750
rect 50513 48704 50571 48750
rect 50617 48704 50674 48750
rect 50720 48704 50777 48750
rect 50823 48704 50880 48750
rect 50926 48704 50983 48750
rect 51029 48704 51086 48750
rect 51132 48704 51189 48750
rect 51235 48704 51292 48750
rect 51338 48704 51395 48750
rect 51441 48704 51454 48750
rect 50454 48675 51454 48704
rect 37896 48439 38556 48452
rect 43695 48451 44325 48544
rect 50454 48526 51454 48555
rect 50454 48480 50467 48526
rect 50513 48480 50571 48526
rect 50617 48480 50674 48526
rect 50720 48480 50777 48526
rect 50823 48480 50880 48526
rect 50926 48480 50983 48526
rect 51029 48480 51086 48526
rect 51132 48480 51189 48526
rect 51235 48480 51292 48526
rect 51338 48480 51395 48526
rect 51441 48480 51454 48526
rect 37896 48393 37909 48439
rect 37955 48393 38026 48439
rect 38072 48393 38143 48439
rect 38189 48393 38261 48439
rect 38307 48393 38379 48439
rect 38425 48393 38497 48439
rect 38543 48393 38556 48439
rect 37896 48364 38556 48393
rect 33671 48302 34671 48331
rect 33671 48256 33684 48302
rect 33730 48256 33787 48302
rect 33833 48256 33890 48302
rect 33936 48256 33993 48302
rect 34039 48256 34096 48302
rect 34142 48256 34199 48302
rect 34245 48256 34302 48302
rect 34348 48256 34405 48302
rect 34451 48256 34508 48302
rect 34554 48256 34612 48302
rect 34658 48256 34671 48302
rect 33671 48195 34671 48256
rect 33671 48043 34671 48075
rect 33671 47997 33816 48043
rect 33862 47997 34002 48043
rect 34048 47997 34189 48043
rect 34235 47997 34376 48043
rect 34422 47997 34562 48043
rect 34608 47997 34671 48043
rect 50454 48451 51454 48480
rect 37896 48215 38556 48244
rect 37896 48169 37909 48215
rect 37955 48169 38026 48215
rect 38072 48169 38143 48215
rect 38189 48169 38261 48215
rect 38307 48169 38379 48215
rect 38425 48169 38497 48215
rect 38543 48169 38556 48215
rect 37896 48140 38556 48169
rect 39598 48215 39730 48228
rect 43695 48227 44325 48331
rect 39598 48169 39641 48215
rect 39687 48169 39730 48215
rect 39598 48140 39730 48169
rect 50454 48302 51454 48331
rect 50454 48256 50467 48302
rect 50513 48256 50571 48302
rect 50617 48256 50674 48302
rect 50720 48256 50777 48302
rect 50823 48256 50880 48302
rect 50926 48256 50983 48302
rect 51029 48256 51086 48302
rect 51132 48256 51189 48302
rect 51235 48256 51292 48302
rect 51338 48256 51395 48302
rect 51441 48256 51454 48302
rect 50454 48195 51454 48256
rect 43695 48057 44325 48107
rect 33671 47951 34671 47997
rect 37896 47991 38556 48020
rect 37896 47945 37909 47991
rect 37955 47945 38026 47991
rect 38072 47945 38143 47991
rect 38189 47945 38261 47991
rect 38307 47945 38379 47991
rect 38425 47945 38497 47991
rect 38543 47945 38556 47991
rect 37896 47932 38556 47945
rect 39598 47991 39730 48020
rect 39598 47945 39641 47991
rect 39687 47945 39730 47991
rect 43695 48011 43739 48057
rect 43785 48011 43906 48057
rect 43952 48011 44071 48057
rect 44117 48011 44236 48057
rect 44282 48011 44325 48057
rect 50454 48043 51454 48075
rect 43695 47964 44325 48011
rect 39598 47932 39730 47945
rect 50454 47997 50516 48043
rect 50562 47997 50703 48043
rect 50749 47997 50890 48043
rect 50936 47997 51076 48043
rect 51122 47997 51263 48043
rect 51309 47997 51454 48043
rect 50454 47951 51454 47997
rect 33671 47657 34671 47703
rect 33671 47611 33816 47657
rect 33862 47611 34002 47657
rect 34048 47611 34189 47657
rect 34235 47611 34376 47657
rect 34422 47611 34562 47657
rect 34608 47611 34671 47657
rect 37896 47709 38556 47722
rect 37896 47663 37909 47709
rect 37955 47663 38026 47709
rect 38072 47663 38143 47709
rect 38189 47663 38261 47709
rect 38307 47663 38379 47709
rect 38425 47663 38497 47709
rect 38543 47663 38556 47709
rect 37896 47634 38556 47663
rect 39598 47709 39730 47722
rect 39598 47663 39641 47709
rect 39687 47663 39730 47709
rect 39598 47634 39730 47663
rect 43695 47643 44325 47690
rect 33671 47579 34671 47611
rect 33671 47398 34671 47459
rect 33671 47352 33684 47398
rect 33730 47352 33787 47398
rect 33833 47352 33890 47398
rect 33936 47352 33993 47398
rect 34039 47352 34096 47398
rect 34142 47352 34199 47398
rect 34245 47352 34302 47398
rect 34348 47352 34405 47398
rect 34451 47352 34508 47398
rect 34554 47352 34612 47398
rect 34658 47352 34671 47398
rect 33671 47323 34671 47352
rect 37896 47485 38556 47514
rect 37896 47439 37909 47485
rect 37955 47439 38026 47485
rect 38072 47439 38143 47485
rect 38189 47439 38261 47485
rect 38307 47439 38379 47485
rect 38425 47439 38497 47485
rect 38543 47439 38556 47485
rect 37896 47410 38556 47439
rect 43695 47597 43739 47643
rect 43785 47597 43906 47643
rect 43952 47597 44071 47643
rect 44117 47597 44236 47643
rect 44282 47597 44325 47643
rect 43695 47547 44325 47597
rect 50454 47657 51454 47703
rect 39598 47485 39730 47514
rect 39598 47439 39641 47485
rect 39687 47439 39730 47485
rect 39598 47426 39730 47439
rect 50454 47611 50516 47657
rect 50562 47611 50703 47657
rect 50749 47611 50890 47657
rect 50936 47611 51076 47657
rect 51122 47611 51263 47657
rect 51309 47611 51454 47657
rect 50454 47579 51454 47611
rect 43695 47323 44325 47427
rect 33671 47174 34671 47203
rect 37896 47261 38556 47290
rect 37896 47215 37909 47261
rect 37955 47215 38026 47261
rect 38072 47215 38143 47261
rect 38189 47215 38261 47261
rect 38307 47215 38379 47261
rect 38425 47215 38497 47261
rect 38543 47215 38556 47261
rect 37896 47202 38556 47215
rect 50454 47398 51454 47459
rect 50454 47352 50467 47398
rect 50513 47352 50571 47398
rect 50617 47352 50674 47398
rect 50720 47352 50777 47398
rect 50823 47352 50880 47398
rect 50926 47352 50983 47398
rect 51029 47352 51086 47398
rect 51132 47352 51189 47398
rect 51235 47352 51292 47398
rect 51338 47352 51395 47398
rect 51441 47352 51454 47398
rect 50454 47323 51454 47352
rect 33671 47128 33684 47174
rect 33730 47128 33787 47174
rect 33833 47128 33890 47174
rect 33936 47128 33993 47174
rect 34039 47128 34096 47174
rect 34142 47128 34199 47174
rect 34245 47128 34302 47174
rect 34348 47128 34405 47174
rect 34451 47128 34508 47174
rect 34554 47128 34612 47174
rect 34658 47128 34671 47174
rect 33671 47099 34671 47128
rect 39727 47174 40167 47187
rect 39727 47128 39740 47174
rect 39786 47128 39862 47174
rect 39908 47128 39985 47174
rect 40031 47128 40108 47174
rect 40154 47128 40167 47174
rect 39727 47099 40167 47128
rect 43695 47110 44325 47203
rect 50454 47174 51454 47203
rect 33671 46950 34671 46979
rect 33671 46904 33684 46950
rect 33730 46904 33787 46950
rect 33833 46904 33890 46950
rect 33936 46904 33993 46950
rect 34039 46904 34096 46950
rect 34142 46904 34199 46950
rect 34245 46904 34302 46950
rect 34348 46904 34405 46950
rect 34451 46904 34508 46950
rect 34554 46904 34612 46950
rect 34658 46904 34671 46950
rect 33671 46875 34671 46904
rect 39727 46950 40167 46979
rect 39727 46904 39740 46950
rect 39786 46904 39862 46950
rect 39908 46904 39985 46950
rect 40031 46904 40108 46950
rect 40154 46904 40167 46950
rect 39727 46875 40167 46904
rect 43695 46950 44325 46990
rect 50454 47128 50467 47174
rect 50513 47128 50571 47174
rect 50617 47128 50674 47174
rect 50720 47128 50777 47174
rect 50823 47128 50880 47174
rect 50926 47128 50983 47174
rect 51029 47128 51086 47174
rect 51132 47128 51189 47174
rect 51235 47128 51292 47174
rect 51338 47128 51395 47174
rect 51441 47128 51454 47174
rect 50454 47099 51454 47128
rect 43695 46904 43739 46950
rect 43785 46904 43906 46950
rect 43952 46904 44071 46950
rect 44117 46904 44236 46950
rect 44282 46904 44325 46950
rect 43695 46864 44325 46904
rect 33671 46726 34671 46755
rect 33671 46680 33684 46726
rect 33730 46680 33787 46726
rect 33833 46680 33890 46726
rect 33936 46680 33993 46726
rect 34039 46680 34096 46726
rect 34142 46680 34199 46726
rect 34245 46680 34302 46726
rect 34348 46680 34405 46726
rect 34451 46680 34508 46726
rect 34554 46680 34612 46726
rect 34658 46680 34671 46726
rect 33671 46651 34671 46680
rect 39727 46726 40167 46755
rect 39727 46680 39740 46726
rect 39786 46680 39862 46726
rect 39908 46680 39985 46726
rect 40031 46680 40108 46726
rect 40154 46680 40167 46726
rect 39727 46667 40167 46680
rect 50454 46950 51454 46979
rect 50454 46904 50467 46950
rect 50513 46904 50571 46950
rect 50617 46904 50674 46950
rect 50720 46904 50777 46950
rect 50823 46904 50880 46950
rect 50926 46904 50983 46950
rect 51029 46904 51086 46950
rect 51132 46904 51189 46950
rect 51235 46904 51292 46950
rect 51338 46904 51395 46950
rect 51441 46904 51454 46950
rect 50454 46875 51454 46904
rect 37896 46639 38556 46652
rect 43695 46651 44325 46744
rect 50454 46726 51454 46755
rect 50454 46680 50467 46726
rect 50513 46680 50571 46726
rect 50617 46680 50674 46726
rect 50720 46680 50777 46726
rect 50823 46680 50880 46726
rect 50926 46680 50983 46726
rect 51029 46680 51086 46726
rect 51132 46680 51189 46726
rect 51235 46680 51292 46726
rect 51338 46680 51395 46726
rect 51441 46680 51454 46726
rect 37896 46593 37909 46639
rect 37955 46593 38026 46639
rect 38072 46593 38143 46639
rect 38189 46593 38261 46639
rect 38307 46593 38379 46639
rect 38425 46593 38497 46639
rect 38543 46593 38556 46639
rect 37896 46564 38556 46593
rect 33671 46502 34671 46531
rect 33671 46456 33684 46502
rect 33730 46456 33787 46502
rect 33833 46456 33890 46502
rect 33936 46456 33993 46502
rect 34039 46456 34096 46502
rect 34142 46456 34199 46502
rect 34245 46456 34302 46502
rect 34348 46456 34405 46502
rect 34451 46456 34508 46502
rect 34554 46456 34612 46502
rect 34658 46456 34671 46502
rect 33671 46395 34671 46456
rect 33671 46243 34671 46275
rect 33671 46197 33816 46243
rect 33862 46197 34002 46243
rect 34048 46197 34189 46243
rect 34235 46197 34376 46243
rect 34422 46197 34562 46243
rect 34608 46197 34671 46243
rect 50454 46651 51454 46680
rect 37896 46415 38556 46444
rect 37896 46369 37909 46415
rect 37955 46369 38026 46415
rect 38072 46369 38143 46415
rect 38189 46369 38261 46415
rect 38307 46369 38379 46415
rect 38425 46369 38497 46415
rect 38543 46369 38556 46415
rect 37896 46340 38556 46369
rect 39598 46415 39730 46428
rect 43695 46427 44325 46531
rect 39598 46369 39641 46415
rect 39687 46369 39730 46415
rect 39598 46340 39730 46369
rect 50454 46502 51454 46531
rect 50454 46456 50467 46502
rect 50513 46456 50571 46502
rect 50617 46456 50674 46502
rect 50720 46456 50777 46502
rect 50823 46456 50880 46502
rect 50926 46456 50983 46502
rect 51029 46456 51086 46502
rect 51132 46456 51189 46502
rect 51235 46456 51292 46502
rect 51338 46456 51395 46502
rect 51441 46456 51454 46502
rect 50454 46395 51454 46456
rect 43695 46257 44325 46307
rect 33671 46151 34671 46197
rect 37896 46191 38556 46220
rect 37896 46145 37909 46191
rect 37955 46145 38026 46191
rect 38072 46145 38143 46191
rect 38189 46145 38261 46191
rect 38307 46145 38379 46191
rect 38425 46145 38497 46191
rect 38543 46145 38556 46191
rect 37896 46132 38556 46145
rect 39598 46191 39730 46220
rect 39598 46145 39641 46191
rect 39687 46145 39730 46191
rect 43695 46211 43739 46257
rect 43785 46211 43906 46257
rect 43952 46211 44071 46257
rect 44117 46211 44236 46257
rect 44282 46211 44325 46257
rect 50454 46243 51454 46275
rect 43695 46164 44325 46211
rect 39598 46132 39730 46145
rect 50454 46197 50516 46243
rect 50562 46197 50703 46243
rect 50749 46197 50890 46243
rect 50936 46197 51076 46243
rect 51122 46197 51263 46243
rect 51309 46197 51454 46243
rect 50454 46151 51454 46197
rect 33671 45857 34671 45903
rect 33671 45811 33816 45857
rect 33862 45811 34002 45857
rect 34048 45811 34189 45857
rect 34235 45811 34376 45857
rect 34422 45811 34562 45857
rect 34608 45811 34671 45857
rect 37896 45909 38556 45922
rect 37896 45863 37909 45909
rect 37955 45863 38026 45909
rect 38072 45863 38143 45909
rect 38189 45863 38261 45909
rect 38307 45863 38379 45909
rect 38425 45863 38497 45909
rect 38543 45863 38556 45909
rect 37896 45834 38556 45863
rect 39598 45909 39730 45922
rect 39598 45863 39641 45909
rect 39687 45863 39730 45909
rect 39598 45834 39730 45863
rect 43695 45843 44325 45890
rect 33671 45779 34671 45811
rect 33671 45598 34671 45659
rect 33671 45552 33684 45598
rect 33730 45552 33787 45598
rect 33833 45552 33890 45598
rect 33936 45552 33993 45598
rect 34039 45552 34096 45598
rect 34142 45552 34199 45598
rect 34245 45552 34302 45598
rect 34348 45552 34405 45598
rect 34451 45552 34508 45598
rect 34554 45552 34612 45598
rect 34658 45552 34671 45598
rect 33671 45523 34671 45552
rect 37896 45685 38556 45714
rect 37896 45639 37909 45685
rect 37955 45639 38026 45685
rect 38072 45639 38143 45685
rect 38189 45639 38261 45685
rect 38307 45639 38379 45685
rect 38425 45639 38497 45685
rect 38543 45639 38556 45685
rect 37896 45610 38556 45639
rect 43695 45797 43739 45843
rect 43785 45797 43906 45843
rect 43952 45797 44071 45843
rect 44117 45797 44236 45843
rect 44282 45797 44325 45843
rect 43695 45747 44325 45797
rect 50454 45857 51454 45903
rect 39598 45685 39730 45714
rect 39598 45639 39641 45685
rect 39687 45639 39730 45685
rect 39598 45626 39730 45639
rect 50454 45811 50516 45857
rect 50562 45811 50703 45857
rect 50749 45811 50890 45857
rect 50936 45811 51076 45857
rect 51122 45811 51263 45857
rect 51309 45811 51454 45857
rect 50454 45779 51454 45811
rect 43695 45523 44325 45627
rect 33671 45374 34671 45403
rect 37896 45461 38556 45490
rect 37896 45415 37909 45461
rect 37955 45415 38026 45461
rect 38072 45415 38143 45461
rect 38189 45415 38261 45461
rect 38307 45415 38379 45461
rect 38425 45415 38497 45461
rect 38543 45415 38556 45461
rect 37896 45402 38556 45415
rect 50454 45598 51454 45659
rect 50454 45552 50467 45598
rect 50513 45552 50571 45598
rect 50617 45552 50674 45598
rect 50720 45552 50777 45598
rect 50823 45552 50880 45598
rect 50926 45552 50983 45598
rect 51029 45552 51086 45598
rect 51132 45552 51189 45598
rect 51235 45552 51292 45598
rect 51338 45552 51395 45598
rect 51441 45552 51454 45598
rect 50454 45523 51454 45552
rect 33671 45328 33684 45374
rect 33730 45328 33787 45374
rect 33833 45328 33890 45374
rect 33936 45328 33993 45374
rect 34039 45328 34096 45374
rect 34142 45328 34199 45374
rect 34245 45328 34302 45374
rect 34348 45328 34405 45374
rect 34451 45328 34508 45374
rect 34554 45328 34612 45374
rect 34658 45328 34671 45374
rect 33671 45299 34671 45328
rect 39727 45374 40167 45387
rect 39727 45328 39740 45374
rect 39786 45328 39862 45374
rect 39908 45328 39985 45374
rect 40031 45328 40108 45374
rect 40154 45328 40167 45374
rect 39727 45299 40167 45328
rect 43695 45310 44325 45403
rect 50454 45374 51454 45403
rect 33671 45150 34671 45179
rect 33671 45104 33684 45150
rect 33730 45104 33787 45150
rect 33833 45104 33890 45150
rect 33936 45104 33993 45150
rect 34039 45104 34096 45150
rect 34142 45104 34199 45150
rect 34245 45104 34302 45150
rect 34348 45104 34405 45150
rect 34451 45104 34508 45150
rect 34554 45104 34612 45150
rect 34658 45104 34671 45150
rect 33671 45075 34671 45104
rect 39727 45150 40167 45179
rect 39727 45104 39740 45150
rect 39786 45104 39862 45150
rect 39908 45104 39985 45150
rect 40031 45104 40108 45150
rect 40154 45104 40167 45150
rect 39727 45075 40167 45104
rect 43695 45150 44325 45190
rect 50454 45328 50467 45374
rect 50513 45328 50571 45374
rect 50617 45328 50674 45374
rect 50720 45328 50777 45374
rect 50823 45328 50880 45374
rect 50926 45328 50983 45374
rect 51029 45328 51086 45374
rect 51132 45328 51189 45374
rect 51235 45328 51292 45374
rect 51338 45328 51395 45374
rect 51441 45328 51454 45374
rect 50454 45299 51454 45328
rect 43695 45104 43739 45150
rect 43785 45104 43906 45150
rect 43952 45104 44071 45150
rect 44117 45104 44236 45150
rect 44282 45104 44325 45150
rect 43695 45064 44325 45104
rect 33671 44926 34671 44955
rect 33671 44880 33684 44926
rect 33730 44880 33787 44926
rect 33833 44880 33890 44926
rect 33936 44880 33993 44926
rect 34039 44880 34096 44926
rect 34142 44880 34199 44926
rect 34245 44880 34302 44926
rect 34348 44880 34405 44926
rect 34451 44880 34508 44926
rect 34554 44880 34612 44926
rect 34658 44880 34671 44926
rect 33671 44851 34671 44880
rect 39727 44926 40167 44955
rect 39727 44880 39740 44926
rect 39786 44880 39862 44926
rect 39908 44880 39985 44926
rect 40031 44880 40108 44926
rect 40154 44880 40167 44926
rect 39727 44867 40167 44880
rect 50454 45150 51454 45179
rect 50454 45104 50467 45150
rect 50513 45104 50571 45150
rect 50617 45104 50674 45150
rect 50720 45104 50777 45150
rect 50823 45104 50880 45150
rect 50926 45104 50983 45150
rect 51029 45104 51086 45150
rect 51132 45104 51189 45150
rect 51235 45104 51292 45150
rect 51338 45104 51395 45150
rect 51441 45104 51454 45150
rect 50454 45075 51454 45104
rect 37896 44839 38556 44852
rect 43695 44851 44325 44944
rect 50454 44926 51454 44955
rect 50454 44880 50467 44926
rect 50513 44880 50571 44926
rect 50617 44880 50674 44926
rect 50720 44880 50777 44926
rect 50823 44880 50880 44926
rect 50926 44880 50983 44926
rect 51029 44880 51086 44926
rect 51132 44880 51189 44926
rect 51235 44880 51292 44926
rect 51338 44880 51395 44926
rect 51441 44880 51454 44926
rect 37896 44793 37909 44839
rect 37955 44793 38026 44839
rect 38072 44793 38143 44839
rect 38189 44793 38261 44839
rect 38307 44793 38379 44839
rect 38425 44793 38497 44839
rect 38543 44793 38556 44839
rect 37896 44764 38556 44793
rect 33671 44702 34671 44731
rect 33671 44656 33684 44702
rect 33730 44656 33787 44702
rect 33833 44656 33890 44702
rect 33936 44656 33993 44702
rect 34039 44656 34096 44702
rect 34142 44656 34199 44702
rect 34245 44656 34302 44702
rect 34348 44656 34405 44702
rect 34451 44656 34508 44702
rect 34554 44656 34612 44702
rect 34658 44656 34671 44702
rect 33671 44595 34671 44656
rect 33671 44443 34671 44475
rect 33671 44397 33816 44443
rect 33862 44397 34002 44443
rect 34048 44397 34189 44443
rect 34235 44397 34376 44443
rect 34422 44397 34562 44443
rect 34608 44397 34671 44443
rect 50454 44851 51454 44880
rect 37896 44615 38556 44644
rect 37896 44569 37909 44615
rect 37955 44569 38026 44615
rect 38072 44569 38143 44615
rect 38189 44569 38261 44615
rect 38307 44569 38379 44615
rect 38425 44569 38497 44615
rect 38543 44569 38556 44615
rect 37896 44540 38556 44569
rect 39598 44615 39730 44628
rect 43695 44627 44325 44731
rect 39598 44569 39641 44615
rect 39687 44569 39730 44615
rect 39598 44540 39730 44569
rect 50454 44702 51454 44731
rect 50454 44656 50467 44702
rect 50513 44656 50571 44702
rect 50617 44656 50674 44702
rect 50720 44656 50777 44702
rect 50823 44656 50880 44702
rect 50926 44656 50983 44702
rect 51029 44656 51086 44702
rect 51132 44656 51189 44702
rect 51235 44656 51292 44702
rect 51338 44656 51395 44702
rect 51441 44656 51454 44702
rect 50454 44595 51454 44656
rect 43695 44457 44325 44507
rect 33671 44351 34671 44397
rect 37896 44391 38556 44420
rect 37896 44345 37909 44391
rect 37955 44345 38026 44391
rect 38072 44345 38143 44391
rect 38189 44345 38261 44391
rect 38307 44345 38379 44391
rect 38425 44345 38497 44391
rect 38543 44345 38556 44391
rect 37896 44332 38556 44345
rect 39598 44391 39730 44420
rect 39598 44345 39641 44391
rect 39687 44345 39730 44391
rect 43695 44411 43739 44457
rect 43785 44411 43906 44457
rect 43952 44411 44071 44457
rect 44117 44411 44236 44457
rect 44282 44411 44325 44457
rect 50454 44443 51454 44475
rect 43695 44364 44325 44411
rect 39598 44332 39730 44345
rect 50454 44397 50516 44443
rect 50562 44397 50703 44443
rect 50749 44397 50890 44443
rect 50936 44397 51076 44443
rect 51122 44397 51263 44443
rect 51309 44397 51454 44443
rect 50454 44351 51454 44397
rect 33671 44057 34671 44103
rect 33671 44011 33816 44057
rect 33862 44011 34002 44057
rect 34048 44011 34189 44057
rect 34235 44011 34376 44057
rect 34422 44011 34562 44057
rect 34608 44011 34671 44057
rect 37896 44109 38556 44122
rect 37896 44063 37909 44109
rect 37955 44063 38026 44109
rect 38072 44063 38143 44109
rect 38189 44063 38261 44109
rect 38307 44063 38379 44109
rect 38425 44063 38497 44109
rect 38543 44063 38556 44109
rect 37896 44034 38556 44063
rect 39598 44109 39730 44122
rect 39598 44063 39641 44109
rect 39687 44063 39730 44109
rect 39598 44034 39730 44063
rect 43695 44043 44325 44090
rect 33671 43979 34671 44011
rect 33671 43798 34671 43859
rect 33671 43752 33684 43798
rect 33730 43752 33787 43798
rect 33833 43752 33890 43798
rect 33936 43752 33993 43798
rect 34039 43752 34096 43798
rect 34142 43752 34199 43798
rect 34245 43752 34302 43798
rect 34348 43752 34405 43798
rect 34451 43752 34508 43798
rect 34554 43752 34612 43798
rect 34658 43752 34671 43798
rect 33671 43723 34671 43752
rect 37896 43885 38556 43914
rect 37896 43839 37909 43885
rect 37955 43839 38026 43885
rect 38072 43839 38143 43885
rect 38189 43839 38261 43885
rect 38307 43839 38379 43885
rect 38425 43839 38497 43885
rect 38543 43839 38556 43885
rect 37896 43810 38556 43839
rect 43695 43997 43739 44043
rect 43785 43997 43906 44043
rect 43952 43997 44071 44043
rect 44117 43997 44236 44043
rect 44282 43997 44325 44043
rect 43695 43947 44325 43997
rect 50454 44057 51454 44103
rect 39598 43885 39730 43914
rect 39598 43839 39641 43885
rect 39687 43839 39730 43885
rect 39598 43826 39730 43839
rect 50454 44011 50516 44057
rect 50562 44011 50703 44057
rect 50749 44011 50890 44057
rect 50936 44011 51076 44057
rect 51122 44011 51263 44057
rect 51309 44011 51454 44057
rect 50454 43979 51454 44011
rect 43695 43723 44325 43827
rect 33671 43574 34671 43603
rect 37896 43661 38556 43690
rect 37896 43615 37909 43661
rect 37955 43615 38026 43661
rect 38072 43615 38143 43661
rect 38189 43615 38261 43661
rect 38307 43615 38379 43661
rect 38425 43615 38497 43661
rect 38543 43615 38556 43661
rect 37896 43602 38556 43615
rect 50454 43798 51454 43859
rect 50454 43752 50467 43798
rect 50513 43752 50571 43798
rect 50617 43752 50674 43798
rect 50720 43752 50777 43798
rect 50823 43752 50880 43798
rect 50926 43752 50983 43798
rect 51029 43752 51086 43798
rect 51132 43752 51189 43798
rect 51235 43752 51292 43798
rect 51338 43752 51395 43798
rect 51441 43752 51454 43798
rect 50454 43723 51454 43752
rect 33671 43528 33684 43574
rect 33730 43528 33787 43574
rect 33833 43528 33890 43574
rect 33936 43528 33993 43574
rect 34039 43528 34096 43574
rect 34142 43528 34199 43574
rect 34245 43528 34302 43574
rect 34348 43528 34405 43574
rect 34451 43528 34508 43574
rect 34554 43528 34612 43574
rect 34658 43528 34671 43574
rect 33671 43499 34671 43528
rect 39727 43574 40167 43587
rect 39727 43528 39740 43574
rect 39786 43528 39862 43574
rect 39908 43528 39985 43574
rect 40031 43528 40108 43574
rect 40154 43528 40167 43574
rect 39727 43499 40167 43528
rect 43695 43510 44325 43603
rect 50454 43574 51454 43603
rect 33671 43350 34671 43379
rect 33671 43304 33684 43350
rect 33730 43304 33787 43350
rect 33833 43304 33890 43350
rect 33936 43304 33993 43350
rect 34039 43304 34096 43350
rect 34142 43304 34199 43350
rect 34245 43304 34302 43350
rect 34348 43304 34405 43350
rect 34451 43304 34508 43350
rect 34554 43304 34612 43350
rect 34658 43304 34671 43350
rect 33671 43275 34671 43304
rect 39727 43350 40167 43379
rect 39727 43304 39740 43350
rect 39786 43304 39862 43350
rect 39908 43304 39985 43350
rect 40031 43304 40108 43350
rect 40154 43304 40167 43350
rect 39727 43275 40167 43304
rect 43695 43350 44325 43390
rect 50454 43528 50467 43574
rect 50513 43528 50571 43574
rect 50617 43528 50674 43574
rect 50720 43528 50777 43574
rect 50823 43528 50880 43574
rect 50926 43528 50983 43574
rect 51029 43528 51086 43574
rect 51132 43528 51189 43574
rect 51235 43528 51292 43574
rect 51338 43528 51395 43574
rect 51441 43528 51454 43574
rect 50454 43499 51454 43528
rect 43695 43304 43739 43350
rect 43785 43304 43906 43350
rect 43952 43304 44071 43350
rect 44117 43304 44236 43350
rect 44282 43304 44325 43350
rect 43695 43264 44325 43304
rect 33671 43126 34671 43155
rect 33671 43080 33684 43126
rect 33730 43080 33787 43126
rect 33833 43080 33890 43126
rect 33936 43080 33993 43126
rect 34039 43080 34096 43126
rect 34142 43080 34199 43126
rect 34245 43080 34302 43126
rect 34348 43080 34405 43126
rect 34451 43080 34508 43126
rect 34554 43080 34612 43126
rect 34658 43080 34671 43126
rect 33671 43051 34671 43080
rect 39727 43126 40167 43155
rect 39727 43080 39740 43126
rect 39786 43080 39862 43126
rect 39908 43080 39985 43126
rect 40031 43080 40108 43126
rect 40154 43080 40167 43126
rect 39727 43067 40167 43080
rect 50454 43350 51454 43379
rect 50454 43304 50467 43350
rect 50513 43304 50571 43350
rect 50617 43304 50674 43350
rect 50720 43304 50777 43350
rect 50823 43304 50880 43350
rect 50926 43304 50983 43350
rect 51029 43304 51086 43350
rect 51132 43304 51189 43350
rect 51235 43304 51292 43350
rect 51338 43304 51395 43350
rect 51441 43304 51454 43350
rect 50454 43275 51454 43304
rect 37896 43039 38556 43052
rect 43695 43051 44325 43144
rect 50454 43126 51454 43155
rect 50454 43080 50467 43126
rect 50513 43080 50571 43126
rect 50617 43080 50674 43126
rect 50720 43080 50777 43126
rect 50823 43080 50880 43126
rect 50926 43080 50983 43126
rect 51029 43080 51086 43126
rect 51132 43080 51189 43126
rect 51235 43080 51292 43126
rect 51338 43080 51395 43126
rect 51441 43080 51454 43126
rect 37896 42993 37909 43039
rect 37955 42993 38026 43039
rect 38072 42993 38143 43039
rect 38189 42993 38261 43039
rect 38307 42993 38379 43039
rect 38425 42993 38497 43039
rect 38543 42993 38556 43039
rect 37896 42964 38556 42993
rect 33671 42902 34671 42931
rect 33671 42856 33684 42902
rect 33730 42856 33787 42902
rect 33833 42856 33890 42902
rect 33936 42856 33993 42902
rect 34039 42856 34096 42902
rect 34142 42856 34199 42902
rect 34245 42856 34302 42902
rect 34348 42856 34405 42902
rect 34451 42856 34508 42902
rect 34554 42856 34612 42902
rect 34658 42856 34671 42902
rect 33671 42795 34671 42856
rect 33671 42643 34671 42675
rect 33671 42597 33816 42643
rect 33862 42597 34002 42643
rect 34048 42597 34189 42643
rect 34235 42597 34376 42643
rect 34422 42597 34562 42643
rect 34608 42597 34671 42643
rect 50454 43051 51454 43080
rect 37896 42815 38556 42844
rect 37896 42769 37909 42815
rect 37955 42769 38026 42815
rect 38072 42769 38143 42815
rect 38189 42769 38261 42815
rect 38307 42769 38379 42815
rect 38425 42769 38497 42815
rect 38543 42769 38556 42815
rect 37896 42740 38556 42769
rect 39598 42815 39730 42828
rect 43695 42827 44325 42931
rect 39598 42769 39641 42815
rect 39687 42769 39730 42815
rect 39598 42740 39730 42769
rect 50454 42902 51454 42931
rect 50454 42856 50467 42902
rect 50513 42856 50571 42902
rect 50617 42856 50674 42902
rect 50720 42856 50777 42902
rect 50823 42856 50880 42902
rect 50926 42856 50983 42902
rect 51029 42856 51086 42902
rect 51132 42856 51189 42902
rect 51235 42856 51292 42902
rect 51338 42856 51395 42902
rect 51441 42856 51454 42902
rect 50454 42795 51454 42856
rect 43695 42657 44325 42707
rect 33671 42551 34671 42597
rect 37896 42591 38556 42620
rect 37896 42545 37909 42591
rect 37955 42545 38026 42591
rect 38072 42545 38143 42591
rect 38189 42545 38261 42591
rect 38307 42545 38379 42591
rect 38425 42545 38497 42591
rect 38543 42545 38556 42591
rect 37896 42532 38556 42545
rect 39598 42591 39730 42620
rect 39598 42545 39641 42591
rect 39687 42545 39730 42591
rect 43695 42611 43739 42657
rect 43785 42611 43906 42657
rect 43952 42611 44071 42657
rect 44117 42611 44236 42657
rect 44282 42611 44325 42657
rect 50454 42643 51454 42675
rect 43695 42564 44325 42611
rect 39598 42532 39730 42545
rect 50454 42597 50516 42643
rect 50562 42597 50703 42643
rect 50749 42597 50890 42643
rect 50936 42597 51076 42643
rect 51122 42597 51263 42643
rect 51309 42597 51454 42643
rect 50454 42551 51454 42597
rect 33671 42257 34671 42303
rect 33671 42211 33816 42257
rect 33862 42211 34002 42257
rect 34048 42211 34189 42257
rect 34235 42211 34376 42257
rect 34422 42211 34562 42257
rect 34608 42211 34671 42257
rect 37896 42309 38556 42322
rect 37896 42263 37909 42309
rect 37955 42263 38026 42309
rect 38072 42263 38143 42309
rect 38189 42263 38261 42309
rect 38307 42263 38379 42309
rect 38425 42263 38497 42309
rect 38543 42263 38556 42309
rect 37896 42234 38556 42263
rect 39598 42309 39730 42322
rect 39598 42263 39641 42309
rect 39687 42263 39730 42309
rect 39598 42234 39730 42263
rect 43695 42243 44325 42290
rect 33671 42179 34671 42211
rect 33671 41998 34671 42059
rect 33671 41952 33684 41998
rect 33730 41952 33787 41998
rect 33833 41952 33890 41998
rect 33936 41952 33993 41998
rect 34039 41952 34096 41998
rect 34142 41952 34199 41998
rect 34245 41952 34302 41998
rect 34348 41952 34405 41998
rect 34451 41952 34508 41998
rect 34554 41952 34612 41998
rect 34658 41952 34671 41998
rect 33671 41923 34671 41952
rect 37896 42085 38556 42114
rect 37896 42039 37909 42085
rect 37955 42039 38026 42085
rect 38072 42039 38143 42085
rect 38189 42039 38261 42085
rect 38307 42039 38379 42085
rect 38425 42039 38497 42085
rect 38543 42039 38556 42085
rect 37896 42010 38556 42039
rect 43695 42197 43739 42243
rect 43785 42197 43906 42243
rect 43952 42197 44071 42243
rect 44117 42197 44236 42243
rect 44282 42197 44325 42243
rect 43695 42147 44325 42197
rect 50454 42257 51454 42303
rect 39598 42085 39730 42114
rect 39598 42039 39641 42085
rect 39687 42039 39730 42085
rect 39598 42026 39730 42039
rect 50454 42211 50516 42257
rect 50562 42211 50703 42257
rect 50749 42211 50890 42257
rect 50936 42211 51076 42257
rect 51122 42211 51263 42257
rect 51309 42211 51454 42257
rect 50454 42179 51454 42211
rect 43695 41923 44325 42027
rect 33671 41774 34671 41803
rect 37896 41861 38556 41890
rect 37896 41815 37909 41861
rect 37955 41815 38026 41861
rect 38072 41815 38143 41861
rect 38189 41815 38261 41861
rect 38307 41815 38379 41861
rect 38425 41815 38497 41861
rect 38543 41815 38556 41861
rect 37896 41802 38556 41815
rect 50454 41998 51454 42059
rect 50454 41952 50467 41998
rect 50513 41952 50571 41998
rect 50617 41952 50674 41998
rect 50720 41952 50777 41998
rect 50823 41952 50880 41998
rect 50926 41952 50983 41998
rect 51029 41952 51086 41998
rect 51132 41952 51189 41998
rect 51235 41952 51292 41998
rect 51338 41952 51395 41998
rect 51441 41952 51454 41998
rect 50454 41923 51454 41952
rect 33671 41728 33684 41774
rect 33730 41728 33787 41774
rect 33833 41728 33890 41774
rect 33936 41728 33993 41774
rect 34039 41728 34096 41774
rect 34142 41728 34199 41774
rect 34245 41728 34302 41774
rect 34348 41728 34405 41774
rect 34451 41728 34508 41774
rect 34554 41728 34612 41774
rect 34658 41728 34671 41774
rect 33671 41699 34671 41728
rect 39727 41774 40167 41787
rect 39727 41728 39740 41774
rect 39786 41728 39862 41774
rect 39908 41728 39985 41774
rect 40031 41728 40108 41774
rect 40154 41728 40167 41774
rect 39727 41699 40167 41728
rect 43695 41710 44325 41803
rect 50454 41774 51454 41803
rect 33671 41550 34671 41579
rect 33671 41504 33684 41550
rect 33730 41504 33787 41550
rect 33833 41504 33890 41550
rect 33936 41504 33993 41550
rect 34039 41504 34096 41550
rect 34142 41504 34199 41550
rect 34245 41504 34302 41550
rect 34348 41504 34405 41550
rect 34451 41504 34508 41550
rect 34554 41504 34612 41550
rect 34658 41504 34671 41550
rect 33671 41475 34671 41504
rect 39727 41550 40167 41579
rect 39727 41504 39740 41550
rect 39786 41504 39862 41550
rect 39908 41504 39985 41550
rect 40031 41504 40108 41550
rect 40154 41504 40167 41550
rect 39727 41475 40167 41504
rect 43695 41550 44325 41590
rect 50454 41728 50467 41774
rect 50513 41728 50571 41774
rect 50617 41728 50674 41774
rect 50720 41728 50777 41774
rect 50823 41728 50880 41774
rect 50926 41728 50983 41774
rect 51029 41728 51086 41774
rect 51132 41728 51189 41774
rect 51235 41728 51292 41774
rect 51338 41728 51395 41774
rect 51441 41728 51454 41774
rect 50454 41699 51454 41728
rect 43695 41504 43739 41550
rect 43785 41504 43906 41550
rect 43952 41504 44071 41550
rect 44117 41504 44236 41550
rect 44282 41504 44325 41550
rect 43695 41464 44325 41504
rect 33671 41326 34671 41355
rect 33671 41280 33684 41326
rect 33730 41280 33787 41326
rect 33833 41280 33890 41326
rect 33936 41280 33993 41326
rect 34039 41280 34096 41326
rect 34142 41280 34199 41326
rect 34245 41280 34302 41326
rect 34348 41280 34405 41326
rect 34451 41280 34508 41326
rect 34554 41280 34612 41326
rect 34658 41280 34671 41326
rect 33671 41251 34671 41280
rect 39727 41326 40167 41355
rect 39727 41280 39740 41326
rect 39786 41280 39862 41326
rect 39908 41280 39985 41326
rect 40031 41280 40108 41326
rect 40154 41280 40167 41326
rect 39727 41267 40167 41280
rect 50454 41550 51454 41579
rect 50454 41504 50467 41550
rect 50513 41504 50571 41550
rect 50617 41504 50674 41550
rect 50720 41504 50777 41550
rect 50823 41504 50880 41550
rect 50926 41504 50983 41550
rect 51029 41504 51086 41550
rect 51132 41504 51189 41550
rect 51235 41504 51292 41550
rect 51338 41504 51395 41550
rect 51441 41504 51454 41550
rect 50454 41475 51454 41504
rect 37896 41239 38556 41252
rect 43695 41251 44325 41344
rect 50454 41326 51454 41355
rect 50454 41280 50467 41326
rect 50513 41280 50571 41326
rect 50617 41280 50674 41326
rect 50720 41280 50777 41326
rect 50823 41280 50880 41326
rect 50926 41280 50983 41326
rect 51029 41280 51086 41326
rect 51132 41280 51189 41326
rect 51235 41280 51292 41326
rect 51338 41280 51395 41326
rect 51441 41280 51454 41326
rect 37896 41193 37909 41239
rect 37955 41193 38026 41239
rect 38072 41193 38143 41239
rect 38189 41193 38261 41239
rect 38307 41193 38379 41239
rect 38425 41193 38497 41239
rect 38543 41193 38556 41239
rect 37896 41164 38556 41193
rect 33671 41102 34671 41131
rect 33671 41056 33684 41102
rect 33730 41056 33787 41102
rect 33833 41056 33890 41102
rect 33936 41056 33993 41102
rect 34039 41056 34096 41102
rect 34142 41056 34199 41102
rect 34245 41056 34302 41102
rect 34348 41056 34405 41102
rect 34451 41056 34508 41102
rect 34554 41056 34612 41102
rect 34658 41056 34671 41102
rect 33671 40995 34671 41056
rect 33671 40843 34671 40875
rect 33671 40797 33816 40843
rect 33862 40797 34002 40843
rect 34048 40797 34189 40843
rect 34235 40797 34376 40843
rect 34422 40797 34562 40843
rect 34608 40797 34671 40843
rect 50454 41251 51454 41280
rect 37896 41015 38556 41044
rect 37896 40969 37909 41015
rect 37955 40969 38026 41015
rect 38072 40969 38143 41015
rect 38189 40969 38261 41015
rect 38307 40969 38379 41015
rect 38425 40969 38497 41015
rect 38543 40969 38556 41015
rect 37896 40940 38556 40969
rect 39598 41015 39730 41028
rect 43695 41027 44325 41131
rect 39598 40969 39641 41015
rect 39687 40969 39730 41015
rect 39598 40940 39730 40969
rect 50454 41102 51454 41131
rect 50454 41056 50467 41102
rect 50513 41056 50571 41102
rect 50617 41056 50674 41102
rect 50720 41056 50777 41102
rect 50823 41056 50880 41102
rect 50926 41056 50983 41102
rect 51029 41056 51086 41102
rect 51132 41056 51189 41102
rect 51235 41056 51292 41102
rect 51338 41056 51395 41102
rect 51441 41056 51454 41102
rect 50454 40995 51454 41056
rect 43695 40857 44325 40907
rect 33671 40751 34671 40797
rect 37896 40791 38556 40820
rect 37896 40745 37909 40791
rect 37955 40745 38026 40791
rect 38072 40745 38143 40791
rect 38189 40745 38261 40791
rect 38307 40745 38379 40791
rect 38425 40745 38497 40791
rect 38543 40745 38556 40791
rect 37896 40732 38556 40745
rect 39598 40791 39730 40820
rect 39598 40745 39641 40791
rect 39687 40745 39730 40791
rect 43695 40811 43739 40857
rect 43785 40811 43906 40857
rect 43952 40811 44071 40857
rect 44117 40811 44236 40857
rect 44282 40811 44325 40857
rect 50454 40843 51454 40875
rect 43695 40764 44325 40811
rect 39598 40732 39730 40745
rect 50454 40797 50516 40843
rect 50562 40797 50703 40843
rect 50749 40797 50890 40843
rect 50936 40797 51076 40843
rect 51122 40797 51263 40843
rect 51309 40797 51454 40843
rect 50454 40751 51454 40797
rect 33671 40457 34671 40503
rect 33671 40411 33816 40457
rect 33862 40411 34002 40457
rect 34048 40411 34189 40457
rect 34235 40411 34376 40457
rect 34422 40411 34562 40457
rect 34608 40411 34671 40457
rect 37896 40509 38556 40522
rect 37896 40463 37909 40509
rect 37955 40463 38026 40509
rect 38072 40463 38143 40509
rect 38189 40463 38261 40509
rect 38307 40463 38379 40509
rect 38425 40463 38497 40509
rect 38543 40463 38556 40509
rect 37896 40434 38556 40463
rect 39598 40509 39730 40522
rect 39598 40463 39641 40509
rect 39687 40463 39730 40509
rect 39598 40434 39730 40463
rect 43695 40443 44325 40490
rect 33671 40379 34671 40411
rect 33671 40198 34671 40259
rect 33671 40152 33684 40198
rect 33730 40152 33787 40198
rect 33833 40152 33890 40198
rect 33936 40152 33993 40198
rect 34039 40152 34096 40198
rect 34142 40152 34199 40198
rect 34245 40152 34302 40198
rect 34348 40152 34405 40198
rect 34451 40152 34508 40198
rect 34554 40152 34612 40198
rect 34658 40152 34671 40198
rect 33671 40123 34671 40152
rect 37896 40285 38556 40314
rect 37896 40239 37909 40285
rect 37955 40239 38026 40285
rect 38072 40239 38143 40285
rect 38189 40239 38261 40285
rect 38307 40239 38379 40285
rect 38425 40239 38497 40285
rect 38543 40239 38556 40285
rect 37896 40210 38556 40239
rect 43695 40397 43739 40443
rect 43785 40397 43906 40443
rect 43952 40397 44071 40443
rect 44117 40397 44236 40443
rect 44282 40397 44325 40443
rect 43695 40347 44325 40397
rect 50454 40457 51454 40503
rect 39598 40285 39730 40314
rect 39598 40239 39641 40285
rect 39687 40239 39730 40285
rect 39598 40226 39730 40239
rect 50454 40411 50516 40457
rect 50562 40411 50703 40457
rect 50749 40411 50890 40457
rect 50936 40411 51076 40457
rect 51122 40411 51263 40457
rect 51309 40411 51454 40457
rect 50454 40379 51454 40411
rect 43695 40123 44325 40227
rect 33671 39974 34671 40003
rect 37896 40061 38556 40090
rect 37896 40015 37909 40061
rect 37955 40015 38026 40061
rect 38072 40015 38143 40061
rect 38189 40015 38261 40061
rect 38307 40015 38379 40061
rect 38425 40015 38497 40061
rect 38543 40015 38556 40061
rect 37896 40002 38556 40015
rect 50454 40198 51454 40259
rect 50454 40152 50467 40198
rect 50513 40152 50571 40198
rect 50617 40152 50674 40198
rect 50720 40152 50777 40198
rect 50823 40152 50880 40198
rect 50926 40152 50983 40198
rect 51029 40152 51086 40198
rect 51132 40152 51189 40198
rect 51235 40152 51292 40198
rect 51338 40152 51395 40198
rect 51441 40152 51454 40198
rect 50454 40123 51454 40152
rect 33671 39928 33684 39974
rect 33730 39928 33787 39974
rect 33833 39928 33890 39974
rect 33936 39928 33993 39974
rect 34039 39928 34096 39974
rect 34142 39928 34199 39974
rect 34245 39928 34302 39974
rect 34348 39928 34405 39974
rect 34451 39928 34508 39974
rect 34554 39928 34612 39974
rect 34658 39928 34671 39974
rect 33671 39899 34671 39928
rect 39727 39974 40167 39987
rect 39727 39928 39740 39974
rect 39786 39928 39862 39974
rect 39908 39928 39985 39974
rect 40031 39928 40108 39974
rect 40154 39928 40167 39974
rect 39727 39899 40167 39928
rect 43695 39910 44325 40003
rect 50454 39974 51454 40003
rect 33671 39750 34671 39779
rect 33671 39704 33684 39750
rect 33730 39704 33787 39750
rect 33833 39704 33890 39750
rect 33936 39704 33993 39750
rect 34039 39704 34096 39750
rect 34142 39704 34199 39750
rect 34245 39704 34302 39750
rect 34348 39704 34405 39750
rect 34451 39704 34508 39750
rect 34554 39704 34612 39750
rect 34658 39704 34671 39750
rect 33671 39675 34671 39704
rect 39727 39750 40167 39779
rect 39727 39704 39740 39750
rect 39786 39704 39862 39750
rect 39908 39704 39985 39750
rect 40031 39704 40108 39750
rect 40154 39704 40167 39750
rect 39727 39675 40167 39704
rect 43695 39750 44325 39790
rect 50454 39928 50467 39974
rect 50513 39928 50571 39974
rect 50617 39928 50674 39974
rect 50720 39928 50777 39974
rect 50823 39928 50880 39974
rect 50926 39928 50983 39974
rect 51029 39928 51086 39974
rect 51132 39928 51189 39974
rect 51235 39928 51292 39974
rect 51338 39928 51395 39974
rect 51441 39928 51454 39974
rect 50454 39899 51454 39928
rect 43695 39704 43739 39750
rect 43785 39704 43906 39750
rect 43952 39704 44071 39750
rect 44117 39704 44236 39750
rect 44282 39704 44325 39750
rect 43695 39664 44325 39704
rect 33671 39526 34671 39555
rect 33671 39480 33684 39526
rect 33730 39480 33787 39526
rect 33833 39480 33890 39526
rect 33936 39480 33993 39526
rect 34039 39480 34096 39526
rect 34142 39480 34199 39526
rect 34245 39480 34302 39526
rect 34348 39480 34405 39526
rect 34451 39480 34508 39526
rect 34554 39480 34612 39526
rect 34658 39480 34671 39526
rect 33671 39451 34671 39480
rect 39727 39526 40167 39555
rect 39727 39480 39740 39526
rect 39786 39480 39862 39526
rect 39908 39480 39985 39526
rect 40031 39480 40108 39526
rect 40154 39480 40167 39526
rect 39727 39467 40167 39480
rect 50454 39750 51454 39779
rect 50454 39704 50467 39750
rect 50513 39704 50571 39750
rect 50617 39704 50674 39750
rect 50720 39704 50777 39750
rect 50823 39704 50880 39750
rect 50926 39704 50983 39750
rect 51029 39704 51086 39750
rect 51132 39704 51189 39750
rect 51235 39704 51292 39750
rect 51338 39704 51395 39750
rect 51441 39704 51454 39750
rect 50454 39675 51454 39704
rect 37896 39439 38556 39452
rect 43695 39451 44325 39544
rect 50454 39526 51454 39555
rect 50454 39480 50467 39526
rect 50513 39480 50571 39526
rect 50617 39480 50674 39526
rect 50720 39480 50777 39526
rect 50823 39480 50880 39526
rect 50926 39480 50983 39526
rect 51029 39480 51086 39526
rect 51132 39480 51189 39526
rect 51235 39480 51292 39526
rect 51338 39480 51395 39526
rect 51441 39480 51454 39526
rect 37896 39393 37909 39439
rect 37955 39393 38026 39439
rect 38072 39393 38143 39439
rect 38189 39393 38261 39439
rect 38307 39393 38379 39439
rect 38425 39393 38497 39439
rect 38543 39393 38556 39439
rect 37896 39364 38556 39393
rect 33671 39302 34671 39331
rect 33671 39256 33684 39302
rect 33730 39256 33787 39302
rect 33833 39256 33890 39302
rect 33936 39256 33993 39302
rect 34039 39256 34096 39302
rect 34142 39256 34199 39302
rect 34245 39256 34302 39302
rect 34348 39256 34405 39302
rect 34451 39256 34508 39302
rect 34554 39256 34612 39302
rect 34658 39256 34671 39302
rect 33671 39195 34671 39256
rect 33671 39043 34671 39075
rect 33671 38997 33816 39043
rect 33862 38997 34002 39043
rect 34048 38997 34189 39043
rect 34235 38997 34376 39043
rect 34422 38997 34562 39043
rect 34608 38997 34671 39043
rect 50454 39451 51454 39480
rect 37896 39215 38556 39244
rect 37896 39169 37909 39215
rect 37955 39169 38026 39215
rect 38072 39169 38143 39215
rect 38189 39169 38261 39215
rect 38307 39169 38379 39215
rect 38425 39169 38497 39215
rect 38543 39169 38556 39215
rect 37896 39140 38556 39169
rect 39598 39215 39730 39228
rect 43695 39227 44325 39331
rect 39598 39169 39641 39215
rect 39687 39169 39730 39215
rect 39598 39140 39730 39169
rect 50454 39302 51454 39331
rect 50454 39256 50467 39302
rect 50513 39256 50571 39302
rect 50617 39256 50674 39302
rect 50720 39256 50777 39302
rect 50823 39256 50880 39302
rect 50926 39256 50983 39302
rect 51029 39256 51086 39302
rect 51132 39256 51189 39302
rect 51235 39256 51292 39302
rect 51338 39256 51395 39302
rect 51441 39256 51454 39302
rect 50454 39195 51454 39256
rect 43695 39057 44325 39107
rect 33671 38951 34671 38997
rect 37896 38991 38556 39020
rect 37896 38945 37909 38991
rect 37955 38945 38026 38991
rect 38072 38945 38143 38991
rect 38189 38945 38261 38991
rect 38307 38945 38379 38991
rect 38425 38945 38497 38991
rect 38543 38945 38556 38991
rect 37896 38932 38556 38945
rect 39598 38991 39730 39020
rect 39598 38945 39641 38991
rect 39687 38945 39730 38991
rect 43695 39011 43739 39057
rect 43785 39011 43906 39057
rect 43952 39011 44071 39057
rect 44117 39011 44236 39057
rect 44282 39011 44325 39057
rect 50454 39043 51454 39075
rect 43695 38964 44325 39011
rect 39598 38932 39730 38945
rect 50454 38997 50516 39043
rect 50562 38997 50703 39043
rect 50749 38997 50890 39043
rect 50936 38997 51076 39043
rect 51122 38997 51263 39043
rect 51309 38997 51454 39043
rect 50454 38951 51454 38997
rect 33671 38657 34671 38703
rect 33671 38611 33816 38657
rect 33862 38611 34002 38657
rect 34048 38611 34189 38657
rect 34235 38611 34376 38657
rect 34422 38611 34562 38657
rect 34608 38611 34671 38657
rect 37896 38709 38556 38722
rect 37896 38663 37909 38709
rect 37955 38663 38026 38709
rect 38072 38663 38143 38709
rect 38189 38663 38261 38709
rect 38307 38663 38379 38709
rect 38425 38663 38497 38709
rect 38543 38663 38556 38709
rect 37896 38634 38556 38663
rect 39598 38709 39730 38722
rect 39598 38663 39641 38709
rect 39687 38663 39730 38709
rect 39598 38634 39730 38663
rect 43695 38643 44325 38690
rect 33671 38579 34671 38611
rect 33671 38398 34671 38459
rect 33671 38352 33684 38398
rect 33730 38352 33787 38398
rect 33833 38352 33890 38398
rect 33936 38352 33993 38398
rect 34039 38352 34096 38398
rect 34142 38352 34199 38398
rect 34245 38352 34302 38398
rect 34348 38352 34405 38398
rect 34451 38352 34508 38398
rect 34554 38352 34612 38398
rect 34658 38352 34671 38398
rect 33671 38323 34671 38352
rect 37896 38485 38556 38514
rect 37896 38439 37909 38485
rect 37955 38439 38026 38485
rect 38072 38439 38143 38485
rect 38189 38439 38261 38485
rect 38307 38439 38379 38485
rect 38425 38439 38497 38485
rect 38543 38439 38556 38485
rect 37896 38410 38556 38439
rect 43695 38597 43739 38643
rect 43785 38597 43906 38643
rect 43952 38597 44071 38643
rect 44117 38597 44236 38643
rect 44282 38597 44325 38643
rect 43695 38547 44325 38597
rect 50454 38657 51454 38703
rect 39598 38485 39730 38514
rect 39598 38439 39641 38485
rect 39687 38439 39730 38485
rect 39598 38426 39730 38439
rect 50454 38611 50516 38657
rect 50562 38611 50703 38657
rect 50749 38611 50890 38657
rect 50936 38611 51076 38657
rect 51122 38611 51263 38657
rect 51309 38611 51454 38657
rect 50454 38579 51454 38611
rect 43695 38323 44325 38427
rect 33671 38174 34671 38203
rect 37896 38261 38556 38290
rect 37896 38215 37909 38261
rect 37955 38215 38026 38261
rect 38072 38215 38143 38261
rect 38189 38215 38261 38261
rect 38307 38215 38379 38261
rect 38425 38215 38497 38261
rect 38543 38215 38556 38261
rect 37896 38202 38556 38215
rect 50454 38398 51454 38459
rect 50454 38352 50467 38398
rect 50513 38352 50571 38398
rect 50617 38352 50674 38398
rect 50720 38352 50777 38398
rect 50823 38352 50880 38398
rect 50926 38352 50983 38398
rect 51029 38352 51086 38398
rect 51132 38352 51189 38398
rect 51235 38352 51292 38398
rect 51338 38352 51395 38398
rect 51441 38352 51454 38398
rect 50454 38323 51454 38352
rect 33671 38128 33684 38174
rect 33730 38128 33787 38174
rect 33833 38128 33890 38174
rect 33936 38128 33993 38174
rect 34039 38128 34096 38174
rect 34142 38128 34199 38174
rect 34245 38128 34302 38174
rect 34348 38128 34405 38174
rect 34451 38128 34508 38174
rect 34554 38128 34612 38174
rect 34658 38128 34671 38174
rect 33671 38099 34671 38128
rect 39727 38174 40167 38187
rect 39727 38128 39740 38174
rect 39786 38128 39862 38174
rect 39908 38128 39985 38174
rect 40031 38128 40108 38174
rect 40154 38128 40167 38174
rect 39727 38099 40167 38128
rect 43695 38110 44325 38203
rect 50454 38174 51454 38203
rect 33671 37950 34671 37979
rect 33671 37904 33684 37950
rect 33730 37904 33787 37950
rect 33833 37904 33890 37950
rect 33936 37904 33993 37950
rect 34039 37904 34096 37950
rect 34142 37904 34199 37950
rect 34245 37904 34302 37950
rect 34348 37904 34405 37950
rect 34451 37904 34508 37950
rect 34554 37904 34612 37950
rect 34658 37904 34671 37950
rect 33671 37875 34671 37904
rect 39727 37950 40167 37979
rect 39727 37904 39740 37950
rect 39786 37904 39862 37950
rect 39908 37904 39985 37950
rect 40031 37904 40108 37950
rect 40154 37904 40167 37950
rect 39727 37875 40167 37904
rect 43695 37950 44325 37990
rect 50454 38128 50467 38174
rect 50513 38128 50571 38174
rect 50617 38128 50674 38174
rect 50720 38128 50777 38174
rect 50823 38128 50880 38174
rect 50926 38128 50983 38174
rect 51029 38128 51086 38174
rect 51132 38128 51189 38174
rect 51235 38128 51292 38174
rect 51338 38128 51395 38174
rect 51441 38128 51454 38174
rect 50454 38099 51454 38128
rect 43695 37904 43739 37950
rect 43785 37904 43906 37950
rect 43952 37904 44071 37950
rect 44117 37904 44236 37950
rect 44282 37904 44325 37950
rect 43695 37864 44325 37904
rect 33671 37726 34671 37755
rect 33671 37680 33684 37726
rect 33730 37680 33787 37726
rect 33833 37680 33890 37726
rect 33936 37680 33993 37726
rect 34039 37680 34096 37726
rect 34142 37680 34199 37726
rect 34245 37680 34302 37726
rect 34348 37680 34405 37726
rect 34451 37680 34508 37726
rect 34554 37680 34612 37726
rect 34658 37680 34671 37726
rect 33671 37651 34671 37680
rect 39727 37726 40167 37755
rect 39727 37680 39740 37726
rect 39786 37680 39862 37726
rect 39908 37680 39985 37726
rect 40031 37680 40108 37726
rect 40154 37680 40167 37726
rect 39727 37667 40167 37680
rect 50454 37950 51454 37979
rect 50454 37904 50467 37950
rect 50513 37904 50571 37950
rect 50617 37904 50674 37950
rect 50720 37904 50777 37950
rect 50823 37904 50880 37950
rect 50926 37904 50983 37950
rect 51029 37904 51086 37950
rect 51132 37904 51189 37950
rect 51235 37904 51292 37950
rect 51338 37904 51395 37950
rect 51441 37904 51454 37950
rect 50454 37875 51454 37904
rect 37896 37639 38556 37652
rect 43695 37651 44325 37744
rect 50454 37726 51454 37755
rect 50454 37680 50467 37726
rect 50513 37680 50571 37726
rect 50617 37680 50674 37726
rect 50720 37680 50777 37726
rect 50823 37680 50880 37726
rect 50926 37680 50983 37726
rect 51029 37680 51086 37726
rect 51132 37680 51189 37726
rect 51235 37680 51292 37726
rect 51338 37680 51395 37726
rect 51441 37680 51454 37726
rect 37896 37593 37909 37639
rect 37955 37593 38026 37639
rect 38072 37593 38143 37639
rect 38189 37593 38261 37639
rect 38307 37593 38379 37639
rect 38425 37593 38497 37639
rect 38543 37593 38556 37639
rect 37896 37564 38556 37593
rect 33671 37502 34671 37531
rect 33671 37456 33684 37502
rect 33730 37456 33787 37502
rect 33833 37456 33890 37502
rect 33936 37456 33993 37502
rect 34039 37456 34096 37502
rect 34142 37456 34199 37502
rect 34245 37456 34302 37502
rect 34348 37456 34405 37502
rect 34451 37456 34508 37502
rect 34554 37456 34612 37502
rect 34658 37456 34671 37502
rect 33671 37395 34671 37456
rect 33671 37243 34671 37275
rect 33671 37197 33816 37243
rect 33862 37197 34002 37243
rect 34048 37197 34189 37243
rect 34235 37197 34376 37243
rect 34422 37197 34562 37243
rect 34608 37197 34671 37243
rect 50454 37651 51454 37680
rect 37896 37415 38556 37444
rect 37896 37369 37909 37415
rect 37955 37369 38026 37415
rect 38072 37369 38143 37415
rect 38189 37369 38261 37415
rect 38307 37369 38379 37415
rect 38425 37369 38497 37415
rect 38543 37369 38556 37415
rect 37896 37340 38556 37369
rect 39598 37415 39730 37428
rect 43695 37427 44325 37531
rect 39598 37369 39641 37415
rect 39687 37369 39730 37415
rect 39598 37340 39730 37369
rect 50454 37502 51454 37531
rect 50454 37456 50467 37502
rect 50513 37456 50571 37502
rect 50617 37456 50674 37502
rect 50720 37456 50777 37502
rect 50823 37456 50880 37502
rect 50926 37456 50983 37502
rect 51029 37456 51086 37502
rect 51132 37456 51189 37502
rect 51235 37456 51292 37502
rect 51338 37456 51395 37502
rect 51441 37456 51454 37502
rect 50454 37395 51454 37456
rect 43695 37257 44325 37307
rect 33671 37151 34671 37197
rect 37896 37191 38556 37220
rect 37896 37145 37909 37191
rect 37955 37145 38026 37191
rect 38072 37145 38143 37191
rect 38189 37145 38261 37191
rect 38307 37145 38379 37191
rect 38425 37145 38497 37191
rect 38543 37145 38556 37191
rect 37896 37132 38556 37145
rect 39598 37191 39730 37220
rect 39598 37145 39641 37191
rect 39687 37145 39730 37191
rect 43695 37211 43739 37257
rect 43785 37211 43906 37257
rect 43952 37211 44071 37257
rect 44117 37211 44236 37257
rect 44282 37211 44325 37257
rect 50454 37243 51454 37275
rect 43695 37164 44325 37211
rect 39598 37132 39730 37145
rect 50454 37197 50516 37243
rect 50562 37197 50703 37243
rect 50749 37197 50890 37243
rect 50936 37197 51076 37243
rect 51122 37197 51263 37243
rect 51309 37197 51454 37243
rect 50454 37151 51454 37197
rect 33671 36857 34671 36903
rect 33671 36811 33816 36857
rect 33862 36811 34002 36857
rect 34048 36811 34189 36857
rect 34235 36811 34376 36857
rect 34422 36811 34562 36857
rect 34608 36811 34671 36857
rect 37896 36909 38556 36922
rect 37896 36863 37909 36909
rect 37955 36863 38026 36909
rect 38072 36863 38143 36909
rect 38189 36863 38261 36909
rect 38307 36863 38379 36909
rect 38425 36863 38497 36909
rect 38543 36863 38556 36909
rect 37896 36834 38556 36863
rect 39598 36909 39730 36922
rect 39598 36863 39641 36909
rect 39687 36863 39730 36909
rect 39598 36834 39730 36863
rect 43695 36843 44325 36890
rect 33671 36779 34671 36811
rect 33671 36598 34671 36659
rect 33671 36552 33684 36598
rect 33730 36552 33787 36598
rect 33833 36552 33890 36598
rect 33936 36552 33993 36598
rect 34039 36552 34096 36598
rect 34142 36552 34199 36598
rect 34245 36552 34302 36598
rect 34348 36552 34405 36598
rect 34451 36552 34508 36598
rect 34554 36552 34612 36598
rect 34658 36552 34671 36598
rect 33671 36523 34671 36552
rect 37896 36685 38556 36714
rect 37896 36639 37909 36685
rect 37955 36639 38026 36685
rect 38072 36639 38143 36685
rect 38189 36639 38261 36685
rect 38307 36639 38379 36685
rect 38425 36639 38497 36685
rect 38543 36639 38556 36685
rect 37896 36610 38556 36639
rect 43695 36797 43739 36843
rect 43785 36797 43906 36843
rect 43952 36797 44071 36843
rect 44117 36797 44236 36843
rect 44282 36797 44325 36843
rect 43695 36747 44325 36797
rect 50454 36857 51454 36903
rect 39598 36685 39730 36714
rect 39598 36639 39641 36685
rect 39687 36639 39730 36685
rect 39598 36626 39730 36639
rect 50454 36811 50516 36857
rect 50562 36811 50703 36857
rect 50749 36811 50890 36857
rect 50936 36811 51076 36857
rect 51122 36811 51263 36857
rect 51309 36811 51454 36857
rect 50454 36779 51454 36811
rect 43695 36523 44325 36627
rect 33671 36374 34671 36403
rect 37896 36461 38556 36490
rect 37896 36415 37909 36461
rect 37955 36415 38026 36461
rect 38072 36415 38143 36461
rect 38189 36415 38261 36461
rect 38307 36415 38379 36461
rect 38425 36415 38497 36461
rect 38543 36415 38556 36461
rect 37896 36402 38556 36415
rect 50454 36598 51454 36659
rect 50454 36552 50467 36598
rect 50513 36552 50571 36598
rect 50617 36552 50674 36598
rect 50720 36552 50777 36598
rect 50823 36552 50880 36598
rect 50926 36552 50983 36598
rect 51029 36552 51086 36598
rect 51132 36552 51189 36598
rect 51235 36552 51292 36598
rect 51338 36552 51395 36598
rect 51441 36552 51454 36598
rect 50454 36523 51454 36552
rect 33671 36328 33684 36374
rect 33730 36328 33787 36374
rect 33833 36328 33890 36374
rect 33936 36328 33993 36374
rect 34039 36328 34096 36374
rect 34142 36328 34199 36374
rect 34245 36328 34302 36374
rect 34348 36328 34405 36374
rect 34451 36328 34508 36374
rect 34554 36328 34612 36374
rect 34658 36328 34671 36374
rect 33671 36299 34671 36328
rect 39727 36374 40167 36387
rect 39727 36328 39740 36374
rect 39786 36328 39862 36374
rect 39908 36328 39985 36374
rect 40031 36328 40108 36374
rect 40154 36328 40167 36374
rect 39727 36299 40167 36328
rect 43695 36310 44325 36403
rect 50454 36374 51454 36403
rect 33671 36150 34671 36179
rect 33671 36104 33684 36150
rect 33730 36104 33787 36150
rect 33833 36104 33890 36150
rect 33936 36104 33993 36150
rect 34039 36104 34096 36150
rect 34142 36104 34199 36150
rect 34245 36104 34302 36150
rect 34348 36104 34405 36150
rect 34451 36104 34508 36150
rect 34554 36104 34612 36150
rect 34658 36104 34671 36150
rect 33671 36091 34671 36104
rect 39727 36150 40167 36179
rect 39727 36104 39740 36150
rect 39786 36104 39862 36150
rect 39908 36104 39985 36150
rect 40031 36104 40108 36150
rect 40154 36104 40167 36150
rect 39727 36091 40167 36104
rect 43695 36150 44325 36190
rect 50454 36328 50467 36374
rect 50513 36328 50571 36374
rect 50617 36328 50674 36374
rect 50720 36328 50777 36374
rect 50823 36328 50880 36374
rect 50926 36328 50983 36374
rect 51029 36328 51086 36374
rect 51132 36328 51189 36374
rect 51235 36328 51292 36374
rect 51338 36328 51395 36374
rect 51441 36328 51454 36374
rect 50454 36299 51454 36328
rect 43695 36104 43739 36150
rect 43785 36104 43906 36150
rect 43952 36104 44071 36150
rect 44117 36104 44236 36150
rect 44282 36104 44325 36150
rect 43695 36058 44325 36104
rect 50454 36150 51454 36179
rect 50454 36104 50467 36150
rect 50513 36104 50571 36150
rect 50617 36104 50674 36150
rect 50720 36104 50777 36150
rect 50823 36104 50880 36150
rect 50926 36104 50983 36150
rect 51029 36104 51086 36150
rect 51132 36104 51189 36150
rect 51235 36104 51292 36150
rect 51338 36104 51395 36150
rect 51441 36104 51454 36150
rect 50454 36091 51454 36104
<< mvpdiff >>
rect 29274 65850 30373 65896
rect 29274 65804 29317 65850
rect 29363 65804 29478 65850
rect 29524 65804 29638 65850
rect 29684 65804 29798 65850
rect 29844 65804 29959 65850
rect 30005 65804 30121 65850
rect 30167 65804 30284 65850
rect 30330 65804 30373 65850
rect 29274 65771 30373 65804
rect 35396 65818 37922 65831
rect 35396 65772 35409 65818
rect 37291 65772 37348 65818
rect 37394 65772 37451 65818
rect 37497 65772 37554 65818
rect 37600 65772 37657 65818
rect 37703 65772 37760 65818
rect 37806 65772 37863 65818
rect 37909 65772 37922 65818
rect 35396 65743 37922 65772
rect 35396 65594 37922 65623
rect 35396 65548 35409 65594
rect 37291 65548 37348 65594
rect 37394 65548 37451 65594
rect 37497 65548 37554 65594
rect 37600 65548 37657 65594
rect 37703 65548 37760 65594
rect 37806 65548 37863 65594
rect 37909 65548 37922 65594
rect 35396 65519 37922 65548
rect 38363 65594 39681 65607
rect 38363 65548 38376 65594
rect 38422 65548 38479 65594
rect 38525 65548 38582 65594
rect 38628 65548 38686 65594
rect 38732 65548 38790 65594
rect 38836 65548 38894 65594
rect 38940 65548 38998 65594
rect 39044 65548 39102 65594
rect 39148 65548 39206 65594
rect 39252 65548 39310 65594
rect 39356 65548 39414 65594
rect 39460 65548 39518 65594
rect 39564 65548 39622 65594
rect 39668 65548 39681 65594
rect 38363 65519 39681 65548
rect 42663 65594 43981 65607
rect 42663 65548 42676 65594
rect 42722 65548 42779 65594
rect 42825 65548 42882 65594
rect 42928 65548 42986 65594
rect 43032 65548 43090 65594
rect 43136 65548 43194 65594
rect 43240 65548 43298 65594
rect 43344 65548 43402 65594
rect 43448 65548 43506 65594
rect 43552 65548 43610 65594
rect 43656 65548 43714 65594
rect 43760 65548 43818 65594
rect 43864 65548 43922 65594
rect 43968 65548 43981 65594
rect 42663 65519 43981 65548
rect 47101 65818 49627 65831
rect 47101 65772 47114 65818
rect 48996 65772 49053 65818
rect 49099 65772 49156 65818
rect 49202 65772 49259 65818
rect 49305 65772 49362 65818
rect 49408 65772 49465 65818
rect 49511 65772 49568 65818
rect 49614 65772 49627 65818
rect 47101 65743 49627 65772
rect 35396 65370 37922 65399
rect 35396 65324 35409 65370
rect 37291 65324 37348 65370
rect 37394 65324 37451 65370
rect 37497 65324 37554 65370
rect 37600 65324 37657 65370
rect 37703 65324 37760 65370
rect 37806 65324 37863 65370
rect 37909 65324 37922 65370
rect 35396 65311 37922 65324
rect 38363 65370 39681 65399
rect 38363 65324 38376 65370
rect 38422 65324 38479 65370
rect 38525 65324 38582 65370
rect 38628 65324 38686 65370
rect 38732 65324 38790 65370
rect 38836 65324 38894 65370
rect 38940 65324 38998 65370
rect 39044 65324 39102 65370
rect 39148 65324 39206 65370
rect 39252 65324 39310 65370
rect 39356 65324 39414 65370
rect 39460 65324 39518 65370
rect 39564 65324 39622 65370
rect 39668 65324 39681 65370
rect 38363 65311 39681 65324
rect 45333 65594 46651 65607
rect 45333 65548 45346 65594
rect 45392 65548 45449 65594
rect 45495 65548 45552 65594
rect 45598 65548 45656 65594
rect 45702 65548 45760 65594
rect 45806 65548 45864 65594
rect 45910 65548 45968 65594
rect 46014 65548 46072 65594
rect 46118 65548 46176 65594
rect 46222 65548 46280 65594
rect 46326 65548 46384 65594
rect 46430 65548 46488 65594
rect 46534 65548 46592 65594
rect 46638 65548 46651 65594
rect 45333 65519 46651 65548
rect 47101 65594 49627 65623
rect 47101 65548 47114 65594
rect 48996 65548 49053 65594
rect 49099 65548 49156 65594
rect 49202 65548 49259 65594
rect 49305 65548 49362 65594
rect 49408 65548 49465 65594
rect 49511 65548 49568 65594
rect 49614 65548 49627 65594
rect 47101 65519 49627 65548
rect 54750 65850 55849 65896
rect 54750 65804 54793 65850
rect 54839 65804 54956 65850
rect 55002 65804 55118 65850
rect 55164 65804 55279 65850
rect 55325 65804 55439 65850
rect 55485 65804 55599 65850
rect 55645 65804 55760 65850
rect 55806 65804 55849 65850
rect 54750 65771 55849 65804
rect 42663 65370 43981 65399
rect 42663 65324 42676 65370
rect 42722 65324 42779 65370
rect 42825 65324 42882 65370
rect 42928 65324 42986 65370
rect 43032 65324 43090 65370
rect 43136 65324 43194 65370
rect 43240 65324 43298 65370
rect 43344 65324 43402 65370
rect 43448 65324 43506 65370
rect 43552 65324 43610 65370
rect 43656 65324 43714 65370
rect 43760 65324 43818 65370
rect 43864 65324 43922 65370
rect 43968 65324 43981 65370
rect 42663 65311 43981 65324
rect 45333 65370 46651 65399
rect 45333 65324 45346 65370
rect 45392 65324 45449 65370
rect 45495 65324 45552 65370
rect 45598 65324 45656 65370
rect 45702 65324 45760 65370
rect 45806 65324 45864 65370
rect 45910 65324 45968 65370
rect 46014 65324 46072 65370
rect 46118 65324 46176 65370
rect 46222 65324 46280 65370
rect 46326 65324 46384 65370
rect 46430 65324 46488 65370
rect 46534 65324 46592 65370
rect 46638 65324 46651 65370
rect 45333 65311 46651 65324
rect 47101 65370 49627 65399
rect 47101 65324 47114 65370
rect 48996 65324 49053 65370
rect 49099 65324 49156 65370
rect 49202 65324 49259 65370
rect 49305 65324 49362 65370
rect 49408 65324 49465 65370
rect 49511 65324 49568 65370
rect 49614 65324 49627 65370
rect 47101 65311 49627 65324
rect 29274 64950 30373 64983
rect 29274 64904 29317 64950
rect 29363 64904 29478 64950
rect 29524 64904 29638 64950
rect 29684 64904 29798 64950
rect 29844 64904 29959 64950
rect 30005 64904 30121 64950
rect 30167 64904 30284 64950
rect 30330 64904 30373 64950
rect 29274 64871 30373 64904
rect 31336 64950 33336 64963
rect 31336 64904 31349 64950
rect 33323 64904 33336 64950
rect 31336 64875 33336 64904
rect 31336 64726 33336 64755
rect 31336 64680 31349 64726
rect 33323 64680 33336 64726
rect 31336 64651 33336 64680
rect 31336 64502 33336 64531
rect 31336 64456 31349 64502
rect 33323 64456 33336 64502
rect 31336 64427 33336 64456
rect 44799 64950 45323 64963
rect 44799 64904 44812 64950
rect 44858 64904 44925 64950
rect 44971 64904 45038 64950
rect 45084 64904 45151 64950
rect 45197 64904 45264 64950
rect 45310 64904 45323 64950
rect 44799 64875 45323 64904
rect 51789 64950 53789 64963
rect 51789 64904 51802 64950
rect 53776 64904 53789 64950
rect 51789 64875 53789 64904
rect 35260 64639 36360 64652
rect 35260 64593 35273 64639
rect 35523 64593 35580 64639
rect 35626 64593 35683 64639
rect 35729 64593 35786 64639
rect 35832 64593 35889 64639
rect 35935 64593 35992 64639
rect 36038 64593 36095 64639
rect 36141 64593 36198 64639
rect 36244 64593 36301 64639
rect 36347 64593 36360 64639
rect 35260 64564 36360 64593
rect 36841 64639 37501 64652
rect 36841 64593 36854 64639
rect 36900 64593 36971 64639
rect 37017 64593 37088 64639
rect 37134 64593 37206 64639
rect 37252 64593 37324 64639
rect 37370 64593 37442 64639
rect 37488 64593 37501 64639
rect 36841 64564 37501 64593
rect 44799 64726 45323 64755
rect 44799 64680 44812 64726
rect 44858 64680 44925 64726
rect 44971 64680 45038 64726
rect 45084 64680 45151 64726
rect 45197 64680 45264 64726
rect 45310 64680 45323 64726
rect 54750 64950 55849 64983
rect 54750 64904 54793 64950
rect 54839 64904 54956 64950
rect 55002 64904 55118 64950
rect 55164 64904 55279 64950
rect 55325 64904 55439 64950
rect 55485 64904 55599 64950
rect 55645 64904 55760 64950
rect 55806 64904 55849 64950
rect 54750 64871 55849 64904
rect 44799 64651 45323 64680
rect 31336 64278 33336 64307
rect 31336 64232 31349 64278
rect 33323 64232 33336 64278
rect 35260 64415 36360 64444
rect 35260 64369 35273 64415
rect 35523 64369 35580 64415
rect 35626 64369 35683 64415
rect 35729 64369 35786 64415
rect 35832 64369 35889 64415
rect 35935 64369 35992 64415
rect 36038 64369 36095 64415
rect 36141 64369 36198 64415
rect 36244 64369 36301 64415
rect 36347 64369 36360 64415
rect 35260 64340 36360 64369
rect 31336 64219 33336 64232
rect 48765 64639 49865 64652
rect 48765 64593 48778 64639
rect 48824 64593 48881 64639
rect 48927 64593 48984 64639
rect 49030 64593 49087 64639
rect 49133 64593 49190 64639
rect 49236 64593 49293 64639
rect 49339 64593 49396 64639
rect 49442 64593 49499 64639
rect 49545 64593 49602 64639
rect 49852 64593 49865 64639
rect 48765 64564 49865 64593
rect 36841 64415 37501 64444
rect 36841 64369 36854 64415
rect 36900 64369 36971 64415
rect 37017 64369 37088 64415
rect 37134 64369 37206 64415
rect 37252 64369 37324 64415
rect 37370 64369 37442 64415
rect 37488 64369 37501 64415
rect 36841 64340 37501 64369
rect 39008 64415 39326 64428
rect 39008 64369 39021 64415
rect 39067 64369 39144 64415
rect 39190 64369 39267 64415
rect 39313 64369 39326 64415
rect 39008 64340 39326 64369
rect 44799 64502 45323 64531
rect 44799 64456 44812 64502
rect 44858 64456 44925 64502
rect 44971 64456 45038 64502
rect 45084 64456 45151 64502
rect 45197 64456 45264 64502
rect 45310 64456 45323 64502
rect 44799 64427 45323 64456
rect 48765 64415 49865 64444
rect 48765 64369 48778 64415
rect 48824 64369 48881 64415
rect 48927 64369 48984 64415
rect 49030 64369 49087 64415
rect 49133 64369 49190 64415
rect 49236 64369 49293 64415
rect 49339 64369 49396 64415
rect 49442 64369 49499 64415
rect 49545 64369 49602 64415
rect 49852 64369 49865 64415
rect 48765 64340 49865 64369
rect 35260 64191 36360 64220
rect 35260 64145 35273 64191
rect 35523 64145 35580 64191
rect 35626 64145 35683 64191
rect 35729 64145 35786 64191
rect 35832 64145 35889 64191
rect 35935 64145 35992 64191
rect 36038 64145 36095 64191
rect 36141 64145 36198 64191
rect 36244 64145 36301 64191
rect 36347 64145 36360 64191
rect 35260 64132 36360 64145
rect 36841 64191 37501 64220
rect 36841 64145 36854 64191
rect 36900 64145 36971 64191
rect 37017 64145 37088 64191
rect 37134 64145 37206 64191
rect 37252 64145 37324 64191
rect 37370 64145 37442 64191
rect 37488 64145 37501 64191
rect 36841 64132 37501 64145
rect 39008 64191 39326 64220
rect 39008 64145 39021 64191
rect 39067 64145 39144 64191
rect 39190 64145 39267 64191
rect 39313 64145 39326 64191
rect 39008 64132 39326 64145
rect 44799 64278 45323 64307
rect 44799 64232 44812 64278
rect 44858 64232 44925 64278
rect 44971 64232 45038 64278
rect 45084 64232 45151 64278
rect 45197 64232 45264 64278
rect 45310 64232 45323 64278
rect 44799 64219 45323 64232
rect 51789 64726 53789 64755
rect 51789 64680 51802 64726
rect 53776 64680 53789 64726
rect 51789 64651 53789 64680
rect 51789 64502 53789 64531
rect 51789 64456 51802 64502
rect 53776 64456 53789 64502
rect 51789 64427 53789 64456
rect 51789 64278 53789 64307
rect 48765 64191 49865 64220
rect 48765 64145 48778 64191
rect 48824 64145 48881 64191
rect 48927 64145 48984 64191
rect 49030 64145 49087 64191
rect 49133 64145 49190 64191
rect 49236 64145 49293 64191
rect 49339 64145 49396 64191
rect 49442 64145 49499 64191
rect 49545 64145 49602 64191
rect 49852 64145 49865 64191
rect 51789 64232 51802 64278
rect 53776 64232 53789 64278
rect 51789 64219 53789 64232
rect 48765 64132 49865 64145
rect 29274 64050 30373 64083
rect 29274 64004 29317 64050
rect 29363 64004 29478 64050
rect 29524 64004 29638 64050
rect 29684 64004 29798 64050
rect 29844 64004 29959 64050
rect 30005 64004 30121 64050
rect 30167 64004 30284 64050
rect 30330 64004 30373 64050
rect 29274 63971 30373 64004
rect 54750 64050 55849 64083
rect 54750 64004 54793 64050
rect 54839 64004 54956 64050
rect 55002 64004 55118 64050
rect 55164 64004 55279 64050
rect 55325 64004 55439 64050
rect 55485 64004 55599 64050
rect 55645 64004 55760 64050
rect 55806 64004 55849 64050
rect 54750 63971 55849 64004
rect 35260 63909 36360 63922
rect 31336 63822 33336 63835
rect 31336 63776 31349 63822
rect 33323 63776 33336 63822
rect 35260 63863 35273 63909
rect 35523 63863 35580 63909
rect 35626 63863 35683 63909
rect 35729 63863 35786 63909
rect 35832 63863 35889 63909
rect 35935 63863 35992 63909
rect 36038 63863 36095 63909
rect 36141 63863 36198 63909
rect 36244 63863 36301 63909
rect 36347 63863 36360 63909
rect 35260 63834 36360 63863
rect 36841 63909 37501 63922
rect 36841 63863 36854 63909
rect 36900 63863 36971 63909
rect 37017 63863 37088 63909
rect 37134 63863 37206 63909
rect 37252 63863 37324 63909
rect 37370 63863 37442 63909
rect 37488 63863 37501 63909
rect 36841 63834 37501 63863
rect 39008 63909 39326 63922
rect 39008 63863 39021 63909
rect 39067 63863 39144 63909
rect 39190 63863 39267 63909
rect 39313 63863 39326 63909
rect 39008 63834 39326 63863
rect 48765 63909 49865 63922
rect 31336 63747 33336 63776
rect 31336 63598 33336 63627
rect 31336 63552 31349 63598
rect 33323 63552 33336 63598
rect 31336 63523 33336 63552
rect 31336 63374 33336 63403
rect 31336 63328 31349 63374
rect 33323 63328 33336 63374
rect 31336 63299 33336 63328
rect 29274 63150 30373 63183
rect 29274 63104 29317 63150
rect 29363 63104 29478 63150
rect 29524 63104 29638 63150
rect 29684 63104 29798 63150
rect 29844 63104 29959 63150
rect 30005 63104 30121 63150
rect 30167 63104 30284 63150
rect 30330 63104 30373 63150
rect 29274 63071 30373 63104
rect 35260 63685 36360 63714
rect 35260 63639 35273 63685
rect 35523 63639 35580 63685
rect 35626 63639 35683 63685
rect 35729 63639 35786 63685
rect 35832 63639 35889 63685
rect 35935 63639 35992 63685
rect 36038 63639 36095 63685
rect 36141 63639 36198 63685
rect 36244 63639 36301 63685
rect 36347 63639 36360 63685
rect 35260 63610 36360 63639
rect 36841 63685 37501 63714
rect 36841 63639 36854 63685
rect 36900 63639 36971 63685
rect 37017 63639 37088 63685
rect 37134 63639 37206 63685
rect 37252 63639 37324 63685
rect 37370 63639 37442 63685
rect 37488 63639 37501 63685
rect 36841 63610 37501 63639
rect 48765 63863 48778 63909
rect 48824 63863 48881 63909
rect 48927 63863 48984 63909
rect 49030 63863 49087 63909
rect 49133 63863 49190 63909
rect 49236 63863 49293 63909
rect 49339 63863 49396 63909
rect 49442 63863 49499 63909
rect 49545 63863 49602 63909
rect 49852 63863 49865 63909
rect 44799 63822 45323 63835
rect 48765 63834 49865 63863
rect 44799 63776 44812 63822
rect 44858 63776 44925 63822
rect 44971 63776 45038 63822
rect 45084 63776 45151 63822
rect 45197 63776 45264 63822
rect 45310 63776 45323 63822
rect 44799 63747 45323 63776
rect 39008 63685 39326 63714
rect 39008 63639 39021 63685
rect 39067 63639 39144 63685
rect 39190 63639 39267 63685
rect 39313 63639 39326 63685
rect 39008 63626 39326 63639
rect 51789 63822 53789 63835
rect 44799 63598 45323 63627
rect 44799 63552 44812 63598
rect 44858 63552 44925 63598
rect 44971 63552 45038 63598
rect 45084 63552 45151 63598
rect 45197 63552 45264 63598
rect 45310 63552 45323 63598
rect 44799 63523 45323 63552
rect 48765 63685 49865 63714
rect 48765 63639 48778 63685
rect 48824 63639 48881 63685
rect 48927 63639 48984 63685
rect 49030 63639 49087 63685
rect 49133 63639 49190 63685
rect 49236 63639 49293 63685
rect 49339 63639 49396 63685
rect 49442 63639 49499 63685
rect 49545 63639 49602 63685
rect 49852 63639 49865 63685
rect 48765 63610 49865 63639
rect 51789 63776 51802 63822
rect 53776 63776 53789 63822
rect 51789 63747 53789 63776
rect 35260 63461 36360 63490
rect 35260 63415 35273 63461
rect 35523 63415 35580 63461
rect 35626 63415 35683 63461
rect 35729 63415 35786 63461
rect 35832 63415 35889 63461
rect 35935 63415 35992 63461
rect 36038 63415 36095 63461
rect 36141 63415 36198 63461
rect 36244 63415 36301 63461
rect 36347 63415 36360 63461
rect 35260 63402 36360 63415
rect 36841 63461 37501 63490
rect 36841 63415 36854 63461
rect 36900 63415 36971 63461
rect 37017 63415 37088 63461
rect 37134 63415 37206 63461
rect 37252 63415 37324 63461
rect 37370 63415 37442 63461
rect 37488 63415 37501 63461
rect 36841 63402 37501 63415
rect 48765 63461 49865 63490
rect 48765 63415 48778 63461
rect 48824 63415 48881 63461
rect 48927 63415 48984 63461
rect 49030 63415 49087 63461
rect 49133 63415 49190 63461
rect 49236 63415 49293 63461
rect 49339 63415 49396 63461
rect 49442 63415 49499 63461
rect 49545 63415 49602 63461
rect 49852 63415 49865 63461
rect 44799 63374 45323 63403
rect 48765 63402 49865 63415
rect 44799 63328 44812 63374
rect 44858 63328 44925 63374
rect 44971 63328 45038 63374
rect 45084 63328 45151 63374
rect 45197 63328 45264 63374
rect 45310 63328 45323 63374
rect 31336 63150 33336 63179
rect 31336 63104 31349 63150
rect 33323 63104 33336 63150
rect 31336 63075 33336 63104
rect 31336 62926 33336 62955
rect 31336 62880 31349 62926
rect 33323 62880 33336 62926
rect 31336 62851 33336 62880
rect 31336 62702 33336 62731
rect 31336 62656 31349 62702
rect 33323 62656 33336 62702
rect 31336 62627 33336 62656
rect 44799 63299 45323 63328
rect 51789 63598 53789 63627
rect 51789 63552 51802 63598
rect 53776 63552 53789 63598
rect 51789 63523 53789 63552
rect 51789 63374 53789 63403
rect 51789 63328 51802 63374
rect 53776 63328 53789 63374
rect 51789 63299 53789 63328
rect 44799 63150 45323 63179
rect 44799 63104 44812 63150
rect 44858 63104 44925 63150
rect 44971 63104 45038 63150
rect 45084 63104 45151 63150
rect 45197 63104 45264 63150
rect 45310 63104 45323 63150
rect 44799 63075 45323 63104
rect 51789 63150 53789 63179
rect 51789 63104 51802 63150
rect 53776 63104 53789 63150
rect 51789 63075 53789 63104
rect 35260 62839 36360 62852
rect 35260 62793 35273 62839
rect 35523 62793 35580 62839
rect 35626 62793 35683 62839
rect 35729 62793 35786 62839
rect 35832 62793 35889 62839
rect 35935 62793 35992 62839
rect 36038 62793 36095 62839
rect 36141 62793 36198 62839
rect 36244 62793 36301 62839
rect 36347 62793 36360 62839
rect 35260 62764 36360 62793
rect 36841 62839 37501 62852
rect 36841 62793 36854 62839
rect 36900 62793 36971 62839
rect 37017 62793 37088 62839
rect 37134 62793 37206 62839
rect 37252 62793 37324 62839
rect 37370 62793 37442 62839
rect 37488 62793 37501 62839
rect 36841 62764 37501 62793
rect 44799 62926 45323 62955
rect 44799 62880 44812 62926
rect 44858 62880 44925 62926
rect 44971 62880 45038 62926
rect 45084 62880 45151 62926
rect 45197 62880 45264 62926
rect 45310 62880 45323 62926
rect 54750 63150 55849 63183
rect 54750 63104 54793 63150
rect 54839 63104 54956 63150
rect 55002 63104 55118 63150
rect 55164 63104 55279 63150
rect 55325 63104 55439 63150
rect 55485 63104 55599 63150
rect 55645 63104 55760 63150
rect 55806 63104 55849 63150
rect 54750 63071 55849 63104
rect 44799 62851 45323 62880
rect 31336 62478 33336 62507
rect 31336 62432 31349 62478
rect 33323 62432 33336 62478
rect 35260 62615 36360 62644
rect 35260 62569 35273 62615
rect 35523 62569 35580 62615
rect 35626 62569 35683 62615
rect 35729 62569 35786 62615
rect 35832 62569 35889 62615
rect 35935 62569 35992 62615
rect 36038 62569 36095 62615
rect 36141 62569 36198 62615
rect 36244 62569 36301 62615
rect 36347 62569 36360 62615
rect 35260 62540 36360 62569
rect 31336 62419 33336 62432
rect 48765 62839 49865 62852
rect 48765 62793 48778 62839
rect 48824 62793 48881 62839
rect 48927 62793 48984 62839
rect 49030 62793 49087 62839
rect 49133 62793 49190 62839
rect 49236 62793 49293 62839
rect 49339 62793 49396 62839
rect 49442 62793 49499 62839
rect 49545 62793 49602 62839
rect 49852 62793 49865 62839
rect 48765 62764 49865 62793
rect 36841 62615 37501 62644
rect 36841 62569 36854 62615
rect 36900 62569 36971 62615
rect 37017 62569 37088 62615
rect 37134 62569 37206 62615
rect 37252 62569 37324 62615
rect 37370 62569 37442 62615
rect 37488 62569 37501 62615
rect 36841 62540 37501 62569
rect 39008 62615 39326 62628
rect 39008 62569 39021 62615
rect 39067 62569 39144 62615
rect 39190 62569 39267 62615
rect 39313 62569 39326 62615
rect 39008 62540 39326 62569
rect 44799 62702 45323 62731
rect 44799 62656 44812 62702
rect 44858 62656 44925 62702
rect 44971 62656 45038 62702
rect 45084 62656 45151 62702
rect 45197 62656 45264 62702
rect 45310 62656 45323 62702
rect 44799 62627 45323 62656
rect 48765 62615 49865 62644
rect 48765 62569 48778 62615
rect 48824 62569 48881 62615
rect 48927 62569 48984 62615
rect 49030 62569 49087 62615
rect 49133 62569 49190 62615
rect 49236 62569 49293 62615
rect 49339 62569 49396 62615
rect 49442 62569 49499 62615
rect 49545 62569 49602 62615
rect 49852 62569 49865 62615
rect 48765 62540 49865 62569
rect 35260 62391 36360 62420
rect 35260 62345 35273 62391
rect 35523 62345 35580 62391
rect 35626 62345 35683 62391
rect 35729 62345 35786 62391
rect 35832 62345 35889 62391
rect 35935 62345 35992 62391
rect 36038 62345 36095 62391
rect 36141 62345 36198 62391
rect 36244 62345 36301 62391
rect 36347 62345 36360 62391
rect 35260 62332 36360 62345
rect 36841 62391 37501 62420
rect 36841 62345 36854 62391
rect 36900 62345 36971 62391
rect 37017 62345 37088 62391
rect 37134 62345 37206 62391
rect 37252 62345 37324 62391
rect 37370 62345 37442 62391
rect 37488 62345 37501 62391
rect 36841 62332 37501 62345
rect 39008 62391 39326 62420
rect 39008 62345 39021 62391
rect 39067 62345 39144 62391
rect 39190 62345 39267 62391
rect 39313 62345 39326 62391
rect 39008 62332 39326 62345
rect 44799 62478 45323 62507
rect 44799 62432 44812 62478
rect 44858 62432 44925 62478
rect 44971 62432 45038 62478
rect 45084 62432 45151 62478
rect 45197 62432 45264 62478
rect 45310 62432 45323 62478
rect 44799 62419 45323 62432
rect 51789 62926 53789 62955
rect 51789 62880 51802 62926
rect 53776 62880 53789 62926
rect 51789 62851 53789 62880
rect 51789 62702 53789 62731
rect 51789 62656 51802 62702
rect 53776 62656 53789 62702
rect 51789 62627 53789 62656
rect 51789 62478 53789 62507
rect 48765 62391 49865 62420
rect 48765 62345 48778 62391
rect 48824 62345 48881 62391
rect 48927 62345 48984 62391
rect 49030 62345 49087 62391
rect 49133 62345 49190 62391
rect 49236 62345 49293 62391
rect 49339 62345 49396 62391
rect 49442 62345 49499 62391
rect 49545 62345 49602 62391
rect 49852 62345 49865 62391
rect 51789 62432 51802 62478
rect 53776 62432 53789 62478
rect 51789 62419 53789 62432
rect 48765 62332 49865 62345
rect 29274 62250 30373 62283
rect 29274 62204 29317 62250
rect 29363 62204 29478 62250
rect 29524 62204 29638 62250
rect 29684 62204 29798 62250
rect 29844 62204 29959 62250
rect 30005 62204 30121 62250
rect 30167 62204 30284 62250
rect 30330 62204 30373 62250
rect 29274 62171 30373 62204
rect 54750 62250 55849 62283
rect 54750 62204 54793 62250
rect 54839 62204 54956 62250
rect 55002 62204 55118 62250
rect 55164 62204 55279 62250
rect 55325 62204 55439 62250
rect 55485 62204 55599 62250
rect 55645 62204 55760 62250
rect 55806 62204 55849 62250
rect 54750 62171 55849 62204
rect 35260 62109 36360 62122
rect 31336 62022 33336 62035
rect 31336 61976 31349 62022
rect 33323 61976 33336 62022
rect 35260 62063 35273 62109
rect 35523 62063 35580 62109
rect 35626 62063 35683 62109
rect 35729 62063 35786 62109
rect 35832 62063 35889 62109
rect 35935 62063 35992 62109
rect 36038 62063 36095 62109
rect 36141 62063 36198 62109
rect 36244 62063 36301 62109
rect 36347 62063 36360 62109
rect 35260 62034 36360 62063
rect 36841 62109 37501 62122
rect 36841 62063 36854 62109
rect 36900 62063 36971 62109
rect 37017 62063 37088 62109
rect 37134 62063 37206 62109
rect 37252 62063 37324 62109
rect 37370 62063 37442 62109
rect 37488 62063 37501 62109
rect 36841 62034 37501 62063
rect 39008 62109 39326 62122
rect 39008 62063 39021 62109
rect 39067 62063 39144 62109
rect 39190 62063 39267 62109
rect 39313 62063 39326 62109
rect 39008 62034 39326 62063
rect 48765 62109 49865 62122
rect 31336 61947 33336 61976
rect 31336 61798 33336 61827
rect 31336 61752 31349 61798
rect 33323 61752 33336 61798
rect 31336 61723 33336 61752
rect 31336 61574 33336 61603
rect 31336 61528 31349 61574
rect 33323 61528 33336 61574
rect 31336 61499 33336 61528
rect 29274 61350 30373 61383
rect 29274 61304 29317 61350
rect 29363 61304 29478 61350
rect 29524 61304 29638 61350
rect 29684 61304 29798 61350
rect 29844 61304 29959 61350
rect 30005 61304 30121 61350
rect 30167 61304 30284 61350
rect 30330 61304 30373 61350
rect 29274 61271 30373 61304
rect 35260 61885 36360 61914
rect 35260 61839 35273 61885
rect 35523 61839 35580 61885
rect 35626 61839 35683 61885
rect 35729 61839 35786 61885
rect 35832 61839 35889 61885
rect 35935 61839 35992 61885
rect 36038 61839 36095 61885
rect 36141 61839 36198 61885
rect 36244 61839 36301 61885
rect 36347 61839 36360 61885
rect 35260 61810 36360 61839
rect 36841 61885 37501 61914
rect 36841 61839 36854 61885
rect 36900 61839 36971 61885
rect 37017 61839 37088 61885
rect 37134 61839 37206 61885
rect 37252 61839 37324 61885
rect 37370 61839 37442 61885
rect 37488 61839 37501 61885
rect 36841 61810 37501 61839
rect 48765 62063 48778 62109
rect 48824 62063 48881 62109
rect 48927 62063 48984 62109
rect 49030 62063 49087 62109
rect 49133 62063 49190 62109
rect 49236 62063 49293 62109
rect 49339 62063 49396 62109
rect 49442 62063 49499 62109
rect 49545 62063 49602 62109
rect 49852 62063 49865 62109
rect 44799 62022 45323 62035
rect 48765 62034 49865 62063
rect 44799 61976 44812 62022
rect 44858 61976 44925 62022
rect 44971 61976 45038 62022
rect 45084 61976 45151 62022
rect 45197 61976 45264 62022
rect 45310 61976 45323 62022
rect 44799 61947 45323 61976
rect 39008 61885 39326 61914
rect 39008 61839 39021 61885
rect 39067 61839 39144 61885
rect 39190 61839 39267 61885
rect 39313 61839 39326 61885
rect 39008 61826 39326 61839
rect 51789 62022 53789 62035
rect 44799 61798 45323 61827
rect 44799 61752 44812 61798
rect 44858 61752 44925 61798
rect 44971 61752 45038 61798
rect 45084 61752 45151 61798
rect 45197 61752 45264 61798
rect 45310 61752 45323 61798
rect 44799 61723 45323 61752
rect 48765 61885 49865 61914
rect 48765 61839 48778 61885
rect 48824 61839 48881 61885
rect 48927 61839 48984 61885
rect 49030 61839 49087 61885
rect 49133 61839 49190 61885
rect 49236 61839 49293 61885
rect 49339 61839 49396 61885
rect 49442 61839 49499 61885
rect 49545 61839 49602 61885
rect 49852 61839 49865 61885
rect 48765 61810 49865 61839
rect 51789 61976 51802 62022
rect 53776 61976 53789 62022
rect 51789 61947 53789 61976
rect 35260 61661 36360 61690
rect 35260 61615 35273 61661
rect 35523 61615 35580 61661
rect 35626 61615 35683 61661
rect 35729 61615 35786 61661
rect 35832 61615 35889 61661
rect 35935 61615 35992 61661
rect 36038 61615 36095 61661
rect 36141 61615 36198 61661
rect 36244 61615 36301 61661
rect 36347 61615 36360 61661
rect 35260 61602 36360 61615
rect 36841 61661 37501 61690
rect 36841 61615 36854 61661
rect 36900 61615 36971 61661
rect 37017 61615 37088 61661
rect 37134 61615 37206 61661
rect 37252 61615 37324 61661
rect 37370 61615 37442 61661
rect 37488 61615 37501 61661
rect 36841 61602 37501 61615
rect 48765 61661 49865 61690
rect 48765 61615 48778 61661
rect 48824 61615 48881 61661
rect 48927 61615 48984 61661
rect 49030 61615 49087 61661
rect 49133 61615 49190 61661
rect 49236 61615 49293 61661
rect 49339 61615 49396 61661
rect 49442 61615 49499 61661
rect 49545 61615 49602 61661
rect 49852 61615 49865 61661
rect 44799 61574 45323 61603
rect 48765 61602 49865 61615
rect 44799 61528 44812 61574
rect 44858 61528 44925 61574
rect 44971 61528 45038 61574
rect 45084 61528 45151 61574
rect 45197 61528 45264 61574
rect 45310 61528 45323 61574
rect 31336 61350 33336 61379
rect 31336 61304 31349 61350
rect 33323 61304 33336 61350
rect 31336 61275 33336 61304
rect 31336 61126 33336 61155
rect 31336 61080 31349 61126
rect 33323 61080 33336 61126
rect 31336 61051 33336 61080
rect 31336 60902 33336 60931
rect 31336 60856 31349 60902
rect 33323 60856 33336 60902
rect 31336 60827 33336 60856
rect 44799 61499 45323 61528
rect 51789 61798 53789 61827
rect 51789 61752 51802 61798
rect 53776 61752 53789 61798
rect 51789 61723 53789 61752
rect 51789 61574 53789 61603
rect 51789 61528 51802 61574
rect 53776 61528 53789 61574
rect 51789 61499 53789 61528
rect 44799 61350 45323 61379
rect 44799 61304 44812 61350
rect 44858 61304 44925 61350
rect 44971 61304 45038 61350
rect 45084 61304 45151 61350
rect 45197 61304 45264 61350
rect 45310 61304 45323 61350
rect 44799 61275 45323 61304
rect 51789 61350 53789 61379
rect 51789 61304 51802 61350
rect 53776 61304 53789 61350
rect 51789 61275 53789 61304
rect 35260 61039 36360 61052
rect 35260 60993 35273 61039
rect 35523 60993 35580 61039
rect 35626 60993 35683 61039
rect 35729 60993 35786 61039
rect 35832 60993 35889 61039
rect 35935 60993 35992 61039
rect 36038 60993 36095 61039
rect 36141 60993 36198 61039
rect 36244 60993 36301 61039
rect 36347 60993 36360 61039
rect 35260 60964 36360 60993
rect 36841 61039 37501 61052
rect 36841 60993 36854 61039
rect 36900 60993 36971 61039
rect 37017 60993 37088 61039
rect 37134 60993 37206 61039
rect 37252 60993 37324 61039
rect 37370 60993 37442 61039
rect 37488 60993 37501 61039
rect 36841 60964 37501 60993
rect 44799 61126 45323 61155
rect 44799 61080 44812 61126
rect 44858 61080 44925 61126
rect 44971 61080 45038 61126
rect 45084 61080 45151 61126
rect 45197 61080 45264 61126
rect 45310 61080 45323 61126
rect 54750 61350 55849 61383
rect 54750 61304 54793 61350
rect 54839 61304 54956 61350
rect 55002 61304 55118 61350
rect 55164 61304 55279 61350
rect 55325 61304 55439 61350
rect 55485 61304 55599 61350
rect 55645 61304 55760 61350
rect 55806 61304 55849 61350
rect 54750 61271 55849 61304
rect 44799 61051 45323 61080
rect 31336 60678 33336 60707
rect 31336 60632 31349 60678
rect 33323 60632 33336 60678
rect 35260 60815 36360 60844
rect 35260 60769 35273 60815
rect 35523 60769 35580 60815
rect 35626 60769 35683 60815
rect 35729 60769 35786 60815
rect 35832 60769 35889 60815
rect 35935 60769 35992 60815
rect 36038 60769 36095 60815
rect 36141 60769 36198 60815
rect 36244 60769 36301 60815
rect 36347 60769 36360 60815
rect 35260 60740 36360 60769
rect 31336 60619 33336 60632
rect 48765 61039 49865 61052
rect 48765 60993 48778 61039
rect 48824 60993 48881 61039
rect 48927 60993 48984 61039
rect 49030 60993 49087 61039
rect 49133 60993 49190 61039
rect 49236 60993 49293 61039
rect 49339 60993 49396 61039
rect 49442 60993 49499 61039
rect 49545 60993 49602 61039
rect 49852 60993 49865 61039
rect 48765 60964 49865 60993
rect 36841 60815 37501 60844
rect 36841 60769 36854 60815
rect 36900 60769 36971 60815
rect 37017 60769 37088 60815
rect 37134 60769 37206 60815
rect 37252 60769 37324 60815
rect 37370 60769 37442 60815
rect 37488 60769 37501 60815
rect 36841 60740 37501 60769
rect 39008 60815 39326 60828
rect 39008 60769 39021 60815
rect 39067 60769 39144 60815
rect 39190 60769 39267 60815
rect 39313 60769 39326 60815
rect 39008 60740 39326 60769
rect 44799 60902 45323 60931
rect 44799 60856 44812 60902
rect 44858 60856 44925 60902
rect 44971 60856 45038 60902
rect 45084 60856 45151 60902
rect 45197 60856 45264 60902
rect 45310 60856 45323 60902
rect 44799 60827 45323 60856
rect 48765 60815 49865 60844
rect 48765 60769 48778 60815
rect 48824 60769 48881 60815
rect 48927 60769 48984 60815
rect 49030 60769 49087 60815
rect 49133 60769 49190 60815
rect 49236 60769 49293 60815
rect 49339 60769 49396 60815
rect 49442 60769 49499 60815
rect 49545 60769 49602 60815
rect 49852 60769 49865 60815
rect 48765 60740 49865 60769
rect 35260 60591 36360 60620
rect 35260 60545 35273 60591
rect 35523 60545 35580 60591
rect 35626 60545 35683 60591
rect 35729 60545 35786 60591
rect 35832 60545 35889 60591
rect 35935 60545 35992 60591
rect 36038 60545 36095 60591
rect 36141 60545 36198 60591
rect 36244 60545 36301 60591
rect 36347 60545 36360 60591
rect 35260 60532 36360 60545
rect 36841 60591 37501 60620
rect 36841 60545 36854 60591
rect 36900 60545 36971 60591
rect 37017 60545 37088 60591
rect 37134 60545 37206 60591
rect 37252 60545 37324 60591
rect 37370 60545 37442 60591
rect 37488 60545 37501 60591
rect 36841 60532 37501 60545
rect 39008 60591 39326 60620
rect 39008 60545 39021 60591
rect 39067 60545 39144 60591
rect 39190 60545 39267 60591
rect 39313 60545 39326 60591
rect 39008 60532 39326 60545
rect 44799 60678 45323 60707
rect 44799 60632 44812 60678
rect 44858 60632 44925 60678
rect 44971 60632 45038 60678
rect 45084 60632 45151 60678
rect 45197 60632 45264 60678
rect 45310 60632 45323 60678
rect 44799 60619 45323 60632
rect 51789 61126 53789 61155
rect 51789 61080 51802 61126
rect 53776 61080 53789 61126
rect 51789 61051 53789 61080
rect 51789 60902 53789 60931
rect 51789 60856 51802 60902
rect 53776 60856 53789 60902
rect 51789 60827 53789 60856
rect 51789 60678 53789 60707
rect 48765 60591 49865 60620
rect 48765 60545 48778 60591
rect 48824 60545 48881 60591
rect 48927 60545 48984 60591
rect 49030 60545 49087 60591
rect 49133 60545 49190 60591
rect 49236 60545 49293 60591
rect 49339 60545 49396 60591
rect 49442 60545 49499 60591
rect 49545 60545 49602 60591
rect 49852 60545 49865 60591
rect 51789 60632 51802 60678
rect 53776 60632 53789 60678
rect 51789 60619 53789 60632
rect 48765 60532 49865 60545
rect 29274 60450 30373 60483
rect 29274 60404 29317 60450
rect 29363 60404 29478 60450
rect 29524 60404 29638 60450
rect 29684 60404 29798 60450
rect 29844 60404 29959 60450
rect 30005 60404 30121 60450
rect 30167 60404 30284 60450
rect 30330 60404 30373 60450
rect 29274 60371 30373 60404
rect 54750 60450 55849 60483
rect 54750 60404 54793 60450
rect 54839 60404 54956 60450
rect 55002 60404 55118 60450
rect 55164 60404 55279 60450
rect 55325 60404 55439 60450
rect 55485 60404 55599 60450
rect 55645 60404 55760 60450
rect 55806 60404 55849 60450
rect 54750 60371 55849 60404
rect 35260 60309 36360 60322
rect 31336 60222 33336 60235
rect 31336 60176 31349 60222
rect 33323 60176 33336 60222
rect 35260 60263 35273 60309
rect 35523 60263 35580 60309
rect 35626 60263 35683 60309
rect 35729 60263 35786 60309
rect 35832 60263 35889 60309
rect 35935 60263 35992 60309
rect 36038 60263 36095 60309
rect 36141 60263 36198 60309
rect 36244 60263 36301 60309
rect 36347 60263 36360 60309
rect 35260 60234 36360 60263
rect 36841 60309 37501 60322
rect 36841 60263 36854 60309
rect 36900 60263 36971 60309
rect 37017 60263 37088 60309
rect 37134 60263 37206 60309
rect 37252 60263 37324 60309
rect 37370 60263 37442 60309
rect 37488 60263 37501 60309
rect 36841 60234 37501 60263
rect 39008 60309 39326 60322
rect 39008 60263 39021 60309
rect 39067 60263 39144 60309
rect 39190 60263 39267 60309
rect 39313 60263 39326 60309
rect 39008 60234 39326 60263
rect 48765 60309 49865 60322
rect 31336 60147 33336 60176
rect 31336 59998 33336 60027
rect 31336 59952 31349 59998
rect 33323 59952 33336 59998
rect 31336 59923 33336 59952
rect 31336 59774 33336 59803
rect 31336 59728 31349 59774
rect 33323 59728 33336 59774
rect 31336 59699 33336 59728
rect 29274 59550 30373 59583
rect 29274 59504 29317 59550
rect 29363 59504 29478 59550
rect 29524 59504 29638 59550
rect 29684 59504 29798 59550
rect 29844 59504 29959 59550
rect 30005 59504 30121 59550
rect 30167 59504 30284 59550
rect 30330 59504 30373 59550
rect 29274 59471 30373 59504
rect 35260 60085 36360 60114
rect 35260 60039 35273 60085
rect 35523 60039 35580 60085
rect 35626 60039 35683 60085
rect 35729 60039 35786 60085
rect 35832 60039 35889 60085
rect 35935 60039 35992 60085
rect 36038 60039 36095 60085
rect 36141 60039 36198 60085
rect 36244 60039 36301 60085
rect 36347 60039 36360 60085
rect 35260 60010 36360 60039
rect 36841 60085 37501 60114
rect 36841 60039 36854 60085
rect 36900 60039 36971 60085
rect 37017 60039 37088 60085
rect 37134 60039 37206 60085
rect 37252 60039 37324 60085
rect 37370 60039 37442 60085
rect 37488 60039 37501 60085
rect 36841 60010 37501 60039
rect 48765 60263 48778 60309
rect 48824 60263 48881 60309
rect 48927 60263 48984 60309
rect 49030 60263 49087 60309
rect 49133 60263 49190 60309
rect 49236 60263 49293 60309
rect 49339 60263 49396 60309
rect 49442 60263 49499 60309
rect 49545 60263 49602 60309
rect 49852 60263 49865 60309
rect 44799 60222 45323 60235
rect 48765 60234 49865 60263
rect 44799 60176 44812 60222
rect 44858 60176 44925 60222
rect 44971 60176 45038 60222
rect 45084 60176 45151 60222
rect 45197 60176 45264 60222
rect 45310 60176 45323 60222
rect 44799 60147 45323 60176
rect 39008 60085 39326 60114
rect 39008 60039 39021 60085
rect 39067 60039 39144 60085
rect 39190 60039 39267 60085
rect 39313 60039 39326 60085
rect 39008 60026 39326 60039
rect 51789 60222 53789 60235
rect 44799 59998 45323 60027
rect 44799 59952 44812 59998
rect 44858 59952 44925 59998
rect 44971 59952 45038 59998
rect 45084 59952 45151 59998
rect 45197 59952 45264 59998
rect 45310 59952 45323 59998
rect 44799 59923 45323 59952
rect 48765 60085 49865 60114
rect 48765 60039 48778 60085
rect 48824 60039 48881 60085
rect 48927 60039 48984 60085
rect 49030 60039 49087 60085
rect 49133 60039 49190 60085
rect 49236 60039 49293 60085
rect 49339 60039 49396 60085
rect 49442 60039 49499 60085
rect 49545 60039 49602 60085
rect 49852 60039 49865 60085
rect 48765 60010 49865 60039
rect 51789 60176 51802 60222
rect 53776 60176 53789 60222
rect 51789 60147 53789 60176
rect 35260 59861 36360 59890
rect 35260 59815 35273 59861
rect 35523 59815 35580 59861
rect 35626 59815 35683 59861
rect 35729 59815 35786 59861
rect 35832 59815 35889 59861
rect 35935 59815 35992 59861
rect 36038 59815 36095 59861
rect 36141 59815 36198 59861
rect 36244 59815 36301 59861
rect 36347 59815 36360 59861
rect 35260 59802 36360 59815
rect 36841 59861 37501 59890
rect 36841 59815 36854 59861
rect 36900 59815 36971 59861
rect 37017 59815 37088 59861
rect 37134 59815 37206 59861
rect 37252 59815 37324 59861
rect 37370 59815 37442 59861
rect 37488 59815 37501 59861
rect 36841 59802 37501 59815
rect 48765 59861 49865 59890
rect 48765 59815 48778 59861
rect 48824 59815 48881 59861
rect 48927 59815 48984 59861
rect 49030 59815 49087 59861
rect 49133 59815 49190 59861
rect 49236 59815 49293 59861
rect 49339 59815 49396 59861
rect 49442 59815 49499 59861
rect 49545 59815 49602 59861
rect 49852 59815 49865 59861
rect 44799 59774 45323 59803
rect 48765 59802 49865 59815
rect 44799 59728 44812 59774
rect 44858 59728 44925 59774
rect 44971 59728 45038 59774
rect 45084 59728 45151 59774
rect 45197 59728 45264 59774
rect 45310 59728 45323 59774
rect 31336 59550 33336 59579
rect 31336 59504 31349 59550
rect 33323 59504 33336 59550
rect 31336 59475 33336 59504
rect 31336 59326 33336 59355
rect 31336 59280 31349 59326
rect 33323 59280 33336 59326
rect 31336 59251 33336 59280
rect 31336 59102 33336 59131
rect 31336 59056 31349 59102
rect 33323 59056 33336 59102
rect 31336 59027 33336 59056
rect 44799 59699 45323 59728
rect 51789 59998 53789 60027
rect 51789 59952 51802 59998
rect 53776 59952 53789 59998
rect 51789 59923 53789 59952
rect 51789 59774 53789 59803
rect 51789 59728 51802 59774
rect 53776 59728 53789 59774
rect 51789 59699 53789 59728
rect 44799 59550 45323 59579
rect 44799 59504 44812 59550
rect 44858 59504 44925 59550
rect 44971 59504 45038 59550
rect 45084 59504 45151 59550
rect 45197 59504 45264 59550
rect 45310 59504 45323 59550
rect 44799 59475 45323 59504
rect 51789 59550 53789 59579
rect 51789 59504 51802 59550
rect 53776 59504 53789 59550
rect 51789 59475 53789 59504
rect 35260 59239 36360 59252
rect 35260 59193 35273 59239
rect 35523 59193 35580 59239
rect 35626 59193 35683 59239
rect 35729 59193 35786 59239
rect 35832 59193 35889 59239
rect 35935 59193 35992 59239
rect 36038 59193 36095 59239
rect 36141 59193 36198 59239
rect 36244 59193 36301 59239
rect 36347 59193 36360 59239
rect 35260 59164 36360 59193
rect 36841 59239 37501 59252
rect 36841 59193 36854 59239
rect 36900 59193 36971 59239
rect 37017 59193 37088 59239
rect 37134 59193 37206 59239
rect 37252 59193 37324 59239
rect 37370 59193 37442 59239
rect 37488 59193 37501 59239
rect 36841 59164 37501 59193
rect 44799 59326 45323 59355
rect 44799 59280 44812 59326
rect 44858 59280 44925 59326
rect 44971 59280 45038 59326
rect 45084 59280 45151 59326
rect 45197 59280 45264 59326
rect 45310 59280 45323 59326
rect 54750 59550 55849 59583
rect 54750 59504 54793 59550
rect 54839 59504 54956 59550
rect 55002 59504 55118 59550
rect 55164 59504 55279 59550
rect 55325 59504 55439 59550
rect 55485 59504 55599 59550
rect 55645 59504 55760 59550
rect 55806 59504 55849 59550
rect 54750 59471 55849 59504
rect 44799 59251 45323 59280
rect 31336 58878 33336 58907
rect 31336 58832 31349 58878
rect 33323 58832 33336 58878
rect 35260 59015 36360 59044
rect 35260 58969 35273 59015
rect 35523 58969 35580 59015
rect 35626 58969 35683 59015
rect 35729 58969 35786 59015
rect 35832 58969 35889 59015
rect 35935 58969 35992 59015
rect 36038 58969 36095 59015
rect 36141 58969 36198 59015
rect 36244 58969 36301 59015
rect 36347 58969 36360 59015
rect 35260 58940 36360 58969
rect 31336 58819 33336 58832
rect 48765 59239 49865 59252
rect 48765 59193 48778 59239
rect 48824 59193 48881 59239
rect 48927 59193 48984 59239
rect 49030 59193 49087 59239
rect 49133 59193 49190 59239
rect 49236 59193 49293 59239
rect 49339 59193 49396 59239
rect 49442 59193 49499 59239
rect 49545 59193 49602 59239
rect 49852 59193 49865 59239
rect 48765 59164 49865 59193
rect 36841 59015 37501 59044
rect 36841 58969 36854 59015
rect 36900 58969 36971 59015
rect 37017 58969 37088 59015
rect 37134 58969 37206 59015
rect 37252 58969 37324 59015
rect 37370 58969 37442 59015
rect 37488 58969 37501 59015
rect 36841 58940 37501 58969
rect 39008 59015 39326 59028
rect 39008 58969 39021 59015
rect 39067 58969 39144 59015
rect 39190 58969 39267 59015
rect 39313 58969 39326 59015
rect 39008 58940 39326 58969
rect 44799 59102 45323 59131
rect 44799 59056 44812 59102
rect 44858 59056 44925 59102
rect 44971 59056 45038 59102
rect 45084 59056 45151 59102
rect 45197 59056 45264 59102
rect 45310 59056 45323 59102
rect 44799 59027 45323 59056
rect 48765 59015 49865 59044
rect 48765 58969 48778 59015
rect 48824 58969 48881 59015
rect 48927 58969 48984 59015
rect 49030 58969 49087 59015
rect 49133 58969 49190 59015
rect 49236 58969 49293 59015
rect 49339 58969 49396 59015
rect 49442 58969 49499 59015
rect 49545 58969 49602 59015
rect 49852 58969 49865 59015
rect 48765 58940 49865 58969
rect 35260 58791 36360 58820
rect 35260 58745 35273 58791
rect 35523 58745 35580 58791
rect 35626 58745 35683 58791
rect 35729 58745 35786 58791
rect 35832 58745 35889 58791
rect 35935 58745 35992 58791
rect 36038 58745 36095 58791
rect 36141 58745 36198 58791
rect 36244 58745 36301 58791
rect 36347 58745 36360 58791
rect 35260 58732 36360 58745
rect 36841 58791 37501 58820
rect 36841 58745 36854 58791
rect 36900 58745 36971 58791
rect 37017 58745 37088 58791
rect 37134 58745 37206 58791
rect 37252 58745 37324 58791
rect 37370 58745 37442 58791
rect 37488 58745 37501 58791
rect 36841 58732 37501 58745
rect 39008 58791 39326 58820
rect 39008 58745 39021 58791
rect 39067 58745 39144 58791
rect 39190 58745 39267 58791
rect 39313 58745 39326 58791
rect 39008 58732 39326 58745
rect 44799 58878 45323 58907
rect 44799 58832 44812 58878
rect 44858 58832 44925 58878
rect 44971 58832 45038 58878
rect 45084 58832 45151 58878
rect 45197 58832 45264 58878
rect 45310 58832 45323 58878
rect 44799 58819 45323 58832
rect 51789 59326 53789 59355
rect 51789 59280 51802 59326
rect 53776 59280 53789 59326
rect 51789 59251 53789 59280
rect 51789 59102 53789 59131
rect 51789 59056 51802 59102
rect 53776 59056 53789 59102
rect 51789 59027 53789 59056
rect 51789 58878 53789 58907
rect 48765 58791 49865 58820
rect 48765 58745 48778 58791
rect 48824 58745 48881 58791
rect 48927 58745 48984 58791
rect 49030 58745 49087 58791
rect 49133 58745 49190 58791
rect 49236 58745 49293 58791
rect 49339 58745 49396 58791
rect 49442 58745 49499 58791
rect 49545 58745 49602 58791
rect 49852 58745 49865 58791
rect 51789 58832 51802 58878
rect 53776 58832 53789 58878
rect 51789 58819 53789 58832
rect 48765 58732 49865 58745
rect 29274 58650 30373 58683
rect 29274 58604 29317 58650
rect 29363 58604 29478 58650
rect 29524 58604 29638 58650
rect 29684 58604 29798 58650
rect 29844 58604 29959 58650
rect 30005 58604 30121 58650
rect 30167 58604 30284 58650
rect 30330 58604 30373 58650
rect 29274 58571 30373 58604
rect 54750 58650 55849 58683
rect 54750 58604 54793 58650
rect 54839 58604 54956 58650
rect 55002 58604 55118 58650
rect 55164 58604 55279 58650
rect 55325 58604 55439 58650
rect 55485 58604 55599 58650
rect 55645 58604 55760 58650
rect 55806 58604 55849 58650
rect 54750 58571 55849 58604
rect 35260 58509 36360 58522
rect 31336 58422 33336 58435
rect 31336 58376 31349 58422
rect 33323 58376 33336 58422
rect 35260 58463 35273 58509
rect 35523 58463 35580 58509
rect 35626 58463 35683 58509
rect 35729 58463 35786 58509
rect 35832 58463 35889 58509
rect 35935 58463 35992 58509
rect 36038 58463 36095 58509
rect 36141 58463 36198 58509
rect 36244 58463 36301 58509
rect 36347 58463 36360 58509
rect 35260 58434 36360 58463
rect 36841 58509 37501 58522
rect 36841 58463 36854 58509
rect 36900 58463 36971 58509
rect 37017 58463 37088 58509
rect 37134 58463 37206 58509
rect 37252 58463 37324 58509
rect 37370 58463 37442 58509
rect 37488 58463 37501 58509
rect 36841 58434 37501 58463
rect 39008 58509 39326 58522
rect 39008 58463 39021 58509
rect 39067 58463 39144 58509
rect 39190 58463 39267 58509
rect 39313 58463 39326 58509
rect 39008 58434 39326 58463
rect 48765 58509 49865 58522
rect 31336 58347 33336 58376
rect 31336 58198 33336 58227
rect 31336 58152 31349 58198
rect 33323 58152 33336 58198
rect 31336 58123 33336 58152
rect 31336 57974 33336 58003
rect 31336 57928 31349 57974
rect 33323 57928 33336 57974
rect 31336 57899 33336 57928
rect 29274 57750 30373 57783
rect 29274 57704 29317 57750
rect 29363 57704 29478 57750
rect 29524 57704 29638 57750
rect 29684 57704 29798 57750
rect 29844 57704 29959 57750
rect 30005 57704 30121 57750
rect 30167 57704 30284 57750
rect 30330 57704 30373 57750
rect 29274 57671 30373 57704
rect 35260 58285 36360 58314
rect 35260 58239 35273 58285
rect 35523 58239 35580 58285
rect 35626 58239 35683 58285
rect 35729 58239 35786 58285
rect 35832 58239 35889 58285
rect 35935 58239 35992 58285
rect 36038 58239 36095 58285
rect 36141 58239 36198 58285
rect 36244 58239 36301 58285
rect 36347 58239 36360 58285
rect 35260 58210 36360 58239
rect 36841 58285 37501 58314
rect 36841 58239 36854 58285
rect 36900 58239 36971 58285
rect 37017 58239 37088 58285
rect 37134 58239 37206 58285
rect 37252 58239 37324 58285
rect 37370 58239 37442 58285
rect 37488 58239 37501 58285
rect 36841 58210 37501 58239
rect 48765 58463 48778 58509
rect 48824 58463 48881 58509
rect 48927 58463 48984 58509
rect 49030 58463 49087 58509
rect 49133 58463 49190 58509
rect 49236 58463 49293 58509
rect 49339 58463 49396 58509
rect 49442 58463 49499 58509
rect 49545 58463 49602 58509
rect 49852 58463 49865 58509
rect 44799 58422 45323 58435
rect 48765 58434 49865 58463
rect 44799 58376 44812 58422
rect 44858 58376 44925 58422
rect 44971 58376 45038 58422
rect 45084 58376 45151 58422
rect 45197 58376 45264 58422
rect 45310 58376 45323 58422
rect 44799 58347 45323 58376
rect 39008 58285 39326 58314
rect 39008 58239 39021 58285
rect 39067 58239 39144 58285
rect 39190 58239 39267 58285
rect 39313 58239 39326 58285
rect 39008 58226 39326 58239
rect 51789 58422 53789 58435
rect 44799 58198 45323 58227
rect 44799 58152 44812 58198
rect 44858 58152 44925 58198
rect 44971 58152 45038 58198
rect 45084 58152 45151 58198
rect 45197 58152 45264 58198
rect 45310 58152 45323 58198
rect 44799 58123 45323 58152
rect 48765 58285 49865 58314
rect 48765 58239 48778 58285
rect 48824 58239 48881 58285
rect 48927 58239 48984 58285
rect 49030 58239 49087 58285
rect 49133 58239 49190 58285
rect 49236 58239 49293 58285
rect 49339 58239 49396 58285
rect 49442 58239 49499 58285
rect 49545 58239 49602 58285
rect 49852 58239 49865 58285
rect 48765 58210 49865 58239
rect 51789 58376 51802 58422
rect 53776 58376 53789 58422
rect 51789 58347 53789 58376
rect 35260 58061 36360 58090
rect 35260 58015 35273 58061
rect 35523 58015 35580 58061
rect 35626 58015 35683 58061
rect 35729 58015 35786 58061
rect 35832 58015 35889 58061
rect 35935 58015 35992 58061
rect 36038 58015 36095 58061
rect 36141 58015 36198 58061
rect 36244 58015 36301 58061
rect 36347 58015 36360 58061
rect 35260 58002 36360 58015
rect 36841 58061 37501 58090
rect 36841 58015 36854 58061
rect 36900 58015 36971 58061
rect 37017 58015 37088 58061
rect 37134 58015 37206 58061
rect 37252 58015 37324 58061
rect 37370 58015 37442 58061
rect 37488 58015 37501 58061
rect 36841 58002 37501 58015
rect 48765 58061 49865 58090
rect 48765 58015 48778 58061
rect 48824 58015 48881 58061
rect 48927 58015 48984 58061
rect 49030 58015 49087 58061
rect 49133 58015 49190 58061
rect 49236 58015 49293 58061
rect 49339 58015 49396 58061
rect 49442 58015 49499 58061
rect 49545 58015 49602 58061
rect 49852 58015 49865 58061
rect 44799 57974 45323 58003
rect 48765 58002 49865 58015
rect 44799 57928 44812 57974
rect 44858 57928 44925 57974
rect 44971 57928 45038 57974
rect 45084 57928 45151 57974
rect 45197 57928 45264 57974
rect 45310 57928 45323 57974
rect 31336 57750 33336 57779
rect 31336 57704 31349 57750
rect 33323 57704 33336 57750
rect 31336 57675 33336 57704
rect 31336 57526 33336 57555
rect 31336 57480 31349 57526
rect 33323 57480 33336 57526
rect 31336 57451 33336 57480
rect 31336 57302 33336 57331
rect 31336 57256 31349 57302
rect 33323 57256 33336 57302
rect 31336 57227 33336 57256
rect 44799 57899 45323 57928
rect 51789 58198 53789 58227
rect 51789 58152 51802 58198
rect 53776 58152 53789 58198
rect 51789 58123 53789 58152
rect 51789 57974 53789 58003
rect 51789 57928 51802 57974
rect 53776 57928 53789 57974
rect 51789 57899 53789 57928
rect 44799 57750 45323 57779
rect 44799 57704 44812 57750
rect 44858 57704 44925 57750
rect 44971 57704 45038 57750
rect 45084 57704 45151 57750
rect 45197 57704 45264 57750
rect 45310 57704 45323 57750
rect 44799 57675 45323 57704
rect 51789 57750 53789 57779
rect 51789 57704 51802 57750
rect 53776 57704 53789 57750
rect 51789 57675 53789 57704
rect 35260 57439 36360 57452
rect 35260 57393 35273 57439
rect 35523 57393 35580 57439
rect 35626 57393 35683 57439
rect 35729 57393 35786 57439
rect 35832 57393 35889 57439
rect 35935 57393 35992 57439
rect 36038 57393 36095 57439
rect 36141 57393 36198 57439
rect 36244 57393 36301 57439
rect 36347 57393 36360 57439
rect 35260 57364 36360 57393
rect 36841 57439 37501 57452
rect 36841 57393 36854 57439
rect 36900 57393 36971 57439
rect 37017 57393 37088 57439
rect 37134 57393 37206 57439
rect 37252 57393 37324 57439
rect 37370 57393 37442 57439
rect 37488 57393 37501 57439
rect 36841 57364 37501 57393
rect 44799 57526 45323 57555
rect 44799 57480 44812 57526
rect 44858 57480 44925 57526
rect 44971 57480 45038 57526
rect 45084 57480 45151 57526
rect 45197 57480 45264 57526
rect 45310 57480 45323 57526
rect 54750 57750 55849 57783
rect 54750 57704 54793 57750
rect 54839 57704 54956 57750
rect 55002 57704 55118 57750
rect 55164 57704 55279 57750
rect 55325 57704 55439 57750
rect 55485 57704 55599 57750
rect 55645 57704 55760 57750
rect 55806 57704 55849 57750
rect 54750 57671 55849 57704
rect 44799 57451 45323 57480
rect 31336 57078 33336 57107
rect 31336 57032 31349 57078
rect 33323 57032 33336 57078
rect 35260 57215 36360 57244
rect 35260 57169 35273 57215
rect 35523 57169 35580 57215
rect 35626 57169 35683 57215
rect 35729 57169 35786 57215
rect 35832 57169 35889 57215
rect 35935 57169 35992 57215
rect 36038 57169 36095 57215
rect 36141 57169 36198 57215
rect 36244 57169 36301 57215
rect 36347 57169 36360 57215
rect 35260 57140 36360 57169
rect 31336 57019 33336 57032
rect 48765 57439 49865 57452
rect 48765 57393 48778 57439
rect 48824 57393 48881 57439
rect 48927 57393 48984 57439
rect 49030 57393 49087 57439
rect 49133 57393 49190 57439
rect 49236 57393 49293 57439
rect 49339 57393 49396 57439
rect 49442 57393 49499 57439
rect 49545 57393 49602 57439
rect 49852 57393 49865 57439
rect 48765 57364 49865 57393
rect 36841 57215 37501 57244
rect 36841 57169 36854 57215
rect 36900 57169 36971 57215
rect 37017 57169 37088 57215
rect 37134 57169 37206 57215
rect 37252 57169 37324 57215
rect 37370 57169 37442 57215
rect 37488 57169 37501 57215
rect 36841 57140 37501 57169
rect 39008 57215 39326 57228
rect 39008 57169 39021 57215
rect 39067 57169 39144 57215
rect 39190 57169 39267 57215
rect 39313 57169 39326 57215
rect 39008 57140 39326 57169
rect 44799 57302 45323 57331
rect 44799 57256 44812 57302
rect 44858 57256 44925 57302
rect 44971 57256 45038 57302
rect 45084 57256 45151 57302
rect 45197 57256 45264 57302
rect 45310 57256 45323 57302
rect 44799 57227 45323 57256
rect 48765 57215 49865 57244
rect 48765 57169 48778 57215
rect 48824 57169 48881 57215
rect 48927 57169 48984 57215
rect 49030 57169 49087 57215
rect 49133 57169 49190 57215
rect 49236 57169 49293 57215
rect 49339 57169 49396 57215
rect 49442 57169 49499 57215
rect 49545 57169 49602 57215
rect 49852 57169 49865 57215
rect 48765 57140 49865 57169
rect 35260 56991 36360 57020
rect 35260 56945 35273 56991
rect 35523 56945 35580 56991
rect 35626 56945 35683 56991
rect 35729 56945 35786 56991
rect 35832 56945 35889 56991
rect 35935 56945 35992 56991
rect 36038 56945 36095 56991
rect 36141 56945 36198 56991
rect 36244 56945 36301 56991
rect 36347 56945 36360 56991
rect 35260 56932 36360 56945
rect 36841 56991 37501 57020
rect 36841 56945 36854 56991
rect 36900 56945 36971 56991
rect 37017 56945 37088 56991
rect 37134 56945 37206 56991
rect 37252 56945 37324 56991
rect 37370 56945 37442 56991
rect 37488 56945 37501 56991
rect 36841 56932 37501 56945
rect 39008 56991 39326 57020
rect 39008 56945 39021 56991
rect 39067 56945 39144 56991
rect 39190 56945 39267 56991
rect 39313 56945 39326 56991
rect 39008 56932 39326 56945
rect 44799 57078 45323 57107
rect 44799 57032 44812 57078
rect 44858 57032 44925 57078
rect 44971 57032 45038 57078
rect 45084 57032 45151 57078
rect 45197 57032 45264 57078
rect 45310 57032 45323 57078
rect 44799 57019 45323 57032
rect 51789 57526 53789 57555
rect 51789 57480 51802 57526
rect 53776 57480 53789 57526
rect 51789 57451 53789 57480
rect 51789 57302 53789 57331
rect 51789 57256 51802 57302
rect 53776 57256 53789 57302
rect 51789 57227 53789 57256
rect 51789 57078 53789 57107
rect 48765 56991 49865 57020
rect 48765 56945 48778 56991
rect 48824 56945 48881 56991
rect 48927 56945 48984 56991
rect 49030 56945 49087 56991
rect 49133 56945 49190 56991
rect 49236 56945 49293 56991
rect 49339 56945 49396 56991
rect 49442 56945 49499 56991
rect 49545 56945 49602 56991
rect 49852 56945 49865 56991
rect 51789 57032 51802 57078
rect 53776 57032 53789 57078
rect 51789 57019 53789 57032
rect 48765 56932 49865 56945
rect 29274 56850 30373 56883
rect 29274 56804 29317 56850
rect 29363 56804 29478 56850
rect 29524 56804 29638 56850
rect 29684 56804 29798 56850
rect 29844 56804 29959 56850
rect 30005 56804 30121 56850
rect 30167 56804 30284 56850
rect 30330 56804 30373 56850
rect 29274 56771 30373 56804
rect 54750 56850 55849 56883
rect 54750 56804 54793 56850
rect 54839 56804 54956 56850
rect 55002 56804 55118 56850
rect 55164 56804 55279 56850
rect 55325 56804 55439 56850
rect 55485 56804 55599 56850
rect 55645 56804 55760 56850
rect 55806 56804 55849 56850
rect 54750 56771 55849 56804
rect 35260 56709 36360 56722
rect 31336 56622 33336 56635
rect 31336 56576 31349 56622
rect 33323 56576 33336 56622
rect 35260 56663 35273 56709
rect 35523 56663 35580 56709
rect 35626 56663 35683 56709
rect 35729 56663 35786 56709
rect 35832 56663 35889 56709
rect 35935 56663 35992 56709
rect 36038 56663 36095 56709
rect 36141 56663 36198 56709
rect 36244 56663 36301 56709
rect 36347 56663 36360 56709
rect 35260 56634 36360 56663
rect 36841 56709 37501 56722
rect 36841 56663 36854 56709
rect 36900 56663 36971 56709
rect 37017 56663 37088 56709
rect 37134 56663 37206 56709
rect 37252 56663 37324 56709
rect 37370 56663 37442 56709
rect 37488 56663 37501 56709
rect 36841 56634 37501 56663
rect 39008 56709 39326 56722
rect 39008 56663 39021 56709
rect 39067 56663 39144 56709
rect 39190 56663 39267 56709
rect 39313 56663 39326 56709
rect 39008 56634 39326 56663
rect 48765 56709 49865 56722
rect 31336 56547 33336 56576
rect 31336 56398 33336 56427
rect 31336 56352 31349 56398
rect 33323 56352 33336 56398
rect 31336 56323 33336 56352
rect 31336 56174 33336 56203
rect 31336 56128 31349 56174
rect 33323 56128 33336 56174
rect 31336 56099 33336 56128
rect 29274 55950 30373 55983
rect 29274 55904 29317 55950
rect 29363 55904 29478 55950
rect 29524 55904 29638 55950
rect 29684 55904 29798 55950
rect 29844 55904 29959 55950
rect 30005 55904 30121 55950
rect 30167 55904 30284 55950
rect 30330 55904 30373 55950
rect 29274 55871 30373 55904
rect 35260 56485 36360 56514
rect 35260 56439 35273 56485
rect 35523 56439 35580 56485
rect 35626 56439 35683 56485
rect 35729 56439 35786 56485
rect 35832 56439 35889 56485
rect 35935 56439 35992 56485
rect 36038 56439 36095 56485
rect 36141 56439 36198 56485
rect 36244 56439 36301 56485
rect 36347 56439 36360 56485
rect 35260 56410 36360 56439
rect 36841 56485 37501 56514
rect 36841 56439 36854 56485
rect 36900 56439 36971 56485
rect 37017 56439 37088 56485
rect 37134 56439 37206 56485
rect 37252 56439 37324 56485
rect 37370 56439 37442 56485
rect 37488 56439 37501 56485
rect 36841 56410 37501 56439
rect 48765 56663 48778 56709
rect 48824 56663 48881 56709
rect 48927 56663 48984 56709
rect 49030 56663 49087 56709
rect 49133 56663 49190 56709
rect 49236 56663 49293 56709
rect 49339 56663 49396 56709
rect 49442 56663 49499 56709
rect 49545 56663 49602 56709
rect 49852 56663 49865 56709
rect 44799 56622 45323 56635
rect 48765 56634 49865 56663
rect 44799 56576 44812 56622
rect 44858 56576 44925 56622
rect 44971 56576 45038 56622
rect 45084 56576 45151 56622
rect 45197 56576 45264 56622
rect 45310 56576 45323 56622
rect 44799 56547 45323 56576
rect 39008 56485 39326 56514
rect 39008 56439 39021 56485
rect 39067 56439 39144 56485
rect 39190 56439 39267 56485
rect 39313 56439 39326 56485
rect 39008 56426 39326 56439
rect 51789 56622 53789 56635
rect 44799 56398 45323 56427
rect 44799 56352 44812 56398
rect 44858 56352 44925 56398
rect 44971 56352 45038 56398
rect 45084 56352 45151 56398
rect 45197 56352 45264 56398
rect 45310 56352 45323 56398
rect 44799 56323 45323 56352
rect 48765 56485 49865 56514
rect 48765 56439 48778 56485
rect 48824 56439 48881 56485
rect 48927 56439 48984 56485
rect 49030 56439 49087 56485
rect 49133 56439 49190 56485
rect 49236 56439 49293 56485
rect 49339 56439 49396 56485
rect 49442 56439 49499 56485
rect 49545 56439 49602 56485
rect 49852 56439 49865 56485
rect 48765 56410 49865 56439
rect 51789 56576 51802 56622
rect 53776 56576 53789 56622
rect 51789 56547 53789 56576
rect 35260 56261 36360 56290
rect 35260 56215 35273 56261
rect 35523 56215 35580 56261
rect 35626 56215 35683 56261
rect 35729 56215 35786 56261
rect 35832 56215 35889 56261
rect 35935 56215 35992 56261
rect 36038 56215 36095 56261
rect 36141 56215 36198 56261
rect 36244 56215 36301 56261
rect 36347 56215 36360 56261
rect 35260 56202 36360 56215
rect 36841 56261 37501 56290
rect 36841 56215 36854 56261
rect 36900 56215 36971 56261
rect 37017 56215 37088 56261
rect 37134 56215 37206 56261
rect 37252 56215 37324 56261
rect 37370 56215 37442 56261
rect 37488 56215 37501 56261
rect 36841 56202 37501 56215
rect 48765 56261 49865 56290
rect 48765 56215 48778 56261
rect 48824 56215 48881 56261
rect 48927 56215 48984 56261
rect 49030 56215 49087 56261
rect 49133 56215 49190 56261
rect 49236 56215 49293 56261
rect 49339 56215 49396 56261
rect 49442 56215 49499 56261
rect 49545 56215 49602 56261
rect 49852 56215 49865 56261
rect 44799 56174 45323 56203
rect 48765 56202 49865 56215
rect 44799 56128 44812 56174
rect 44858 56128 44925 56174
rect 44971 56128 45038 56174
rect 45084 56128 45151 56174
rect 45197 56128 45264 56174
rect 45310 56128 45323 56174
rect 31336 55950 33336 55979
rect 31336 55904 31349 55950
rect 33323 55904 33336 55950
rect 31336 55875 33336 55904
rect 31336 55726 33336 55755
rect 31336 55680 31349 55726
rect 33323 55680 33336 55726
rect 31336 55651 33336 55680
rect 31336 55502 33336 55531
rect 31336 55456 31349 55502
rect 33323 55456 33336 55502
rect 31336 55427 33336 55456
rect 44799 56099 45323 56128
rect 51789 56398 53789 56427
rect 51789 56352 51802 56398
rect 53776 56352 53789 56398
rect 51789 56323 53789 56352
rect 51789 56174 53789 56203
rect 51789 56128 51802 56174
rect 53776 56128 53789 56174
rect 51789 56099 53789 56128
rect 44799 55950 45323 55979
rect 44799 55904 44812 55950
rect 44858 55904 44925 55950
rect 44971 55904 45038 55950
rect 45084 55904 45151 55950
rect 45197 55904 45264 55950
rect 45310 55904 45323 55950
rect 44799 55875 45323 55904
rect 51789 55950 53789 55979
rect 51789 55904 51802 55950
rect 53776 55904 53789 55950
rect 51789 55875 53789 55904
rect 35260 55639 36360 55652
rect 35260 55593 35273 55639
rect 35523 55593 35580 55639
rect 35626 55593 35683 55639
rect 35729 55593 35786 55639
rect 35832 55593 35889 55639
rect 35935 55593 35992 55639
rect 36038 55593 36095 55639
rect 36141 55593 36198 55639
rect 36244 55593 36301 55639
rect 36347 55593 36360 55639
rect 35260 55564 36360 55593
rect 36841 55639 37501 55652
rect 36841 55593 36854 55639
rect 36900 55593 36971 55639
rect 37017 55593 37088 55639
rect 37134 55593 37206 55639
rect 37252 55593 37324 55639
rect 37370 55593 37442 55639
rect 37488 55593 37501 55639
rect 36841 55564 37501 55593
rect 44799 55726 45323 55755
rect 44799 55680 44812 55726
rect 44858 55680 44925 55726
rect 44971 55680 45038 55726
rect 45084 55680 45151 55726
rect 45197 55680 45264 55726
rect 45310 55680 45323 55726
rect 54750 55950 55849 55983
rect 54750 55904 54793 55950
rect 54839 55904 54956 55950
rect 55002 55904 55118 55950
rect 55164 55904 55279 55950
rect 55325 55904 55439 55950
rect 55485 55904 55599 55950
rect 55645 55904 55760 55950
rect 55806 55904 55849 55950
rect 54750 55871 55849 55904
rect 44799 55651 45323 55680
rect 31336 55278 33336 55307
rect 31336 55232 31349 55278
rect 33323 55232 33336 55278
rect 35260 55415 36360 55444
rect 35260 55369 35273 55415
rect 35523 55369 35580 55415
rect 35626 55369 35683 55415
rect 35729 55369 35786 55415
rect 35832 55369 35889 55415
rect 35935 55369 35992 55415
rect 36038 55369 36095 55415
rect 36141 55369 36198 55415
rect 36244 55369 36301 55415
rect 36347 55369 36360 55415
rect 35260 55340 36360 55369
rect 31336 55219 33336 55232
rect 48765 55639 49865 55652
rect 48765 55593 48778 55639
rect 48824 55593 48881 55639
rect 48927 55593 48984 55639
rect 49030 55593 49087 55639
rect 49133 55593 49190 55639
rect 49236 55593 49293 55639
rect 49339 55593 49396 55639
rect 49442 55593 49499 55639
rect 49545 55593 49602 55639
rect 49852 55593 49865 55639
rect 48765 55564 49865 55593
rect 36841 55415 37501 55444
rect 36841 55369 36854 55415
rect 36900 55369 36971 55415
rect 37017 55369 37088 55415
rect 37134 55369 37206 55415
rect 37252 55369 37324 55415
rect 37370 55369 37442 55415
rect 37488 55369 37501 55415
rect 36841 55340 37501 55369
rect 39008 55415 39326 55428
rect 39008 55369 39021 55415
rect 39067 55369 39144 55415
rect 39190 55369 39267 55415
rect 39313 55369 39326 55415
rect 39008 55340 39326 55369
rect 44799 55502 45323 55531
rect 44799 55456 44812 55502
rect 44858 55456 44925 55502
rect 44971 55456 45038 55502
rect 45084 55456 45151 55502
rect 45197 55456 45264 55502
rect 45310 55456 45323 55502
rect 44799 55427 45323 55456
rect 48765 55415 49865 55444
rect 48765 55369 48778 55415
rect 48824 55369 48881 55415
rect 48927 55369 48984 55415
rect 49030 55369 49087 55415
rect 49133 55369 49190 55415
rect 49236 55369 49293 55415
rect 49339 55369 49396 55415
rect 49442 55369 49499 55415
rect 49545 55369 49602 55415
rect 49852 55369 49865 55415
rect 48765 55340 49865 55369
rect 35260 55191 36360 55220
rect 35260 55145 35273 55191
rect 35523 55145 35580 55191
rect 35626 55145 35683 55191
rect 35729 55145 35786 55191
rect 35832 55145 35889 55191
rect 35935 55145 35992 55191
rect 36038 55145 36095 55191
rect 36141 55145 36198 55191
rect 36244 55145 36301 55191
rect 36347 55145 36360 55191
rect 35260 55132 36360 55145
rect 36841 55191 37501 55220
rect 36841 55145 36854 55191
rect 36900 55145 36971 55191
rect 37017 55145 37088 55191
rect 37134 55145 37206 55191
rect 37252 55145 37324 55191
rect 37370 55145 37442 55191
rect 37488 55145 37501 55191
rect 36841 55132 37501 55145
rect 39008 55191 39326 55220
rect 39008 55145 39021 55191
rect 39067 55145 39144 55191
rect 39190 55145 39267 55191
rect 39313 55145 39326 55191
rect 39008 55132 39326 55145
rect 44799 55278 45323 55307
rect 44799 55232 44812 55278
rect 44858 55232 44925 55278
rect 44971 55232 45038 55278
rect 45084 55232 45151 55278
rect 45197 55232 45264 55278
rect 45310 55232 45323 55278
rect 44799 55219 45323 55232
rect 51789 55726 53789 55755
rect 51789 55680 51802 55726
rect 53776 55680 53789 55726
rect 51789 55651 53789 55680
rect 51789 55502 53789 55531
rect 51789 55456 51802 55502
rect 53776 55456 53789 55502
rect 51789 55427 53789 55456
rect 51789 55278 53789 55307
rect 48765 55191 49865 55220
rect 48765 55145 48778 55191
rect 48824 55145 48881 55191
rect 48927 55145 48984 55191
rect 49030 55145 49087 55191
rect 49133 55145 49190 55191
rect 49236 55145 49293 55191
rect 49339 55145 49396 55191
rect 49442 55145 49499 55191
rect 49545 55145 49602 55191
rect 49852 55145 49865 55191
rect 51789 55232 51802 55278
rect 53776 55232 53789 55278
rect 51789 55219 53789 55232
rect 48765 55132 49865 55145
rect 29274 55050 30373 55083
rect 29274 55004 29317 55050
rect 29363 55004 29478 55050
rect 29524 55004 29638 55050
rect 29684 55004 29798 55050
rect 29844 55004 29959 55050
rect 30005 55004 30121 55050
rect 30167 55004 30284 55050
rect 30330 55004 30373 55050
rect 29274 54971 30373 55004
rect 54750 55050 55849 55083
rect 54750 55004 54793 55050
rect 54839 55004 54956 55050
rect 55002 55004 55118 55050
rect 55164 55004 55279 55050
rect 55325 55004 55439 55050
rect 55485 55004 55599 55050
rect 55645 55004 55760 55050
rect 55806 55004 55849 55050
rect 54750 54971 55849 55004
rect 35260 54909 36360 54922
rect 31336 54822 33336 54835
rect 31336 54776 31349 54822
rect 33323 54776 33336 54822
rect 35260 54863 35273 54909
rect 35523 54863 35580 54909
rect 35626 54863 35683 54909
rect 35729 54863 35786 54909
rect 35832 54863 35889 54909
rect 35935 54863 35992 54909
rect 36038 54863 36095 54909
rect 36141 54863 36198 54909
rect 36244 54863 36301 54909
rect 36347 54863 36360 54909
rect 35260 54834 36360 54863
rect 36841 54909 37501 54922
rect 36841 54863 36854 54909
rect 36900 54863 36971 54909
rect 37017 54863 37088 54909
rect 37134 54863 37206 54909
rect 37252 54863 37324 54909
rect 37370 54863 37442 54909
rect 37488 54863 37501 54909
rect 36841 54834 37501 54863
rect 39008 54909 39326 54922
rect 39008 54863 39021 54909
rect 39067 54863 39144 54909
rect 39190 54863 39267 54909
rect 39313 54863 39326 54909
rect 39008 54834 39326 54863
rect 48765 54909 49865 54922
rect 31336 54747 33336 54776
rect 31336 54598 33336 54627
rect 31336 54552 31349 54598
rect 33323 54552 33336 54598
rect 31336 54523 33336 54552
rect 31336 54374 33336 54403
rect 31336 54328 31349 54374
rect 33323 54328 33336 54374
rect 31336 54299 33336 54328
rect 29274 54150 30373 54183
rect 29274 54104 29317 54150
rect 29363 54104 29478 54150
rect 29524 54104 29638 54150
rect 29684 54104 29798 54150
rect 29844 54104 29959 54150
rect 30005 54104 30121 54150
rect 30167 54104 30284 54150
rect 30330 54104 30373 54150
rect 29274 54071 30373 54104
rect 35260 54685 36360 54714
rect 35260 54639 35273 54685
rect 35523 54639 35580 54685
rect 35626 54639 35683 54685
rect 35729 54639 35786 54685
rect 35832 54639 35889 54685
rect 35935 54639 35992 54685
rect 36038 54639 36095 54685
rect 36141 54639 36198 54685
rect 36244 54639 36301 54685
rect 36347 54639 36360 54685
rect 35260 54610 36360 54639
rect 36841 54685 37501 54714
rect 36841 54639 36854 54685
rect 36900 54639 36971 54685
rect 37017 54639 37088 54685
rect 37134 54639 37206 54685
rect 37252 54639 37324 54685
rect 37370 54639 37442 54685
rect 37488 54639 37501 54685
rect 36841 54610 37501 54639
rect 48765 54863 48778 54909
rect 48824 54863 48881 54909
rect 48927 54863 48984 54909
rect 49030 54863 49087 54909
rect 49133 54863 49190 54909
rect 49236 54863 49293 54909
rect 49339 54863 49396 54909
rect 49442 54863 49499 54909
rect 49545 54863 49602 54909
rect 49852 54863 49865 54909
rect 44799 54822 45323 54835
rect 48765 54834 49865 54863
rect 44799 54776 44812 54822
rect 44858 54776 44925 54822
rect 44971 54776 45038 54822
rect 45084 54776 45151 54822
rect 45197 54776 45264 54822
rect 45310 54776 45323 54822
rect 44799 54747 45323 54776
rect 39008 54685 39326 54714
rect 39008 54639 39021 54685
rect 39067 54639 39144 54685
rect 39190 54639 39267 54685
rect 39313 54639 39326 54685
rect 39008 54626 39326 54639
rect 51789 54822 53789 54835
rect 44799 54598 45323 54627
rect 44799 54552 44812 54598
rect 44858 54552 44925 54598
rect 44971 54552 45038 54598
rect 45084 54552 45151 54598
rect 45197 54552 45264 54598
rect 45310 54552 45323 54598
rect 44799 54523 45323 54552
rect 48765 54685 49865 54714
rect 48765 54639 48778 54685
rect 48824 54639 48881 54685
rect 48927 54639 48984 54685
rect 49030 54639 49087 54685
rect 49133 54639 49190 54685
rect 49236 54639 49293 54685
rect 49339 54639 49396 54685
rect 49442 54639 49499 54685
rect 49545 54639 49602 54685
rect 49852 54639 49865 54685
rect 48765 54610 49865 54639
rect 51789 54776 51802 54822
rect 53776 54776 53789 54822
rect 51789 54747 53789 54776
rect 35260 54461 36360 54490
rect 35260 54415 35273 54461
rect 35523 54415 35580 54461
rect 35626 54415 35683 54461
rect 35729 54415 35786 54461
rect 35832 54415 35889 54461
rect 35935 54415 35992 54461
rect 36038 54415 36095 54461
rect 36141 54415 36198 54461
rect 36244 54415 36301 54461
rect 36347 54415 36360 54461
rect 35260 54402 36360 54415
rect 36841 54461 37501 54490
rect 36841 54415 36854 54461
rect 36900 54415 36971 54461
rect 37017 54415 37088 54461
rect 37134 54415 37206 54461
rect 37252 54415 37324 54461
rect 37370 54415 37442 54461
rect 37488 54415 37501 54461
rect 36841 54402 37501 54415
rect 48765 54461 49865 54490
rect 48765 54415 48778 54461
rect 48824 54415 48881 54461
rect 48927 54415 48984 54461
rect 49030 54415 49087 54461
rect 49133 54415 49190 54461
rect 49236 54415 49293 54461
rect 49339 54415 49396 54461
rect 49442 54415 49499 54461
rect 49545 54415 49602 54461
rect 49852 54415 49865 54461
rect 44799 54374 45323 54403
rect 48765 54402 49865 54415
rect 44799 54328 44812 54374
rect 44858 54328 44925 54374
rect 44971 54328 45038 54374
rect 45084 54328 45151 54374
rect 45197 54328 45264 54374
rect 45310 54328 45323 54374
rect 31336 54150 33336 54179
rect 31336 54104 31349 54150
rect 33323 54104 33336 54150
rect 31336 54075 33336 54104
rect 31336 53926 33336 53955
rect 31336 53880 31349 53926
rect 33323 53880 33336 53926
rect 31336 53851 33336 53880
rect 31336 53702 33336 53731
rect 31336 53656 31349 53702
rect 33323 53656 33336 53702
rect 31336 53627 33336 53656
rect 44799 54299 45323 54328
rect 51789 54598 53789 54627
rect 51789 54552 51802 54598
rect 53776 54552 53789 54598
rect 51789 54523 53789 54552
rect 51789 54374 53789 54403
rect 51789 54328 51802 54374
rect 53776 54328 53789 54374
rect 51789 54299 53789 54328
rect 44799 54150 45323 54179
rect 44799 54104 44812 54150
rect 44858 54104 44925 54150
rect 44971 54104 45038 54150
rect 45084 54104 45151 54150
rect 45197 54104 45264 54150
rect 45310 54104 45323 54150
rect 44799 54075 45323 54104
rect 51789 54150 53789 54179
rect 51789 54104 51802 54150
rect 53776 54104 53789 54150
rect 51789 54075 53789 54104
rect 35260 53839 36360 53852
rect 35260 53793 35273 53839
rect 35523 53793 35580 53839
rect 35626 53793 35683 53839
rect 35729 53793 35786 53839
rect 35832 53793 35889 53839
rect 35935 53793 35992 53839
rect 36038 53793 36095 53839
rect 36141 53793 36198 53839
rect 36244 53793 36301 53839
rect 36347 53793 36360 53839
rect 35260 53764 36360 53793
rect 36841 53839 37501 53852
rect 36841 53793 36854 53839
rect 36900 53793 36971 53839
rect 37017 53793 37088 53839
rect 37134 53793 37206 53839
rect 37252 53793 37324 53839
rect 37370 53793 37442 53839
rect 37488 53793 37501 53839
rect 36841 53764 37501 53793
rect 44799 53926 45323 53955
rect 44799 53880 44812 53926
rect 44858 53880 44925 53926
rect 44971 53880 45038 53926
rect 45084 53880 45151 53926
rect 45197 53880 45264 53926
rect 45310 53880 45323 53926
rect 54750 54150 55849 54183
rect 54750 54104 54793 54150
rect 54839 54104 54956 54150
rect 55002 54104 55118 54150
rect 55164 54104 55279 54150
rect 55325 54104 55439 54150
rect 55485 54104 55599 54150
rect 55645 54104 55760 54150
rect 55806 54104 55849 54150
rect 54750 54071 55849 54104
rect 44799 53851 45323 53880
rect 31336 53478 33336 53507
rect 31336 53432 31349 53478
rect 33323 53432 33336 53478
rect 35260 53615 36360 53644
rect 35260 53569 35273 53615
rect 35523 53569 35580 53615
rect 35626 53569 35683 53615
rect 35729 53569 35786 53615
rect 35832 53569 35889 53615
rect 35935 53569 35992 53615
rect 36038 53569 36095 53615
rect 36141 53569 36198 53615
rect 36244 53569 36301 53615
rect 36347 53569 36360 53615
rect 35260 53540 36360 53569
rect 31336 53419 33336 53432
rect 48765 53839 49865 53852
rect 48765 53793 48778 53839
rect 48824 53793 48881 53839
rect 48927 53793 48984 53839
rect 49030 53793 49087 53839
rect 49133 53793 49190 53839
rect 49236 53793 49293 53839
rect 49339 53793 49396 53839
rect 49442 53793 49499 53839
rect 49545 53793 49602 53839
rect 49852 53793 49865 53839
rect 48765 53764 49865 53793
rect 36841 53615 37501 53644
rect 36841 53569 36854 53615
rect 36900 53569 36971 53615
rect 37017 53569 37088 53615
rect 37134 53569 37206 53615
rect 37252 53569 37324 53615
rect 37370 53569 37442 53615
rect 37488 53569 37501 53615
rect 36841 53540 37501 53569
rect 39008 53615 39326 53628
rect 39008 53569 39021 53615
rect 39067 53569 39144 53615
rect 39190 53569 39267 53615
rect 39313 53569 39326 53615
rect 39008 53540 39326 53569
rect 44799 53702 45323 53731
rect 44799 53656 44812 53702
rect 44858 53656 44925 53702
rect 44971 53656 45038 53702
rect 45084 53656 45151 53702
rect 45197 53656 45264 53702
rect 45310 53656 45323 53702
rect 44799 53627 45323 53656
rect 48765 53615 49865 53644
rect 48765 53569 48778 53615
rect 48824 53569 48881 53615
rect 48927 53569 48984 53615
rect 49030 53569 49087 53615
rect 49133 53569 49190 53615
rect 49236 53569 49293 53615
rect 49339 53569 49396 53615
rect 49442 53569 49499 53615
rect 49545 53569 49602 53615
rect 49852 53569 49865 53615
rect 48765 53540 49865 53569
rect 35260 53391 36360 53420
rect 35260 53345 35273 53391
rect 35523 53345 35580 53391
rect 35626 53345 35683 53391
rect 35729 53345 35786 53391
rect 35832 53345 35889 53391
rect 35935 53345 35992 53391
rect 36038 53345 36095 53391
rect 36141 53345 36198 53391
rect 36244 53345 36301 53391
rect 36347 53345 36360 53391
rect 35260 53332 36360 53345
rect 36841 53391 37501 53420
rect 36841 53345 36854 53391
rect 36900 53345 36971 53391
rect 37017 53345 37088 53391
rect 37134 53345 37206 53391
rect 37252 53345 37324 53391
rect 37370 53345 37442 53391
rect 37488 53345 37501 53391
rect 36841 53332 37501 53345
rect 39008 53391 39326 53420
rect 39008 53345 39021 53391
rect 39067 53345 39144 53391
rect 39190 53345 39267 53391
rect 39313 53345 39326 53391
rect 39008 53332 39326 53345
rect 44799 53478 45323 53507
rect 44799 53432 44812 53478
rect 44858 53432 44925 53478
rect 44971 53432 45038 53478
rect 45084 53432 45151 53478
rect 45197 53432 45264 53478
rect 45310 53432 45323 53478
rect 44799 53419 45323 53432
rect 51789 53926 53789 53955
rect 51789 53880 51802 53926
rect 53776 53880 53789 53926
rect 51789 53851 53789 53880
rect 51789 53702 53789 53731
rect 51789 53656 51802 53702
rect 53776 53656 53789 53702
rect 51789 53627 53789 53656
rect 51789 53478 53789 53507
rect 48765 53391 49865 53420
rect 48765 53345 48778 53391
rect 48824 53345 48881 53391
rect 48927 53345 48984 53391
rect 49030 53345 49087 53391
rect 49133 53345 49190 53391
rect 49236 53345 49293 53391
rect 49339 53345 49396 53391
rect 49442 53345 49499 53391
rect 49545 53345 49602 53391
rect 49852 53345 49865 53391
rect 51789 53432 51802 53478
rect 53776 53432 53789 53478
rect 51789 53419 53789 53432
rect 48765 53332 49865 53345
rect 29274 53250 30373 53283
rect 29274 53204 29317 53250
rect 29363 53204 29478 53250
rect 29524 53204 29638 53250
rect 29684 53204 29798 53250
rect 29844 53204 29959 53250
rect 30005 53204 30121 53250
rect 30167 53204 30284 53250
rect 30330 53204 30373 53250
rect 29274 53171 30373 53204
rect 54750 53250 55849 53283
rect 54750 53204 54793 53250
rect 54839 53204 54956 53250
rect 55002 53204 55118 53250
rect 55164 53204 55279 53250
rect 55325 53204 55439 53250
rect 55485 53204 55599 53250
rect 55645 53204 55760 53250
rect 55806 53204 55849 53250
rect 54750 53171 55849 53204
rect 35260 53109 36360 53122
rect 31336 53022 33336 53035
rect 31336 52976 31349 53022
rect 33323 52976 33336 53022
rect 35260 53063 35273 53109
rect 35523 53063 35580 53109
rect 35626 53063 35683 53109
rect 35729 53063 35786 53109
rect 35832 53063 35889 53109
rect 35935 53063 35992 53109
rect 36038 53063 36095 53109
rect 36141 53063 36198 53109
rect 36244 53063 36301 53109
rect 36347 53063 36360 53109
rect 35260 53034 36360 53063
rect 36841 53109 37501 53122
rect 36841 53063 36854 53109
rect 36900 53063 36971 53109
rect 37017 53063 37088 53109
rect 37134 53063 37206 53109
rect 37252 53063 37324 53109
rect 37370 53063 37442 53109
rect 37488 53063 37501 53109
rect 36841 53034 37501 53063
rect 39008 53109 39326 53122
rect 39008 53063 39021 53109
rect 39067 53063 39144 53109
rect 39190 53063 39267 53109
rect 39313 53063 39326 53109
rect 39008 53034 39326 53063
rect 48765 53109 49865 53122
rect 31336 52947 33336 52976
rect 31336 52798 33336 52827
rect 31336 52752 31349 52798
rect 33323 52752 33336 52798
rect 31336 52723 33336 52752
rect 31336 52574 33336 52603
rect 31336 52528 31349 52574
rect 33323 52528 33336 52574
rect 31336 52499 33336 52528
rect 29274 52350 30373 52383
rect 29274 52304 29317 52350
rect 29363 52304 29478 52350
rect 29524 52304 29638 52350
rect 29684 52304 29798 52350
rect 29844 52304 29959 52350
rect 30005 52304 30121 52350
rect 30167 52304 30284 52350
rect 30330 52304 30373 52350
rect 29274 52271 30373 52304
rect 35260 52885 36360 52914
rect 35260 52839 35273 52885
rect 35523 52839 35580 52885
rect 35626 52839 35683 52885
rect 35729 52839 35786 52885
rect 35832 52839 35889 52885
rect 35935 52839 35992 52885
rect 36038 52839 36095 52885
rect 36141 52839 36198 52885
rect 36244 52839 36301 52885
rect 36347 52839 36360 52885
rect 35260 52810 36360 52839
rect 36841 52885 37501 52914
rect 36841 52839 36854 52885
rect 36900 52839 36971 52885
rect 37017 52839 37088 52885
rect 37134 52839 37206 52885
rect 37252 52839 37324 52885
rect 37370 52839 37442 52885
rect 37488 52839 37501 52885
rect 36841 52810 37501 52839
rect 48765 53063 48778 53109
rect 48824 53063 48881 53109
rect 48927 53063 48984 53109
rect 49030 53063 49087 53109
rect 49133 53063 49190 53109
rect 49236 53063 49293 53109
rect 49339 53063 49396 53109
rect 49442 53063 49499 53109
rect 49545 53063 49602 53109
rect 49852 53063 49865 53109
rect 44799 53022 45323 53035
rect 48765 53034 49865 53063
rect 44799 52976 44812 53022
rect 44858 52976 44925 53022
rect 44971 52976 45038 53022
rect 45084 52976 45151 53022
rect 45197 52976 45264 53022
rect 45310 52976 45323 53022
rect 44799 52947 45323 52976
rect 39008 52885 39326 52914
rect 39008 52839 39021 52885
rect 39067 52839 39144 52885
rect 39190 52839 39267 52885
rect 39313 52839 39326 52885
rect 39008 52826 39326 52839
rect 51789 53022 53789 53035
rect 44799 52798 45323 52827
rect 44799 52752 44812 52798
rect 44858 52752 44925 52798
rect 44971 52752 45038 52798
rect 45084 52752 45151 52798
rect 45197 52752 45264 52798
rect 45310 52752 45323 52798
rect 44799 52723 45323 52752
rect 48765 52885 49865 52914
rect 48765 52839 48778 52885
rect 48824 52839 48881 52885
rect 48927 52839 48984 52885
rect 49030 52839 49087 52885
rect 49133 52839 49190 52885
rect 49236 52839 49293 52885
rect 49339 52839 49396 52885
rect 49442 52839 49499 52885
rect 49545 52839 49602 52885
rect 49852 52839 49865 52885
rect 48765 52810 49865 52839
rect 51789 52976 51802 53022
rect 53776 52976 53789 53022
rect 51789 52947 53789 52976
rect 35260 52661 36360 52690
rect 35260 52615 35273 52661
rect 35523 52615 35580 52661
rect 35626 52615 35683 52661
rect 35729 52615 35786 52661
rect 35832 52615 35889 52661
rect 35935 52615 35992 52661
rect 36038 52615 36095 52661
rect 36141 52615 36198 52661
rect 36244 52615 36301 52661
rect 36347 52615 36360 52661
rect 35260 52602 36360 52615
rect 36841 52661 37501 52690
rect 36841 52615 36854 52661
rect 36900 52615 36971 52661
rect 37017 52615 37088 52661
rect 37134 52615 37206 52661
rect 37252 52615 37324 52661
rect 37370 52615 37442 52661
rect 37488 52615 37501 52661
rect 36841 52602 37501 52615
rect 48765 52661 49865 52690
rect 48765 52615 48778 52661
rect 48824 52615 48881 52661
rect 48927 52615 48984 52661
rect 49030 52615 49087 52661
rect 49133 52615 49190 52661
rect 49236 52615 49293 52661
rect 49339 52615 49396 52661
rect 49442 52615 49499 52661
rect 49545 52615 49602 52661
rect 49852 52615 49865 52661
rect 44799 52574 45323 52603
rect 48765 52602 49865 52615
rect 44799 52528 44812 52574
rect 44858 52528 44925 52574
rect 44971 52528 45038 52574
rect 45084 52528 45151 52574
rect 45197 52528 45264 52574
rect 45310 52528 45323 52574
rect 31336 52350 33336 52379
rect 31336 52304 31349 52350
rect 33323 52304 33336 52350
rect 31336 52275 33336 52304
rect 31336 52126 33336 52155
rect 31336 52080 31349 52126
rect 33323 52080 33336 52126
rect 31336 52051 33336 52080
rect 31336 51902 33336 51931
rect 31336 51856 31349 51902
rect 33323 51856 33336 51902
rect 31336 51827 33336 51856
rect 44799 52499 45323 52528
rect 51789 52798 53789 52827
rect 51789 52752 51802 52798
rect 53776 52752 53789 52798
rect 51789 52723 53789 52752
rect 51789 52574 53789 52603
rect 51789 52528 51802 52574
rect 53776 52528 53789 52574
rect 51789 52499 53789 52528
rect 44799 52350 45323 52379
rect 44799 52304 44812 52350
rect 44858 52304 44925 52350
rect 44971 52304 45038 52350
rect 45084 52304 45151 52350
rect 45197 52304 45264 52350
rect 45310 52304 45323 52350
rect 44799 52275 45323 52304
rect 51789 52350 53789 52379
rect 51789 52304 51802 52350
rect 53776 52304 53789 52350
rect 51789 52275 53789 52304
rect 35260 52039 36360 52052
rect 35260 51993 35273 52039
rect 35523 51993 35580 52039
rect 35626 51993 35683 52039
rect 35729 51993 35786 52039
rect 35832 51993 35889 52039
rect 35935 51993 35992 52039
rect 36038 51993 36095 52039
rect 36141 51993 36198 52039
rect 36244 51993 36301 52039
rect 36347 51993 36360 52039
rect 35260 51964 36360 51993
rect 36841 52039 37501 52052
rect 36841 51993 36854 52039
rect 36900 51993 36971 52039
rect 37017 51993 37088 52039
rect 37134 51993 37206 52039
rect 37252 51993 37324 52039
rect 37370 51993 37442 52039
rect 37488 51993 37501 52039
rect 36841 51964 37501 51993
rect 44799 52126 45323 52155
rect 44799 52080 44812 52126
rect 44858 52080 44925 52126
rect 44971 52080 45038 52126
rect 45084 52080 45151 52126
rect 45197 52080 45264 52126
rect 45310 52080 45323 52126
rect 54750 52350 55849 52383
rect 54750 52304 54793 52350
rect 54839 52304 54956 52350
rect 55002 52304 55118 52350
rect 55164 52304 55279 52350
rect 55325 52304 55439 52350
rect 55485 52304 55599 52350
rect 55645 52304 55760 52350
rect 55806 52304 55849 52350
rect 54750 52271 55849 52304
rect 44799 52051 45323 52080
rect 31336 51678 33336 51707
rect 31336 51632 31349 51678
rect 33323 51632 33336 51678
rect 35260 51815 36360 51844
rect 35260 51769 35273 51815
rect 35523 51769 35580 51815
rect 35626 51769 35683 51815
rect 35729 51769 35786 51815
rect 35832 51769 35889 51815
rect 35935 51769 35992 51815
rect 36038 51769 36095 51815
rect 36141 51769 36198 51815
rect 36244 51769 36301 51815
rect 36347 51769 36360 51815
rect 35260 51740 36360 51769
rect 31336 51619 33336 51632
rect 48765 52039 49865 52052
rect 48765 51993 48778 52039
rect 48824 51993 48881 52039
rect 48927 51993 48984 52039
rect 49030 51993 49087 52039
rect 49133 51993 49190 52039
rect 49236 51993 49293 52039
rect 49339 51993 49396 52039
rect 49442 51993 49499 52039
rect 49545 51993 49602 52039
rect 49852 51993 49865 52039
rect 48765 51964 49865 51993
rect 36841 51815 37501 51844
rect 36841 51769 36854 51815
rect 36900 51769 36971 51815
rect 37017 51769 37088 51815
rect 37134 51769 37206 51815
rect 37252 51769 37324 51815
rect 37370 51769 37442 51815
rect 37488 51769 37501 51815
rect 36841 51740 37501 51769
rect 39008 51815 39326 51828
rect 39008 51769 39021 51815
rect 39067 51769 39144 51815
rect 39190 51769 39267 51815
rect 39313 51769 39326 51815
rect 39008 51740 39326 51769
rect 44799 51902 45323 51931
rect 44799 51856 44812 51902
rect 44858 51856 44925 51902
rect 44971 51856 45038 51902
rect 45084 51856 45151 51902
rect 45197 51856 45264 51902
rect 45310 51856 45323 51902
rect 44799 51827 45323 51856
rect 48765 51815 49865 51844
rect 48765 51769 48778 51815
rect 48824 51769 48881 51815
rect 48927 51769 48984 51815
rect 49030 51769 49087 51815
rect 49133 51769 49190 51815
rect 49236 51769 49293 51815
rect 49339 51769 49396 51815
rect 49442 51769 49499 51815
rect 49545 51769 49602 51815
rect 49852 51769 49865 51815
rect 48765 51740 49865 51769
rect 35260 51591 36360 51620
rect 35260 51545 35273 51591
rect 35523 51545 35580 51591
rect 35626 51545 35683 51591
rect 35729 51545 35786 51591
rect 35832 51545 35889 51591
rect 35935 51545 35992 51591
rect 36038 51545 36095 51591
rect 36141 51545 36198 51591
rect 36244 51545 36301 51591
rect 36347 51545 36360 51591
rect 35260 51532 36360 51545
rect 36841 51591 37501 51620
rect 36841 51545 36854 51591
rect 36900 51545 36971 51591
rect 37017 51545 37088 51591
rect 37134 51545 37206 51591
rect 37252 51545 37324 51591
rect 37370 51545 37442 51591
rect 37488 51545 37501 51591
rect 36841 51532 37501 51545
rect 39008 51591 39326 51620
rect 39008 51545 39021 51591
rect 39067 51545 39144 51591
rect 39190 51545 39267 51591
rect 39313 51545 39326 51591
rect 39008 51532 39326 51545
rect 44799 51678 45323 51707
rect 44799 51632 44812 51678
rect 44858 51632 44925 51678
rect 44971 51632 45038 51678
rect 45084 51632 45151 51678
rect 45197 51632 45264 51678
rect 45310 51632 45323 51678
rect 44799 51619 45323 51632
rect 51789 52126 53789 52155
rect 51789 52080 51802 52126
rect 53776 52080 53789 52126
rect 51789 52051 53789 52080
rect 51789 51902 53789 51931
rect 51789 51856 51802 51902
rect 53776 51856 53789 51902
rect 51789 51827 53789 51856
rect 51789 51678 53789 51707
rect 48765 51591 49865 51620
rect 48765 51545 48778 51591
rect 48824 51545 48881 51591
rect 48927 51545 48984 51591
rect 49030 51545 49087 51591
rect 49133 51545 49190 51591
rect 49236 51545 49293 51591
rect 49339 51545 49396 51591
rect 49442 51545 49499 51591
rect 49545 51545 49602 51591
rect 49852 51545 49865 51591
rect 51789 51632 51802 51678
rect 53776 51632 53789 51678
rect 51789 51619 53789 51632
rect 48765 51532 49865 51545
rect 29274 51450 30373 51483
rect 29274 51404 29317 51450
rect 29363 51404 29478 51450
rect 29524 51404 29638 51450
rect 29684 51404 29798 51450
rect 29844 51404 29959 51450
rect 30005 51404 30121 51450
rect 30167 51404 30284 51450
rect 30330 51404 30373 51450
rect 29274 51371 30373 51404
rect 54750 51450 55849 51483
rect 54750 51404 54793 51450
rect 54839 51404 54956 51450
rect 55002 51404 55118 51450
rect 55164 51404 55279 51450
rect 55325 51404 55439 51450
rect 55485 51404 55599 51450
rect 55645 51404 55760 51450
rect 55806 51404 55849 51450
rect 54750 51371 55849 51404
rect 35260 51309 36360 51322
rect 31336 51222 33336 51235
rect 31336 51176 31349 51222
rect 33323 51176 33336 51222
rect 35260 51263 35273 51309
rect 35523 51263 35580 51309
rect 35626 51263 35683 51309
rect 35729 51263 35786 51309
rect 35832 51263 35889 51309
rect 35935 51263 35992 51309
rect 36038 51263 36095 51309
rect 36141 51263 36198 51309
rect 36244 51263 36301 51309
rect 36347 51263 36360 51309
rect 35260 51234 36360 51263
rect 36841 51309 37501 51322
rect 36841 51263 36854 51309
rect 36900 51263 36971 51309
rect 37017 51263 37088 51309
rect 37134 51263 37206 51309
rect 37252 51263 37324 51309
rect 37370 51263 37442 51309
rect 37488 51263 37501 51309
rect 36841 51234 37501 51263
rect 39008 51309 39326 51322
rect 39008 51263 39021 51309
rect 39067 51263 39144 51309
rect 39190 51263 39267 51309
rect 39313 51263 39326 51309
rect 39008 51234 39326 51263
rect 48765 51309 49865 51322
rect 31336 51147 33336 51176
rect 31336 50998 33336 51027
rect 31336 50952 31349 50998
rect 33323 50952 33336 50998
rect 31336 50923 33336 50952
rect 31336 50774 33336 50803
rect 31336 50728 31349 50774
rect 33323 50728 33336 50774
rect 31336 50699 33336 50728
rect 29274 50550 30373 50583
rect 29274 50504 29317 50550
rect 29363 50504 29478 50550
rect 29524 50504 29638 50550
rect 29684 50504 29798 50550
rect 29844 50504 29959 50550
rect 30005 50504 30121 50550
rect 30167 50504 30284 50550
rect 30330 50504 30373 50550
rect 29274 50471 30373 50504
rect 35260 51085 36360 51114
rect 35260 51039 35273 51085
rect 35523 51039 35580 51085
rect 35626 51039 35683 51085
rect 35729 51039 35786 51085
rect 35832 51039 35889 51085
rect 35935 51039 35992 51085
rect 36038 51039 36095 51085
rect 36141 51039 36198 51085
rect 36244 51039 36301 51085
rect 36347 51039 36360 51085
rect 35260 51010 36360 51039
rect 36841 51085 37501 51114
rect 36841 51039 36854 51085
rect 36900 51039 36971 51085
rect 37017 51039 37088 51085
rect 37134 51039 37206 51085
rect 37252 51039 37324 51085
rect 37370 51039 37442 51085
rect 37488 51039 37501 51085
rect 36841 51010 37501 51039
rect 48765 51263 48778 51309
rect 48824 51263 48881 51309
rect 48927 51263 48984 51309
rect 49030 51263 49087 51309
rect 49133 51263 49190 51309
rect 49236 51263 49293 51309
rect 49339 51263 49396 51309
rect 49442 51263 49499 51309
rect 49545 51263 49602 51309
rect 49852 51263 49865 51309
rect 44799 51222 45323 51235
rect 48765 51234 49865 51263
rect 44799 51176 44812 51222
rect 44858 51176 44925 51222
rect 44971 51176 45038 51222
rect 45084 51176 45151 51222
rect 45197 51176 45264 51222
rect 45310 51176 45323 51222
rect 44799 51147 45323 51176
rect 39008 51085 39326 51114
rect 39008 51039 39021 51085
rect 39067 51039 39144 51085
rect 39190 51039 39267 51085
rect 39313 51039 39326 51085
rect 39008 51026 39326 51039
rect 51789 51222 53789 51235
rect 44799 50998 45323 51027
rect 44799 50952 44812 50998
rect 44858 50952 44925 50998
rect 44971 50952 45038 50998
rect 45084 50952 45151 50998
rect 45197 50952 45264 50998
rect 45310 50952 45323 50998
rect 44799 50923 45323 50952
rect 48765 51085 49865 51114
rect 48765 51039 48778 51085
rect 48824 51039 48881 51085
rect 48927 51039 48984 51085
rect 49030 51039 49087 51085
rect 49133 51039 49190 51085
rect 49236 51039 49293 51085
rect 49339 51039 49396 51085
rect 49442 51039 49499 51085
rect 49545 51039 49602 51085
rect 49852 51039 49865 51085
rect 48765 51010 49865 51039
rect 51789 51176 51802 51222
rect 53776 51176 53789 51222
rect 51789 51147 53789 51176
rect 35260 50861 36360 50890
rect 35260 50815 35273 50861
rect 35523 50815 35580 50861
rect 35626 50815 35683 50861
rect 35729 50815 35786 50861
rect 35832 50815 35889 50861
rect 35935 50815 35992 50861
rect 36038 50815 36095 50861
rect 36141 50815 36198 50861
rect 36244 50815 36301 50861
rect 36347 50815 36360 50861
rect 35260 50802 36360 50815
rect 36841 50861 37501 50890
rect 36841 50815 36854 50861
rect 36900 50815 36971 50861
rect 37017 50815 37088 50861
rect 37134 50815 37206 50861
rect 37252 50815 37324 50861
rect 37370 50815 37442 50861
rect 37488 50815 37501 50861
rect 36841 50802 37501 50815
rect 48765 50861 49865 50890
rect 48765 50815 48778 50861
rect 48824 50815 48881 50861
rect 48927 50815 48984 50861
rect 49030 50815 49087 50861
rect 49133 50815 49190 50861
rect 49236 50815 49293 50861
rect 49339 50815 49396 50861
rect 49442 50815 49499 50861
rect 49545 50815 49602 50861
rect 49852 50815 49865 50861
rect 44799 50774 45323 50803
rect 48765 50802 49865 50815
rect 44799 50728 44812 50774
rect 44858 50728 44925 50774
rect 44971 50728 45038 50774
rect 45084 50728 45151 50774
rect 45197 50728 45264 50774
rect 45310 50728 45323 50774
rect 31336 50550 33336 50579
rect 31336 50504 31349 50550
rect 33323 50504 33336 50550
rect 31336 50475 33336 50504
rect 31336 50326 33336 50355
rect 31336 50280 31349 50326
rect 33323 50280 33336 50326
rect 31336 50251 33336 50280
rect 31336 50102 33336 50131
rect 31336 50056 31349 50102
rect 33323 50056 33336 50102
rect 31336 50027 33336 50056
rect 44799 50699 45323 50728
rect 51789 50998 53789 51027
rect 51789 50952 51802 50998
rect 53776 50952 53789 50998
rect 51789 50923 53789 50952
rect 51789 50774 53789 50803
rect 51789 50728 51802 50774
rect 53776 50728 53789 50774
rect 51789 50699 53789 50728
rect 44799 50550 45323 50579
rect 44799 50504 44812 50550
rect 44858 50504 44925 50550
rect 44971 50504 45038 50550
rect 45084 50504 45151 50550
rect 45197 50504 45264 50550
rect 45310 50504 45323 50550
rect 44799 50475 45323 50504
rect 51789 50550 53789 50579
rect 51789 50504 51802 50550
rect 53776 50504 53789 50550
rect 51789 50475 53789 50504
rect 35260 50239 36360 50252
rect 35260 50193 35273 50239
rect 35523 50193 35580 50239
rect 35626 50193 35683 50239
rect 35729 50193 35786 50239
rect 35832 50193 35889 50239
rect 35935 50193 35992 50239
rect 36038 50193 36095 50239
rect 36141 50193 36198 50239
rect 36244 50193 36301 50239
rect 36347 50193 36360 50239
rect 35260 50164 36360 50193
rect 36841 50239 37501 50252
rect 36841 50193 36854 50239
rect 36900 50193 36971 50239
rect 37017 50193 37088 50239
rect 37134 50193 37206 50239
rect 37252 50193 37324 50239
rect 37370 50193 37442 50239
rect 37488 50193 37501 50239
rect 36841 50164 37501 50193
rect 44799 50326 45323 50355
rect 44799 50280 44812 50326
rect 44858 50280 44925 50326
rect 44971 50280 45038 50326
rect 45084 50280 45151 50326
rect 45197 50280 45264 50326
rect 45310 50280 45323 50326
rect 54750 50550 55849 50583
rect 54750 50504 54793 50550
rect 54839 50504 54956 50550
rect 55002 50504 55118 50550
rect 55164 50504 55279 50550
rect 55325 50504 55439 50550
rect 55485 50504 55599 50550
rect 55645 50504 55760 50550
rect 55806 50504 55849 50550
rect 54750 50471 55849 50504
rect 44799 50251 45323 50280
rect 31336 49878 33336 49907
rect 31336 49832 31349 49878
rect 33323 49832 33336 49878
rect 35260 50015 36360 50044
rect 35260 49969 35273 50015
rect 35523 49969 35580 50015
rect 35626 49969 35683 50015
rect 35729 49969 35786 50015
rect 35832 49969 35889 50015
rect 35935 49969 35992 50015
rect 36038 49969 36095 50015
rect 36141 49969 36198 50015
rect 36244 49969 36301 50015
rect 36347 49969 36360 50015
rect 35260 49940 36360 49969
rect 31336 49819 33336 49832
rect 48765 50239 49865 50252
rect 48765 50193 48778 50239
rect 48824 50193 48881 50239
rect 48927 50193 48984 50239
rect 49030 50193 49087 50239
rect 49133 50193 49190 50239
rect 49236 50193 49293 50239
rect 49339 50193 49396 50239
rect 49442 50193 49499 50239
rect 49545 50193 49602 50239
rect 49852 50193 49865 50239
rect 48765 50164 49865 50193
rect 36841 50015 37501 50044
rect 36841 49969 36854 50015
rect 36900 49969 36971 50015
rect 37017 49969 37088 50015
rect 37134 49969 37206 50015
rect 37252 49969 37324 50015
rect 37370 49969 37442 50015
rect 37488 49969 37501 50015
rect 36841 49940 37501 49969
rect 39008 50015 39326 50028
rect 39008 49969 39021 50015
rect 39067 49969 39144 50015
rect 39190 49969 39267 50015
rect 39313 49969 39326 50015
rect 39008 49940 39326 49969
rect 44799 50102 45323 50131
rect 44799 50056 44812 50102
rect 44858 50056 44925 50102
rect 44971 50056 45038 50102
rect 45084 50056 45151 50102
rect 45197 50056 45264 50102
rect 45310 50056 45323 50102
rect 44799 50027 45323 50056
rect 48765 50015 49865 50044
rect 48765 49969 48778 50015
rect 48824 49969 48881 50015
rect 48927 49969 48984 50015
rect 49030 49969 49087 50015
rect 49133 49969 49190 50015
rect 49236 49969 49293 50015
rect 49339 49969 49396 50015
rect 49442 49969 49499 50015
rect 49545 49969 49602 50015
rect 49852 49969 49865 50015
rect 48765 49940 49865 49969
rect 35260 49791 36360 49820
rect 35260 49745 35273 49791
rect 35523 49745 35580 49791
rect 35626 49745 35683 49791
rect 35729 49745 35786 49791
rect 35832 49745 35889 49791
rect 35935 49745 35992 49791
rect 36038 49745 36095 49791
rect 36141 49745 36198 49791
rect 36244 49745 36301 49791
rect 36347 49745 36360 49791
rect 35260 49732 36360 49745
rect 36841 49791 37501 49820
rect 36841 49745 36854 49791
rect 36900 49745 36971 49791
rect 37017 49745 37088 49791
rect 37134 49745 37206 49791
rect 37252 49745 37324 49791
rect 37370 49745 37442 49791
rect 37488 49745 37501 49791
rect 36841 49732 37501 49745
rect 39008 49791 39326 49820
rect 39008 49745 39021 49791
rect 39067 49745 39144 49791
rect 39190 49745 39267 49791
rect 39313 49745 39326 49791
rect 39008 49732 39326 49745
rect 44799 49878 45323 49907
rect 44799 49832 44812 49878
rect 44858 49832 44925 49878
rect 44971 49832 45038 49878
rect 45084 49832 45151 49878
rect 45197 49832 45264 49878
rect 45310 49832 45323 49878
rect 44799 49819 45323 49832
rect 51789 50326 53789 50355
rect 51789 50280 51802 50326
rect 53776 50280 53789 50326
rect 51789 50251 53789 50280
rect 51789 50102 53789 50131
rect 51789 50056 51802 50102
rect 53776 50056 53789 50102
rect 51789 50027 53789 50056
rect 51789 49878 53789 49907
rect 48765 49791 49865 49820
rect 48765 49745 48778 49791
rect 48824 49745 48881 49791
rect 48927 49745 48984 49791
rect 49030 49745 49087 49791
rect 49133 49745 49190 49791
rect 49236 49745 49293 49791
rect 49339 49745 49396 49791
rect 49442 49745 49499 49791
rect 49545 49745 49602 49791
rect 49852 49745 49865 49791
rect 51789 49832 51802 49878
rect 53776 49832 53789 49878
rect 51789 49819 53789 49832
rect 48765 49732 49865 49745
rect 29274 49650 30373 49683
rect 29274 49604 29317 49650
rect 29363 49604 29478 49650
rect 29524 49604 29638 49650
rect 29684 49604 29798 49650
rect 29844 49604 29959 49650
rect 30005 49604 30121 49650
rect 30167 49604 30284 49650
rect 30330 49604 30373 49650
rect 29274 49571 30373 49604
rect 54750 49650 55849 49683
rect 54750 49604 54793 49650
rect 54839 49604 54956 49650
rect 55002 49604 55118 49650
rect 55164 49604 55279 49650
rect 55325 49604 55439 49650
rect 55485 49604 55599 49650
rect 55645 49604 55760 49650
rect 55806 49604 55849 49650
rect 54750 49571 55849 49604
rect 35260 49509 36360 49522
rect 31336 49422 33336 49435
rect 31336 49376 31349 49422
rect 33323 49376 33336 49422
rect 35260 49463 35273 49509
rect 35523 49463 35580 49509
rect 35626 49463 35683 49509
rect 35729 49463 35786 49509
rect 35832 49463 35889 49509
rect 35935 49463 35992 49509
rect 36038 49463 36095 49509
rect 36141 49463 36198 49509
rect 36244 49463 36301 49509
rect 36347 49463 36360 49509
rect 35260 49434 36360 49463
rect 36841 49509 37501 49522
rect 36841 49463 36854 49509
rect 36900 49463 36971 49509
rect 37017 49463 37088 49509
rect 37134 49463 37206 49509
rect 37252 49463 37324 49509
rect 37370 49463 37442 49509
rect 37488 49463 37501 49509
rect 36841 49434 37501 49463
rect 39008 49509 39326 49522
rect 39008 49463 39021 49509
rect 39067 49463 39144 49509
rect 39190 49463 39267 49509
rect 39313 49463 39326 49509
rect 39008 49434 39326 49463
rect 48765 49509 49865 49522
rect 31336 49347 33336 49376
rect 31336 49198 33336 49227
rect 31336 49152 31349 49198
rect 33323 49152 33336 49198
rect 31336 49123 33336 49152
rect 31336 48974 33336 49003
rect 31336 48928 31349 48974
rect 33323 48928 33336 48974
rect 31336 48899 33336 48928
rect 29274 48750 30373 48783
rect 29274 48704 29317 48750
rect 29363 48704 29478 48750
rect 29524 48704 29638 48750
rect 29684 48704 29798 48750
rect 29844 48704 29959 48750
rect 30005 48704 30121 48750
rect 30167 48704 30284 48750
rect 30330 48704 30373 48750
rect 29274 48671 30373 48704
rect 35260 49285 36360 49314
rect 35260 49239 35273 49285
rect 35523 49239 35580 49285
rect 35626 49239 35683 49285
rect 35729 49239 35786 49285
rect 35832 49239 35889 49285
rect 35935 49239 35992 49285
rect 36038 49239 36095 49285
rect 36141 49239 36198 49285
rect 36244 49239 36301 49285
rect 36347 49239 36360 49285
rect 35260 49210 36360 49239
rect 36841 49285 37501 49314
rect 36841 49239 36854 49285
rect 36900 49239 36971 49285
rect 37017 49239 37088 49285
rect 37134 49239 37206 49285
rect 37252 49239 37324 49285
rect 37370 49239 37442 49285
rect 37488 49239 37501 49285
rect 36841 49210 37501 49239
rect 48765 49463 48778 49509
rect 48824 49463 48881 49509
rect 48927 49463 48984 49509
rect 49030 49463 49087 49509
rect 49133 49463 49190 49509
rect 49236 49463 49293 49509
rect 49339 49463 49396 49509
rect 49442 49463 49499 49509
rect 49545 49463 49602 49509
rect 49852 49463 49865 49509
rect 44799 49422 45323 49435
rect 48765 49434 49865 49463
rect 44799 49376 44812 49422
rect 44858 49376 44925 49422
rect 44971 49376 45038 49422
rect 45084 49376 45151 49422
rect 45197 49376 45264 49422
rect 45310 49376 45323 49422
rect 44799 49347 45323 49376
rect 39008 49285 39326 49314
rect 39008 49239 39021 49285
rect 39067 49239 39144 49285
rect 39190 49239 39267 49285
rect 39313 49239 39326 49285
rect 39008 49226 39326 49239
rect 51789 49422 53789 49435
rect 44799 49198 45323 49227
rect 44799 49152 44812 49198
rect 44858 49152 44925 49198
rect 44971 49152 45038 49198
rect 45084 49152 45151 49198
rect 45197 49152 45264 49198
rect 45310 49152 45323 49198
rect 44799 49123 45323 49152
rect 48765 49285 49865 49314
rect 48765 49239 48778 49285
rect 48824 49239 48881 49285
rect 48927 49239 48984 49285
rect 49030 49239 49087 49285
rect 49133 49239 49190 49285
rect 49236 49239 49293 49285
rect 49339 49239 49396 49285
rect 49442 49239 49499 49285
rect 49545 49239 49602 49285
rect 49852 49239 49865 49285
rect 48765 49210 49865 49239
rect 51789 49376 51802 49422
rect 53776 49376 53789 49422
rect 51789 49347 53789 49376
rect 35260 49061 36360 49090
rect 35260 49015 35273 49061
rect 35523 49015 35580 49061
rect 35626 49015 35683 49061
rect 35729 49015 35786 49061
rect 35832 49015 35889 49061
rect 35935 49015 35992 49061
rect 36038 49015 36095 49061
rect 36141 49015 36198 49061
rect 36244 49015 36301 49061
rect 36347 49015 36360 49061
rect 35260 49002 36360 49015
rect 36841 49061 37501 49090
rect 36841 49015 36854 49061
rect 36900 49015 36971 49061
rect 37017 49015 37088 49061
rect 37134 49015 37206 49061
rect 37252 49015 37324 49061
rect 37370 49015 37442 49061
rect 37488 49015 37501 49061
rect 36841 49002 37501 49015
rect 48765 49061 49865 49090
rect 48765 49015 48778 49061
rect 48824 49015 48881 49061
rect 48927 49015 48984 49061
rect 49030 49015 49087 49061
rect 49133 49015 49190 49061
rect 49236 49015 49293 49061
rect 49339 49015 49396 49061
rect 49442 49015 49499 49061
rect 49545 49015 49602 49061
rect 49852 49015 49865 49061
rect 44799 48974 45323 49003
rect 48765 49002 49865 49015
rect 44799 48928 44812 48974
rect 44858 48928 44925 48974
rect 44971 48928 45038 48974
rect 45084 48928 45151 48974
rect 45197 48928 45264 48974
rect 45310 48928 45323 48974
rect 31336 48750 33336 48779
rect 31336 48704 31349 48750
rect 33323 48704 33336 48750
rect 31336 48675 33336 48704
rect 31336 48526 33336 48555
rect 31336 48480 31349 48526
rect 33323 48480 33336 48526
rect 31336 48451 33336 48480
rect 31336 48302 33336 48331
rect 31336 48256 31349 48302
rect 33323 48256 33336 48302
rect 31336 48227 33336 48256
rect 44799 48899 45323 48928
rect 51789 49198 53789 49227
rect 51789 49152 51802 49198
rect 53776 49152 53789 49198
rect 51789 49123 53789 49152
rect 51789 48974 53789 49003
rect 51789 48928 51802 48974
rect 53776 48928 53789 48974
rect 51789 48899 53789 48928
rect 44799 48750 45323 48779
rect 44799 48704 44812 48750
rect 44858 48704 44925 48750
rect 44971 48704 45038 48750
rect 45084 48704 45151 48750
rect 45197 48704 45264 48750
rect 45310 48704 45323 48750
rect 44799 48675 45323 48704
rect 51789 48750 53789 48779
rect 51789 48704 51802 48750
rect 53776 48704 53789 48750
rect 51789 48675 53789 48704
rect 35260 48439 36360 48452
rect 35260 48393 35273 48439
rect 35523 48393 35580 48439
rect 35626 48393 35683 48439
rect 35729 48393 35786 48439
rect 35832 48393 35889 48439
rect 35935 48393 35992 48439
rect 36038 48393 36095 48439
rect 36141 48393 36198 48439
rect 36244 48393 36301 48439
rect 36347 48393 36360 48439
rect 35260 48364 36360 48393
rect 36841 48439 37501 48452
rect 36841 48393 36854 48439
rect 36900 48393 36971 48439
rect 37017 48393 37088 48439
rect 37134 48393 37206 48439
rect 37252 48393 37324 48439
rect 37370 48393 37442 48439
rect 37488 48393 37501 48439
rect 36841 48364 37501 48393
rect 44799 48526 45323 48555
rect 44799 48480 44812 48526
rect 44858 48480 44925 48526
rect 44971 48480 45038 48526
rect 45084 48480 45151 48526
rect 45197 48480 45264 48526
rect 45310 48480 45323 48526
rect 54750 48750 55849 48783
rect 54750 48704 54793 48750
rect 54839 48704 54956 48750
rect 55002 48704 55118 48750
rect 55164 48704 55279 48750
rect 55325 48704 55439 48750
rect 55485 48704 55599 48750
rect 55645 48704 55760 48750
rect 55806 48704 55849 48750
rect 54750 48671 55849 48704
rect 44799 48451 45323 48480
rect 31336 48078 33336 48107
rect 31336 48032 31349 48078
rect 33323 48032 33336 48078
rect 35260 48215 36360 48244
rect 35260 48169 35273 48215
rect 35523 48169 35580 48215
rect 35626 48169 35683 48215
rect 35729 48169 35786 48215
rect 35832 48169 35889 48215
rect 35935 48169 35992 48215
rect 36038 48169 36095 48215
rect 36141 48169 36198 48215
rect 36244 48169 36301 48215
rect 36347 48169 36360 48215
rect 35260 48140 36360 48169
rect 31336 48019 33336 48032
rect 48765 48439 49865 48452
rect 48765 48393 48778 48439
rect 48824 48393 48881 48439
rect 48927 48393 48984 48439
rect 49030 48393 49087 48439
rect 49133 48393 49190 48439
rect 49236 48393 49293 48439
rect 49339 48393 49396 48439
rect 49442 48393 49499 48439
rect 49545 48393 49602 48439
rect 49852 48393 49865 48439
rect 48765 48364 49865 48393
rect 36841 48215 37501 48244
rect 36841 48169 36854 48215
rect 36900 48169 36971 48215
rect 37017 48169 37088 48215
rect 37134 48169 37206 48215
rect 37252 48169 37324 48215
rect 37370 48169 37442 48215
rect 37488 48169 37501 48215
rect 36841 48140 37501 48169
rect 39008 48215 39326 48228
rect 39008 48169 39021 48215
rect 39067 48169 39144 48215
rect 39190 48169 39267 48215
rect 39313 48169 39326 48215
rect 39008 48140 39326 48169
rect 44799 48302 45323 48331
rect 44799 48256 44812 48302
rect 44858 48256 44925 48302
rect 44971 48256 45038 48302
rect 45084 48256 45151 48302
rect 45197 48256 45264 48302
rect 45310 48256 45323 48302
rect 44799 48227 45323 48256
rect 48765 48215 49865 48244
rect 48765 48169 48778 48215
rect 48824 48169 48881 48215
rect 48927 48169 48984 48215
rect 49030 48169 49087 48215
rect 49133 48169 49190 48215
rect 49236 48169 49293 48215
rect 49339 48169 49396 48215
rect 49442 48169 49499 48215
rect 49545 48169 49602 48215
rect 49852 48169 49865 48215
rect 48765 48140 49865 48169
rect 35260 47991 36360 48020
rect 35260 47945 35273 47991
rect 35523 47945 35580 47991
rect 35626 47945 35683 47991
rect 35729 47945 35786 47991
rect 35832 47945 35889 47991
rect 35935 47945 35992 47991
rect 36038 47945 36095 47991
rect 36141 47945 36198 47991
rect 36244 47945 36301 47991
rect 36347 47945 36360 47991
rect 35260 47932 36360 47945
rect 36841 47991 37501 48020
rect 36841 47945 36854 47991
rect 36900 47945 36971 47991
rect 37017 47945 37088 47991
rect 37134 47945 37206 47991
rect 37252 47945 37324 47991
rect 37370 47945 37442 47991
rect 37488 47945 37501 47991
rect 36841 47932 37501 47945
rect 39008 47991 39326 48020
rect 39008 47945 39021 47991
rect 39067 47945 39144 47991
rect 39190 47945 39267 47991
rect 39313 47945 39326 47991
rect 39008 47932 39326 47945
rect 44799 48078 45323 48107
rect 44799 48032 44812 48078
rect 44858 48032 44925 48078
rect 44971 48032 45038 48078
rect 45084 48032 45151 48078
rect 45197 48032 45264 48078
rect 45310 48032 45323 48078
rect 44799 48019 45323 48032
rect 51789 48526 53789 48555
rect 51789 48480 51802 48526
rect 53776 48480 53789 48526
rect 51789 48451 53789 48480
rect 51789 48302 53789 48331
rect 51789 48256 51802 48302
rect 53776 48256 53789 48302
rect 51789 48227 53789 48256
rect 51789 48078 53789 48107
rect 48765 47991 49865 48020
rect 48765 47945 48778 47991
rect 48824 47945 48881 47991
rect 48927 47945 48984 47991
rect 49030 47945 49087 47991
rect 49133 47945 49190 47991
rect 49236 47945 49293 47991
rect 49339 47945 49396 47991
rect 49442 47945 49499 47991
rect 49545 47945 49602 47991
rect 49852 47945 49865 47991
rect 51789 48032 51802 48078
rect 53776 48032 53789 48078
rect 51789 48019 53789 48032
rect 48765 47932 49865 47945
rect 29274 47850 30373 47883
rect 29274 47804 29317 47850
rect 29363 47804 29478 47850
rect 29524 47804 29638 47850
rect 29684 47804 29798 47850
rect 29844 47804 29959 47850
rect 30005 47804 30121 47850
rect 30167 47804 30284 47850
rect 30330 47804 30373 47850
rect 29274 47771 30373 47804
rect 54750 47850 55849 47883
rect 54750 47804 54793 47850
rect 54839 47804 54956 47850
rect 55002 47804 55118 47850
rect 55164 47804 55279 47850
rect 55325 47804 55439 47850
rect 55485 47804 55599 47850
rect 55645 47804 55760 47850
rect 55806 47804 55849 47850
rect 54750 47771 55849 47804
rect 35260 47709 36360 47722
rect 31336 47622 33336 47635
rect 31336 47576 31349 47622
rect 33323 47576 33336 47622
rect 35260 47663 35273 47709
rect 35523 47663 35580 47709
rect 35626 47663 35683 47709
rect 35729 47663 35786 47709
rect 35832 47663 35889 47709
rect 35935 47663 35992 47709
rect 36038 47663 36095 47709
rect 36141 47663 36198 47709
rect 36244 47663 36301 47709
rect 36347 47663 36360 47709
rect 35260 47634 36360 47663
rect 36841 47709 37501 47722
rect 36841 47663 36854 47709
rect 36900 47663 36971 47709
rect 37017 47663 37088 47709
rect 37134 47663 37206 47709
rect 37252 47663 37324 47709
rect 37370 47663 37442 47709
rect 37488 47663 37501 47709
rect 36841 47634 37501 47663
rect 39008 47709 39326 47722
rect 39008 47663 39021 47709
rect 39067 47663 39144 47709
rect 39190 47663 39267 47709
rect 39313 47663 39326 47709
rect 39008 47634 39326 47663
rect 48765 47709 49865 47722
rect 31336 47547 33336 47576
rect 31336 47398 33336 47427
rect 31336 47352 31349 47398
rect 33323 47352 33336 47398
rect 31336 47323 33336 47352
rect 31336 47174 33336 47203
rect 31336 47128 31349 47174
rect 33323 47128 33336 47174
rect 31336 47099 33336 47128
rect 29274 46950 30373 46983
rect 29274 46904 29317 46950
rect 29363 46904 29478 46950
rect 29524 46904 29638 46950
rect 29684 46904 29798 46950
rect 29844 46904 29959 46950
rect 30005 46904 30121 46950
rect 30167 46904 30284 46950
rect 30330 46904 30373 46950
rect 29274 46871 30373 46904
rect 35260 47485 36360 47514
rect 35260 47439 35273 47485
rect 35523 47439 35580 47485
rect 35626 47439 35683 47485
rect 35729 47439 35786 47485
rect 35832 47439 35889 47485
rect 35935 47439 35992 47485
rect 36038 47439 36095 47485
rect 36141 47439 36198 47485
rect 36244 47439 36301 47485
rect 36347 47439 36360 47485
rect 35260 47410 36360 47439
rect 36841 47485 37501 47514
rect 36841 47439 36854 47485
rect 36900 47439 36971 47485
rect 37017 47439 37088 47485
rect 37134 47439 37206 47485
rect 37252 47439 37324 47485
rect 37370 47439 37442 47485
rect 37488 47439 37501 47485
rect 36841 47410 37501 47439
rect 48765 47663 48778 47709
rect 48824 47663 48881 47709
rect 48927 47663 48984 47709
rect 49030 47663 49087 47709
rect 49133 47663 49190 47709
rect 49236 47663 49293 47709
rect 49339 47663 49396 47709
rect 49442 47663 49499 47709
rect 49545 47663 49602 47709
rect 49852 47663 49865 47709
rect 44799 47622 45323 47635
rect 48765 47634 49865 47663
rect 44799 47576 44812 47622
rect 44858 47576 44925 47622
rect 44971 47576 45038 47622
rect 45084 47576 45151 47622
rect 45197 47576 45264 47622
rect 45310 47576 45323 47622
rect 44799 47547 45323 47576
rect 39008 47485 39326 47514
rect 39008 47439 39021 47485
rect 39067 47439 39144 47485
rect 39190 47439 39267 47485
rect 39313 47439 39326 47485
rect 39008 47426 39326 47439
rect 51789 47622 53789 47635
rect 44799 47398 45323 47427
rect 44799 47352 44812 47398
rect 44858 47352 44925 47398
rect 44971 47352 45038 47398
rect 45084 47352 45151 47398
rect 45197 47352 45264 47398
rect 45310 47352 45323 47398
rect 44799 47323 45323 47352
rect 48765 47485 49865 47514
rect 48765 47439 48778 47485
rect 48824 47439 48881 47485
rect 48927 47439 48984 47485
rect 49030 47439 49087 47485
rect 49133 47439 49190 47485
rect 49236 47439 49293 47485
rect 49339 47439 49396 47485
rect 49442 47439 49499 47485
rect 49545 47439 49602 47485
rect 49852 47439 49865 47485
rect 48765 47410 49865 47439
rect 51789 47576 51802 47622
rect 53776 47576 53789 47622
rect 51789 47547 53789 47576
rect 35260 47261 36360 47290
rect 35260 47215 35273 47261
rect 35523 47215 35580 47261
rect 35626 47215 35683 47261
rect 35729 47215 35786 47261
rect 35832 47215 35889 47261
rect 35935 47215 35992 47261
rect 36038 47215 36095 47261
rect 36141 47215 36198 47261
rect 36244 47215 36301 47261
rect 36347 47215 36360 47261
rect 35260 47202 36360 47215
rect 36841 47261 37501 47290
rect 36841 47215 36854 47261
rect 36900 47215 36971 47261
rect 37017 47215 37088 47261
rect 37134 47215 37206 47261
rect 37252 47215 37324 47261
rect 37370 47215 37442 47261
rect 37488 47215 37501 47261
rect 36841 47202 37501 47215
rect 48765 47261 49865 47290
rect 48765 47215 48778 47261
rect 48824 47215 48881 47261
rect 48927 47215 48984 47261
rect 49030 47215 49087 47261
rect 49133 47215 49190 47261
rect 49236 47215 49293 47261
rect 49339 47215 49396 47261
rect 49442 47215 49499 47261
rect 49545 47215 49602 47261
rect 49852 47215 49865 47261
rect 44799 47174 45323 47203
rect 48765 47202 49865 47215
rect 44799 47128 44812 47174
rect 44858 47128 44925 47174
rect 44971 47128 45038 47174
rect 45084 47128 45151 47174
rect 45197 47128 45264 47174
rect 45310 47128 45323 47174
rect 31336 46950 33336 46979
rect 31336 46904 31349 46950
rect 33323 46904 33336 46950
rect 31336 46875 33336 46904
rect 31336 46726 33336 46755
rect 31336 46680 31349 46726
rect 33323 46680 33336 46726
rect 31336 46651 33336 46680
rect 31336 46502 33336 46531
rect 31336 46456 31349 46502
rect 33323 46456 33336 46502
rect 31336 46427 33336 46456
rect 44799 47099 45323 47128
rect 51789 47398 53789 47427
rect 51789 47352 51802 47398
rect 53776 47352 53789 47398
rect 51789 47323 53789 47352
rect 51789 47174 53789 47203
rect 51789 47128 51802 47174
rect 53776 47128 53789 47174
rect 51789 47099 53789 47128
rect 44799 46950 45323 46979
rect 44799 46904 44812 46950
rect 44858 46904 44925 46950
rect 44971 46904 45038 46950
rect 45084 46904 45151 46950
rect 45197 46904 45264 46950
rect 45310 46904 45323 46950
rect 44799 46875 45323 46904
rect 51789 46950 53789 46979
rect 51789 46904 51802 46950
rect 53776 46904 53789 46950
rect 51789 46875 53789 46904
rect 35260 46639 36360 46652
rect 35260 46593 35273 46639
rect 35523 46593 35580 46639
rect 35626 46593 35683 46639
rect 35729 46593 35786 46639
rect 35832 46593 35889 46639
rect 35935 46593 35992 46639
rect 36038 46593 36095 46639
rect 36141 46593 36198 46639
rect 36244 46593 36301 46639
rect 36347 46593 36360 46639
rect 35260 46564 36360 46593
rect 36841 46639 37501 46652
rect 36841 46593 36854 46639
rect 36900 46593 36971 46639
rect 37017 46593 37088 46639
rect 37134 46593 37206 46639
rect 37252 46593 37324 46639
rect 37370 46593 37442 46639
rect 37488 46593 37501 46639
rect 36841 46564 37501 46593
rect 44799 46726 45323 46755
rect 44799 46680 44812 46726
rect 44858 46680 44925 46726
rect 44971 46680 45038 46726
rect 45084 46680 45151 46726
rect 45197 46680 45264 46726
rect 45310 46680 45323 46726
rect 54750 46950 55849 46983
rect 54750 46904 54793 46950
rect 54839 46904 54956 46950
rect 55002 46904 55118 46950
rect 55164 46904 55279 46950
rect 55325 46904 55439 46950
rect 55485 46904 55599 46950
rect 55645 46904 55760 46950
rect 55806 46904 55849 46950
rect 54750 46871 55849 46904
rect 44799 46651 45323 46680
rect 31336 46278 33336 46307
rect 31336 46232 31349 46278
rect 33323 46232 33336 46278
rect 35260 46415 36360 46444
rect 35260 46369 35273 46415
rect 35523 46369 35580 46415
rect 35626 46369 35683 46415
rect 35729 46369 35786 46415
rect 35832 46369 35889 46415
rect 35935 46369 35992 46415
rect 36038 46369 36095 46415
rect 36141 46369 36198 46415
rect 36244 46369 36301 46415
rect 36347 46369 36360 46415
rect 35260 46340 36360 46369
rect 31336 46219 33336 46232
rect 48765 46639 49865 46652
rect 48765 46593 48778 46639
rect 48824 46593 48881 46639
rect 48927 46593 48984 46639
rect 49030 46593 49087 46639
rect 49133 46593 49190 46639
rect 49236 46593 49293 46639
rect 49339 46593 49396 46639
rect 49442 46593 49499 46639
rect 49545 46593 49602 46639
rect 49852 46593 49865 46639
rect 48765 46564 49865 46593
rect 36841 46415 37501 46444
rect 36841 46369 36854 46415
rect 36900 46369 36971 46415
rect 37017 46369 37088 46415
rect 37134 46369 37206 46415
rect 37252 46369 37324 46415
rect 37370 46369 37442 46415
rect 37488 46369 37501 46415
rect 36841 46340 37501 46369
rect 39008 46415 39326 46428
rect 39008 46369 39021 46415
rect 39067 46369 39144 46415
rect 39190 46369 39267 46415
rect 39313 46369 39326 46415
rect 39008 46340 39326 46369
rect 44799 46502 45323 46531
rect 44799 46456 44812 46502
rect 44858 46456 44925 46502
rect 44971 46456 45038 46502
rect 45084 46456 45151 46502
rect 45197 46456 45264 46502
rect 45310 46456 45323 46502
rect 44799 46427 45323 46456
rect 48765 46415 49865 46444
rect 48765 46369 48778 46415
rect 48824 46369 48881 46415
rect 48927 46369 48984 46415
rect 49030 46369 49087 46415
rect 49133 46369 49190 46415
rect 49236 46369 49293 46415
rect 49339 46369 49396 46415
rect 49442 46369 49499 46415
rect 49545 46369 49602 46415
rect 49852 46369 49865 46415
rect 48765 46340 49865 46369
rect 35260 46191 36360 46220
rect 35260 46145 35273 46191
rect 35523 46145 35580 46191
rect 35626 46145 35683 46191
rect 35729 46145 35786 46191
rect 35832 46145 35889 46191
rect 35935 46145 35992 46191
rect 36038 46145 36095 46191
rect 36141 46145 36198 46191
rect 36244 46145 36301 46191
rect 36347 46145 36360 46191
rect 35260 46132 36360 46145
rect 36841 46191 37501 46220
rect 36841 46145 36854 46191
rect 36900 46145 36971 46191
rect 37017 46145 37088 46191
rect 37134 46145 37206 46191
rect 37252 46145 37324 46191
rect 37370 46145 37442 46191
rect 37488 46145 37501 46191
rect 36841 46132 37501 46145
rect 39008 46191 39326 46220
rect 39008 46145 39021 46191
rect 39067 46145 39144 46191
rect 39190 46145 39267 46191
rect 39313 46145 39326 46191
rect 39008 46132 39326 46145
rect 44799 46278 45323 46307
rect 44799 46232 44812 46278
rect 44858 46232 44925 46278
rect 44971 46232 45038 46278
rect 45084 46232 45151 46278
rect 45197 46232 45264 46278
rect 45310 46232 45323 46278
rect 44799 46219 45323 46232
rect 51789 46726 53789 46755
rect 51789 46680 51802 46726
rect 53776 46680 53789 46726
rect 51789 46651 53789 46680
rect 51789 46502 53789 46531
rect 51789 46456 51802 46502
rect 53776 46456 53789 46502
rect 51789 46427 53789 46456
rect 51789 46278 53789 46307
rect 48765 46191 49865 46220
rect 48765 46145 48778 46191
rect 48824 46145 48881 46191
rect 48927 46145 48984 46191
rect 49030 46145 49087 46191
rect 49133 46145 49190 46191
rect 49236 46145 49293 46191
rect 49339 46145 49396 46191
rect 49442 46145 49499 46191
rect 49545 46145 49602 46191
rect 49852 46145 49865 46191
rect 51789 46232 51802 46278
rect 53776 46232 53789 46278
rect 51789 46219 53789 46232
rect 48765 46132 49865 46145
rect 29274 46050 30373 46083
rect 29274 46004 29317 46050
rect 29363 46004 29478 46050
rect 29524 46004 29638 46050
rect 29684 46004 29798 46050
rect 29844 46004 29959 46050
rect 30005 46004 30121 46050
rect 30167 46004 30284 46050
rect 30330 46004 30373 46050
rect 29274 45971 30373 46004
rect 54750 46050 55849 46083
rect 54750 46004 54793 46050
rect 54839 46004 54956 46050
rect 55002 46004 55118 46050
rect 55164 46004 55279 46050
rect 55325 46004 55439 46050
rect 55485 46004 55599 46050
rect 55645 46004 55760 46050
rect 55806 46004 55849 46050
rect 54750 45971 55849 46004
rect 35260 45909 36360 45922
rect 31336 45822 33336 45835
rect 31336 45776 31349 45822
rect 33323 45776 33336 45822
rect 35260 45863 35273 45909
rect 35523 45863 35580 45909
rect 35626 45863 35683 45909
rect 35729 45863 35786 45909
rect 35832 45863 35889 45909
rect 35935 45863 35992 45909
rect 36038 45863 36095 45909
rect 36141 45863 36198 45909
rect 36244 45863 36301 45909
rect 36347 45863 36360 45909
rect 35260 45834 36360 45863
rect 36841 45909 37501 45922
rect 36841 45863 36854 45909
rect 36900 45863 36971 45909
rect 37017 45863 37088 45909
rect 37134 45863 37206 45909
rect 37252 45863 37324 45909
rect 37370 45863 37442 45909
rect 37488 45863 37501 45909
rect 36841 45834 37501 45863
rect 39008 45909 39326 45922
rect 39008 45863 39021 45909
rect 39067 45863 39144 45909
rect 39190 45863 39267 45909
rect 39313 45863 39326 45909
rect 39008 45834 39326 45863
rect 48765 45909 49865 45922
rect 31336 45747 33336 45776
rect 31336 45598 33336 45627
rect 31336 45552 31349 45598
rect 33323 45552 33336 45598
rect 31336 45523 33336 45552
rect 31336 45374 33336 45403
rect 31336 45328 31349 45374
rect 33323 45328 33336 45374
rect 31336 45299 33336 45328
rect 29274 45150 30373 45183
rect 29274 45104 29317 45150
rect 29363 45104 29478 45150
rect 29524 45104 29638 45150
rect 29684 45104 29798 45150
rect 29844 45104 29959 45150
rect 30005 45104 30121 45150
rect 30167 45104 30284 45150
rect 30330 45104 30373 45150
rect 29274 45071 30373 45104
rect 35260 45685 36360 45714
rect 35260 45639 35273 45685
rect 35523 45639 35580 45685
rect 35626 45639 35683 45685
rect 35729 45639 35786 45685
rect 35832 45639 35889 45685
rect 35935 45639 35992 45685
rect 36038 45639 36095 45685
rect 36141 45639 36198 45685
rect 36244 45639 36301 45685
rect 36347 45639 36360 45685
rect 35260 45610 36360 45639
rect 36841 45685 37501 45714
rect 36841 45639 36854 45685
rect 36900 45639 36971 45685
rect 37017 45639 37088 45685
rect 37134 45639 37206 45685
rect 37252 45639 37324 45685
rect 37370 45639 37442 45685
rect 37488 45639 37501 45685
rect 36841 45610 37501 45639
rect 48765 45863 48778 45909
rect 48824 45863 48881 45909
rect 48927 45863 48984 45909
rect 49030 45863 49087 45909
rect 49133 45863 49190 45909
rect 49236 45863 49293 45909
rect 49339 45863 49396 45909
rect 49442 45863 49499 45909
rect 49545 45863 49602 45909
rect 49852 45863 49865 45909
rect 44799 45822 45323 45835
rect 48765 45834 49865 45863
rect 44799 45776 44812 45822
rect 44858 45776 44925 45822
rect 44971 45776 45038 45822
rect 45084 45776 45151 45822
rect 45197 45776 45264 45822
rect 45310 45776 45323 45822
rect 44799 45747 45323 45776
rect 39008 45685 39326 45714
rect 39008 45639 39021 45685
rect 39067 45639 39144 45685
rect 39190 45639 39267 45685
rect 39313 45639 39326 45685
rect 39008 45626 39326 45639
rect 51789 45822 53789 45835
rect 44799 45598 45323 45627
rect 44799 45552 44812 45598
rect 44858 45552 44925 45598
rect 44971 45552 45038 45598
rect 45084 45552 45151 45598
rect 45197 45552 45264 45598
rect 45310 45552 45323 45598
rect 44799 45523 45323 45552
rect 48765 45685 49865 45714
rect 48765 45639 48778 45685
rect 48824 45639 48881 45685
rect 48927 45639 48984 45685
rect 49030 45639 49087 45685
rect 49133 45639 49190 45685
rect 49236 45639 49293 45685
rect 49339 45639 49396 45685
rect 49442 45639 49499 45685
rect 49545 45639 49602 45685
rect 49852 45639 49865 45685
rect 48765 45610 49865 45639
rect 51789 45776 51802 45822
rect 53776 45776 53789 45822
rect 51789 45747 53789 45776
rect 35260 45461 36360 45490
rect 35260 45415 35273 45461
rect 35523 45415 35580 45461
rect 35626 45415 35683 45461
rect 35729 45415 35786 45461
rect 35832 45415 35889 45461
rect 35935 45415 35992 45461
rect 36038 45415 36095 45461
rect 36141 45415 36198 45461
rect 36244 45415 36301 45461
rect 36347 45415 36360 45461
rect 35260 45402 36360 45415
rect 36841 45461 37501 45490
rect 36841 45415 36854 45461
rect 36900 45415 36971 45461
rect 37017 45415 37088 45461
rect 37134 45415 37206 45461
rect 37252 45415 37324 45461
rect 37370 45415 37442 45461
rect 37488 45415 37501 45461
rect 36841 45402 37501 45415
rect 48765 45461 49865 45490
rect 48765 45415 48778 45461
rect 48824 45415 48881 45461
rect 48927 45415 48984 45461
rect 49030 45415 49087 45461
rect 49133 45415 49190 45461
rect 49236 45415 49293 45461
rect 49339 45415 49396 45461
rect 49442 45415 49499 45461
rect 49545 45415 49602 45461
rect 49852 45415 49865 45461
rect 44799 45374 45323 45403
rect 48765 45402 49865 45415
rect 44799 45328 44812 45374
rect 44858 45328 44925 45374
rect 44971 45328 45038 45374
rect 45084 45328 45151 45374
rect 45197 45328 45264 45374
rect 45310 45328 45323 45374
rect 31336 45150 33336 45179
rect 31336 45104 31349 45150
rect 33323 45104 33336 45150
rect 31336 45075 33336 45104
rect 31336 44926 33336 44955
rect 31336 44880 31349 44926
rect 33323 44880 33336 44926
rect 31336 44851 33336 44880
rect 31336 44702 33336 44731
rect 31336 44656 31349 44702
rect 33323 44656 33336 44702
rect 31336 44627 33336 44656
rect 44799 45299 45323 45328
rect 51789 45598 53789 45627
rect 51789 45552 51802 45598
rect 53776 45552 53789 45598
rect 51789 45523 53789 45552
rect 51789 45374 53789 45403
rect 51789 45328 51802 45374
rect 53776 45328 53789 45374
rect 51789 45299 53789 45328
rect 44799 45150 45323 45179
rect 44799 45104 44812 45150
rect 44858 45104 44925 45150
rect 44971 45104 45038 45150
rect 45084 45104 45151 45150
rect 45197 45104 45264 45150
rect 45310 45104 45323 45150
rect 44799 45075 45323 45104
rect 51789 45150 53789 45179
rect 51789 45104 51802 45150
rect 53776 45104 53789 45150
rect 51789 45075 53789 45104
rect 35260 44839 36360 44852
rect 35260 44793 35273 44839
rect 35523 44793 35580 44839
rect 35626 44793 35683 44839
rect 35729 44793 35786 44839
rect 35832 44793 35889 44839
rect 35935 44793 35992 44839
rect 36038 44793 36095 44839
rect 36141 44793 36198 44839
rect 36244 44793 36301 44839
rect 36347 44793 36360 44839
rect 35260 44764 36360 44793
rect 36841 44839 37501 44852
rect 36841 44793 36854 44839
rect 36900 44793 36971 44839
rect 37017 44793 37088 44839
rect 37134 44793 37206 44839
rect 37252 44793 37324 44839
rect 37370 44793 37442 44839
rect 37488 44793 37501 44839
rect 36841 44764 37501 44793
rect 44799 44926 45323 44955
rect 44799 44880 44812 44926
rect 44858 44880 44925 44926
rect 44971 44880 45038 44926
rect 45084 44880 45151 44926
rect 45197 44880 45264 44926
rect 45310 44880 45323 44926
rect 54750 45150 55849 45183
rect 54750 45104 54793 45150
rect 54839 45104 54956 45150
rect 55002 45104 55118 45150
rect 55164 45104 55279 45150
rect 55325 45104 55439 45150
rect 55485 45104 55599 45150
rect 55645 45104 55760 45150
rect 55806 45104 55849 45150
rect 54750 45071 55849 45104
rect 44799 44851 45323 44880
rect 31336 44478 33336 44507
rect 31336 44432 31349 44478
rect 33323 44432 33336 44478
rect 35260 44615 36360 44644
rect 35260 44569 35273 44615
rect 35523 44569 35580 44615
rect 35626 44569 35683 44615
rect 35729 44569 35786 44615
rect 35832 44569 35889 44615
rect 35935 44569 35992 44615
rect 36038 44569 36095 44615
rect 36141 44569 36198 44615
rect 36244 44569 36301 44615
rect 36347 44569 36360 44615
rect 35260 44540 36360 44569
rect 31336 44419 33336 44432
rect 48765 44839 49865 44852
rect 48765 44793 48778 44839
rect 48824 44793 48881 44839
rect 48927 44793 48984 44839
rect 49030 44793 49087 44839
rect 49133 44793 49190 44839
rect 49236 44793 49293 44839
rect 49339 44793 49396 44839
rect 49442 44793 49499 44839
rect 49545 44793 49602 44839
rect 49852 44793 49865 44839
rect 48765 44764 49865 44793
rect 36841 44615 37501 44644
rect 36841 44569 36854 44615
rect 36900 44569 36971 44615
rect 37017 44569 37088 44615
rect 37134 44569 37206 44615
rect 37252 44569 37324 44615
rect 37370 44569 37442 44615
rect 37488 44569 37501 44615
rect 36841 44540 37501 44569
rect 39008 44615 39326 44628
rect 39008 44569 39021 44615
rect 39067 44569 39144 44615
rect 39190 44569 39267 44615
rect 39313 44569 39326 44615
rect 39008 44540 39326 44569
rect 44799 44702 45323 44731
rect 44799 44656 44812 44702
rect 44858 44656 44925 44702
rect 44971 44656 45038 44702
rect 45084 44656 45151 44702
rect 45197 44656 45264 44702
rect 45310 44656 45323 44702
rect 44799 44627 45323 44656
rect 48765 44615 49865 44644
rect 48765 44569 48778 44615
rect 48824 44569 48881 44615
rect 48927 44569 48984 44615
rect 49030 44569 49087 44615
rect 49133 44569 49190 44615
rect 49236 44569 49293 44615
rect 49339 44569 49396 44615
rect 49442 44569 49499 44615
rect 49545 44569 49602 44615
rect 49852 44569 49865 44615
rect 48765 44540 49865 44569
rect 35260 44391 36360 44420
rect 35260 44345 35273 44391
rect 35523 44345 35580 44391
rect 35626 44345 35683 44391
rect 35729 44345 35786 44391
rect 35832 44345 35889 44391
rect 35935 44345 35992 44391
rect 36038 44345 36095 44391
rect 36141 44345 36198 44391
rect 36244 44345 36301 44391
rect 36347 44345 36360 44391
rect 35260 44332 36360 44345
rect 36841 44391 37501 44420
rect 36841 44345 36854 44391
rect 36900 44345 36971 44391
rect 37017 44345 37088 44391
rect 37134 44345 37206 44391
rect 37252 44345 37324 44391
rect 37370 44345 37442 44391
rect 37488 44345 37501 44391
rect 36841 44332 37501 44345
rect 39008 44391 39326 44420
rect 39008 44345 39021 44391
rect 39067 44345 39144 44391
rect 39190 44345 39267 44391
rect 39313 44345 39326 44391
rect 39008 44332 39326 44345
rect 44799 44478 45323 44507
rect 44799 44432 44812 44478
rect 44858 44432 44925 44478
rect 44971 44432 45038 44478
rect 45084 44432 45151 44478
rect 45197 44432 45264 44478
rect 45310 44432 45323 44478
rect 44799 44419 45323 44432
rect 51789 44926 53789 44955
rect 51789 44880 51802 44926
rect 53776 44880 53789 44926
rect 51789 44851 53789 44880
rect 51789 44702 53789 44731
rect 51789 44656 51802 44702
rect 53776 44656 53789 44702
rect 51789 44627 53789 44656
rect 51789 44478 53789 44507
rect 48765 44391 49865 44420
rect 48765 44345 48778 44391
rect 48824 44345 48881 44391
rect 48927 44345 48984 44391
rect 49030 44345 49087 44391
rect 49133 44345 49190 44391
rect 49236 44345 49293 44391
rect 49339 44345 49396 44391
rect 49442 44345 49499 44391
rect 49545 44345 49602 44391
rect 49852 44345 49865 44391
rect 51789 44432 51802 44478
rect 53776 44432 53789 44478
rect 51789 44419 53789 44432
rect 48765 44332 49865 44345
rect 29274 44250 30373 44283
rect 29274 44204 29317 44250
rect 29363 44204 29478 44250
rect 29524 44204 29638 44250
rect 29684 44204 29798 44250
rect 29844 44204 29959 44250
rect 30005 44204 30121 44250
rect 30167 44204 30284 44250
rect 30330 44204 30373 44250
rect 29274 44171 30373 44204
rect 54750 44250 55849 44283
rect 54750 44204 54793 44250
rect 54839 44204 54956 44250
rect 55002 44204 55118 44250
rect 55164 44204 55279 44250
rect 55325 44204 55439 44250
rect 55485 44204 55599 44250
rect 55645 44204 55760 44250
rect 55806 44204 55849 44250
rect 54750 44171 55849 44204
rect 35260 44109 36360 44122
rect 31336 44022 33336 44035
rect 31336 43976 31349 44022
rect 33323 43976 33336 44022
rect 35260 44063 35273 44109
rect 35523 44063 35580 44109
rect 35626 44063 35683 44109
rect 35729 44063 35786 44109
rect 35832 44063 35889 44109
rect 35935 44063 35992 44109
rect 36038 44063 36095 44109
rect 36141 44063 36198 44109
rect 36244 44063 36301 44109
rect 36347 44063 36360 44109
rect 35260 44034 36360 44063
rect 36841 44109 37501 44122
rect 36841 44063 36854 44109
rect 36900 44063 36971 44109
rect 37017 44063 37088 44109
rect 37134 44063 37206 44109
rect 37252 44063 37324 44109
rect 37370 44063 37442 44109
rect 37488 44063 37501 44109
rect 36841 44034 37501 44063
rect 39008 44109 39326 44122
rect 39008 44063 39021 44109
rect 39067 44063 39144 44109
rect 39190 44063 39267 44109
rect 39313 44063 39326 44109
rect 39008 44034 39326 44063
rect 48765 44109 49865 44122
rect 31336 43947 33336 43976
rect 31336 43798 33336 43827
rect 31336 43752 31349 43798
rect 33323 43752 33336 43798
rect 31336 43723 33336 43752
rect 31336 43574 33336 43603
rect 31336 43528 31349 43574
rect 33323 43528 33336 43574
rect 31336 43499 33336 43528
rect 29274 43350 30373 43383
rect 29274 43304 29317 43350
rect 29363 43304 29478 43350
rect 29524 43304 29638 43350
rect 29684 43304 29798 43350
rect 29844 43304 29959 43350
rect 30005 43304 30121 43350
rect 30167 43304 30284 43350
rect 30330 43304 30373 43350
rect 29274 43271 30373 43304
rect 35260 43885 36360 43914
rect 35260 43839 35273 43885
rect 35523 43839 35580 43885
rect 35626 43839 35683 43885
rect 35729 43839 35786 43885
rect 35832 43839 35889 43885
rect 35935 43839 35992 43885
rect 36038 43839 36095 43885
rect 36141 43839 36198 43885
rect 36244 43839 36301 43885
rect 36347 43839 36360 43885
rect 35260 43810 36360 43839
rect 36841 43885 37501 43914
rect 36841 43839 36854 43885
rect 36900 43839 36971 43885
rect 37017 43839 37088 43885
rect 37134 43839 37206 43885
rect 37252 43839 37324 43885
rect 37370 43839 37442 43885
rect 37488 43839 37501 43885
rect 36841 43810 37501 43839
rect 48765 44063 48778 44109
rect 48824 44063 48881 44109
rect 48927 44063 48984 44109
rect 49030 44063 49087 44109
rect 49133 44063 49190 44109
rect 49236 44063 49293 44109
rect 49339 44063 49396 44109
rect 49442 44063 49499 44109
rect 49545 44063 49602 44109
rect 49852 44063 49865 44109
rect 44799 44022 45323 44035
rect 48765 44034 49865 44063
rect 44799 43976 44812 44022
rect 44858 43976 44925 44022
rect 44971 43976 45038 44022
rect 45084 43976 45151 44022
rect 45197 43976 45264 44022
rect 45310 43976 45323 44022
rect 44799 43947 45323 43976
rect 39008 43885 39326 43914
rect 39008 43839 39021 43885
rect 39067 43839 39144 43885
rect 39190 43839 39267 43885
rect 39313 43839 39326 43885
rect 39008 43826 39326 43839
rect 51789 44022 53789 44035
rect 44799 43798 45323 43827
rect 44799 43752 44812 43798
rect 44858 43752 44925 43798
rect 44971 43752 45038 43798
rect 45084 43752 45151 43798
rect 45197 43752 45264 43798
rect 45310 43752 45323 43798
rect 44799 43723 45323 43752
rect 48765 43885 49865 43914
rect 48765 43839 48778 43885
rect 48824 43839 48881 43885
rect 48927 43839 48984 43885
rect 49030 43839 49087 43885
rect 49133 43839 49190 43885
rect 49236 43839 49293 43885
rect 49339 43839 49396 43885
rect 49442 43839 49499 43885
rect 49545 43839 49602 43885
rect 49852 43839 49865 43885
rect 48765 43810 49865 43839
rect 51789 43976 51802 44022
rect 53776 43976 53789 44022
rect 51789 43947 53789 43976
rect 35260 43661 36360 43690
rect 35260 43615 35273 43661
rect 35523 43615 35580 43661
rect 35626 43615 35683 43661
rect 35729 43615 35786 43661
rect 35832 43615 35889 43661
rect 35935 43615 35992 43661
rect 36038 43615 36095 43661
rect 36141 43615 36198 43661
rect 36244 43615 36301 43661
rect 36347 43615 36360 43661
rect 35260 43602 36360 43615
rect 36841 43661 37501 43690
rect 36841 43615 36854 43661
rect 36900 43615 36971 43661
rect 37017 43615 37088 43661
rect 37134 43615 37206 43661
rect 37252 43615 37324 43661
rect 37370 43615 37442 43661
rect 37488 43615 37501 43661
rect 36841 43602 37501 43615
rect 48765 43661 49865 43690
rect 48765 43615 48778 43661
rect 48824 43615 48881 43661
rect 48927 43615 48984 43661
rect 49030 43615 49087 43661
rect 49133 43615 49190 43661
rect 49236 43615 49293 43661
rect 49339 43615 49396 43661
rect 49442 43615 49499 43661
rect 49545 43615 49602 43661
rect 49852 43615 49865 43661
rect 44799 43574 45323 43603
rect 48765 43602 49865 43615
rect 44799 43528 44812 43574
rect 44858 43528 44925 43574
rect 44971 43528 45038 43574
rect 45084 43528 45151 43574
rect 45197 43528 45264 43574
rect 45310 43528 45323 43574
rect 31336 43350 33336 43379
rect 31336 43304 31349 43350
rect 33323 43304 33336 43350
rect 31336 43275 33336 43304
rect 31336 43126 33336 43155
rect 31336 43080 31349 43126
rect 33323 43080 33336 43126
rect 31336 43051 33336 43080
rect 31336 42902 33336 42931
rect 31336 42856 31349 42902
rect 33323 42856 33336 42902
rect 31336 42827 33336 42856
rect 44799 43499 45323 43528
rect 51789 43798 53789 43827
rect 51789 43752 51802 43798
rect 53776 43752 53789 43798
rect 51789 43723 53789 43752
rect 51789 43574 53789 43603
rect 51789 43528 51802 43574
rect 53776 43528 53789 43574
rect 51789 43499 53789 43528
rect 44799 43350 45323 43379
rect 44799 43304 44812 43350
rect 44858 43304 44925 43350
rect 44971 43304 45038 43350
rect 45084 43304 45151 43350
rect 45197 43304 45264 43350
rect 45310 43304 45323 43350
rect 44799 43275 45323 43304
rect 51789 43350 53789 43379
rect 51789 43304 51802 43350
rect 53776 43304 53789 43350
rect 51789 43275 53789 43304
rect 35260 43039 36360 43052
rect 35260 42993 35273 43039
rect 35523 42993 35580 43039
rect 35626 42993 35683 43039
rect 35729 42993 35786 43039
rect 35832 42993 35889 43039
rect 35935 42993 35992 43039
rect 36038 42993 36095 43039
rect 36141 42993 36198 43039
rect 36244 42993 36301 43039
rect 36347 42993 36360 43039
rect 35260 42964 36360 42993
rect 36841 43039 37501 43052
rect 36841 42993 36854 43039
rect 36900 42993 36971 43039
rect 37017 42993 37088 43039
rect 37134 42993 37206 43039
rect 37252 42993 37324 43039
rect 37370 42993 37442 43039
rect 37488 42993 37501 43039
rect 36841 42964 37501 42993
rect 44799 43126 45323 43155
rect 44799 43080 44812 43126
rect 44858 43080 44925 43126
rect 44971 43080 45038 43126
rect 45084 43080 45151 43126
rect 45197 43080 45264 43126
rect 45310 43080 45323 43126
rect 54750 43350 55849 43383
rect 54750 43304 54793 43350
rect 54839 43304 54956 43350
rect 55002 43304 55118 43350
rect 55164 43304 55279 43350
rect 55325 43304 55439 43350
rect 55485 43304 55599 43350
rect 55645 43304 55760 43350
rect 55806 43304 55849 43350
rect 54750 43271 55849 43304
rect 44799 43051 45323 43080
rect 31336 42678 33336 42707
rect 31336 42632 31349 42678
rect 33323 42632 33336 42678
rect 35260 42815 36360 42844
rect 35260 42769 35273 42815
rect 35523 42769 35580 42815
rect 35626 42769 35683 42815
rect 35729 42769 35786 42815
rect 35832 42769 35889 42815
rect 35935 42769 35992 42815
rect 36038 42769 36095 42815
rect 36141 42769 36198 42815
rect 36244 42769 36301 42815
rect 36347 42769 36360 42815
rect 35260 42740 36360 42769
rect 31336 42619 33336 42632
rect 48765 43039 49865 43052
rect 48765 42993 48778 43039
rect 48824 42993 48881 43039
rect 48927 42993 48984 43039
rect 49030 42993 49087 43039
rect 49133 42993 49190 43039
rect 49236 42993 49293 43039
rect 49339 42993 49396 43039
rect 49442 42993 49499 43039
rect 49545 42993 49602 43039
rect 49852 42993 49865 43039
rect 48765 42964 49865 42993
rect 36841 42815 37501 42844
rect 36841 42769 36854 42815
rect 36900 42769 36971 42815
rect 37017 42769 37088 42815
rect 37134 42769 37206 42815
rect 37252 42769 37324 42815
rect 37370 42769 37442 42815
rect 37488 42769 37501 42815
rect 36841 42740 37501 42769
rect 39008 42815 39326 42828
rect 39008 42769 39021 42815
rect 39067 42769 39144 42815
rect 39190 42769 39267 42815
rect 39313 42769 39326 42815
rect 39008 42740 39326 42769
rect 44799 42902 45323 42931
rect 44799 42856 44812 42902
rect 44858 42856 44925 42902
rect 44971 42856 45038 42902
rect 45084 42856 45151 42902
rect 45197 42856 45264 42902
rect 45310 42856 45323 42902
rect 44799 42827 45323 42856
rect 48765 42815 49865 42844
rect 48765 42769 48778 42815
rect 48824 42769 48881 42815
rect 48927 42769 48984 42815
rect 49030 42769 49087 42815
rect 49133 42769 49190 42815
rect 49236 42769 49293 42815
rect 49339 42769 49396 42815
rect 49442 42769 49499 42815
rect 49545 42769 49602 42815
rect 49852 42769 49865 42815
rect 48765 42740 49865 42769
rect 35260 42591 36360 42620
rect 35260 42545 35273 42591
rect 35523 42545 35580 42591
rect 35626 42545 35683 42591
rect 35729 42545 35786 42591
rect 35832 42545 35889 42591
rect 35935 42545 35992 42591
rect 36038 42545 36095 42591
rect 36141 42545 36198 42591
rect 36244 42545 36301 42591
rect 36347 42545 36360 42591
rect 35260 42532 36360 42545
rect 36841 42591 37501 42620
rect 36841 42545 36854 42591
rect 36900 42545 36971 42591
rect 37017 42545 37088 42591
rect 37134 42545 37206 42591
rect 37252 42545 37324 42591
rect 37370 42545 37442 42591
rect 37488 42545 37501 42591
rect 36841 42532 37501 42545
rect 39008 42591 39326 42620
rect 39008 42545 39021 42591
rect 39067 42545 39144 42591
rect 39190 42545 39267 42591
rect 39313 42545 39326 42591
rect 39008 42532 39326 42545
rect 44799 42678 45323 42707
rect 44799 42632 44812 42678
rect 44858 42632 44925 42678
rect 44971 42632 45038 42678
rect 45084 42632 45151 42678
rect 45197 42632 45264 42678
rect 45310 42632 45323 42678
rect 44799 42619 45323 42632
rect 51789 43126 53789 43155
rect 51789 43080 51802 43126
rect 53776 43080 53789 43126
rect 51789 43051 53789 43080
rect 51789 42902 53789 42931
rect 51789 42856 51802 42902
rect 53776 42856 53789 42902
rect 51789 42827 53789 42856
rect 51789 42678 53789 42707
rect 48765 42591 49865 42620
rect 48765 42545 48778 42591
rect 48824 42545 48881 42591
rect 48927 42545 48984 42591
rect 49030 42545 49087 42591
rect 49133 42545 49190 42591
rect 49236 42545 49293 42591
rect 49339 42545 49396 42591
rect 49442 42545 49499 42591
rect 49545 42545 49602 42591
rect 49852 42545 49865 42591
rect 51789 42632 51802 42678
rect 53776 42632 53789 42678
rect 51789 42619 53789 42632
rect 48765 42532 49865 42545
rect 29274 42450 30373 42483
rect 29274 42404 29317 42450
rect 29363 42404 29478 42450
rect 29524 42404 29638 42450
rect 29684 42404 29798 42450
rect 29844 42404 29959 42450
rect 30005 42404 30121 42450
rect 30167 42404 30284 42450
rect 30330 42404 30373 42450
rect 29274 42371 30373 42404
rect 54750 42450 55849 42483
rect 54750 42404 54793 42450
rect 54839 42404 54956 42450
rect 55002 42404 55118 42450
rect 55164 42404 55279 42450
rect 55325 42404 55439 42450
rect 55485 42404 55599 42450
rect 55645 42404 55760 42450
rect 55806 42404 55849 42450
rect 54750 42371 55849 42404
rect 35260 42309 36360 42322
rect 31336 42222 33336 42235
rect 31336 42176 31349 42222
rect 33323 42176 33336 42222
rect 35260 42263 35273 42309
rect 35523 42263 35580 42309
rect 35626 42263 35683 42309
rect 35729 42263 35786 42309
rect 35832 42263 35889 42309
rect 35935 42263 35992 42309
rect 36038 42263 36095 42309
rect 36141 42263 36198 42309
rect 36244 42263 36301 42309
rect 36347 42263 36360 42309
rect 35260 42234 36360 42263
rect 36841 42309 37501 42322
rect 36841 42263 36854 42309
rect 36900 42263 36971 42309
rect 37017 42263 37088 42309
rect 37134 42263 37206 42309
rect 37252 42263 37324 42309
rect 37370 42263 37442 42309
rect 37488 42263 37501 42309
rect 36841 42234 37501 42263
rect 39008 42309 39326 42322
rect 39008 42263 39021 42309
rect 39067 42263 39144 42309
rect 39190 42263 39267 42309
rect 39313 42263 39326 42309
rect 39008 42234 39326 42263
rect 48765 42309 49865 42322
rect 31336 42147 33336 42176
rect 31336 41998 33336 42027
rect 31336 41952 31349 41998
rect 33323 41952 33336 41998
rect 31336 41923 33336 41952
rect 31336 41774 33336 41803
rect 31336 41728 31349 41774
rect 33323 41728 33336 41774
rect 31336 41699 33336 41728
rect 29274 41550 30373 41583
rect 29274 41504 29317 41550
rect 29363 41504 29478 41550
rect 29524 41504 29638 41550
rect 29684 41504 29798 41550
rect 29844 41504 29959 41550
rect 30005 41504 30121 41550
rect 30167 41504 30284 41550
rect 30330 41504 30373 41550
rect 29274 41471 30373 41504
rect 35260 42085 36360 42114
rect 35260 42039 35273 42085
rect 35523 42039 35580 42085
rect 35626 42039 35683 42085
rect 35729 42039 35786 42085
rect 35832 42039 35889 42085
rect 35935 42039 35992 42085
rect 36038 42039 36095 42085
rect 36141 42039 36198 42085
rect 36244 42039 36301 42085
rect 36347 42039 36360 42085
rect 35260 42010 36360 42039
rect 36841 42085 37501 42114
rect 36841 42039 36854 42085
rect 36900 42039 36971 42085
rect 37017 42039 37088 42085
rect 37134 42039 37206 42085
rect 37252 42039 37324 42085
rect 37370 42039 37442 42085
rect 37488 42039 37501 42085
rect 36841 42010 37501 42039
rect 48765 42263 48778 42309
rect 48824 42263 48881 42309
rect 48927 42263 48984 42309
rect 49030 42263 49087 42309
rect 49133 42263 49190 42309
rect 49236 42263 49293 42309
rect 49339 42263 49396 42309
rect 49442 42263 49499 42309
rect 49545 42263 49602 42309
rect 49852 42263 49865 42309
rect 44799 42222 45323 42235
rect 48765 42234 49865 42263
rect 44799 42176 44812 42222
rect 44858 42176 44925 42222
rect 44971 42176 45038 42222
rect 45084 42176 45151 42222
rect 45197 42176 45264 42222
rect 45310 42176 45323 42222
rect 44799 42147 45323 42176
rect 39008 42085 39326 42114
rect 39008 42039 39021 42085
rect 39067 42039 39144 42085
rect 39190 42039 39267 42085
rect 39313 42039 39326 42085
rect 39008 42026 39326 42039
rect 51789 42222 53789 42235
rect 44799 41998 45323 42027
rect 44799 41952 44812 41998
rect 44858 41952 44925 41998
rect 44971 41952 45038 41998
rect 45084 41952 45151 41998
rect 45197 41952 45264 41998
rect 45310 41952 45323 41998
rect 44799 41923 45323 41952
rect 48765 42085 49865 42114
rect 48765 42039 48778 42085
rect 48824 42039 48881 42085
rect 48927 42039 48984 42085
rect 49030 42039 49087 42085
rect 49133 42039 49190 42085
rect 49236 42039 49293 42085
rect 49339 42039 49396 42085
rect 49442 42039 49499 42085
rect 49545 42039 49602 42085
rect 49852 42039 49865 42085
rect 48765 42010 49865 42039
rect 51789 42176 51802 42222
rect 53776 42176 53789 42222
rect 51789 42147 53789 42176
rect 35260 41861 36360 41890
rect 35260 41815 35273 41861
rect 35523 41815 35580 41861
rect 35626 41815 35683 41861
rect 35729 41815 35786 41861
rect 35832 41815 35889 41861
rect 35935 41815 35992 41861
rect 36038 41815 36095 41861
rect 36141 41815 36198 41861
rect 36244 41815 36301 41861
rect 36347 41815 36360 41861
rect 35260 41802 36360 41815
rect 36841 41861 37501 41890
rect 36841 41815 36854 41861
rect 36900 41815 36971 41861
rect 37017 41815 37088 41861
rect 37134 41815 37206 41861
rect 37252 41815 37324 41861
rect 37370 41815 37442 41861
rect 37488 41815 37501 41861
rect 36841 41802 37501 41815
rect 48765 41861 49865 41890
rect 48765 41815 48778 41861
rect 48824 41815 48881 41861
rect 48927 41815 48984 41861
rect 49030 41815 49087 41861
rect 49133 41815 49190 41861
rect 49236 41815 49293 41861
rect 49339 41815 49396 41861
rect 49442 41815 49499 41861
rect 49545 41815 49602 41861
rect 49852 41815 49865 41861
rect 44799 41774 45323 41803
rect 48765 41802 49865 41815
rect 44799 41728 44812 41774
rect 44858 41728 44925 41774
rect 44971 41728 45038 41774
rect 45084 41728 45151 41774
rect 45197 41728 45264 41774
rect 45310 41728 45323 41774
rect 31336 41550 33336 41579
rect 31336 41504 31349 41550
rect 33323 41504 33336 41550
rect 31336 41475 33336 41504
rect 31336 41326 33336 41355
rect 31336 41280 31349 41326
rect 33323 41280 33336 41326
rect 31336 41251 33336 41280
rect 31336 41102 33336 41131
rect 31336 41056 31349 41102
rect 33323 41056 33336 41102
rect 31336 41027 33336 41056
rect 44799 41699 45323 41728
rect 51789 41998 53789 42027
rect 51789 41952 51802 41998
rect 53776 41952 53789 41998
rect 51789 41923 53789 41952
rect 51789 41774 53789 41803
rect 51789 41728 51802 41774
rect 53776 41728 53789 41774
rect 51789 41699 53789 41728
rect 44799 41550 45323 41579
rect 44799 41504 44812 41550
rect 44858 41504 44925 41550
rect 44971 41504 45038 41550
rect 45084 41504 45151 41550
rect 45197 41504 45264 41550
rect 45310 41504 45323 41550
rect 44799 41475 45323 41504
rect 51789 41550 53789 41579
rect 51789 41504 51802 41550
rect 53776 41504 53789 41550
rect 51789 41475 53789 41504
rect 35260 41239 36360 41252
rect 35260 41193 35273 41239
rect 35523 41193 35580 41239
rect 35626 41193 35683 41239
rect 35729 41193 35786 41239
rect 35832 41193 35889 41239
rect 35935 41193 35992 41239
rect 36038 41193 36095 41239
rect 36141 41193 36198 41239
rect 36244 41193 36301 41239
rect 36347 41193 36360 41239
rect 35260 41164 36360 41193
rect 36841 41239 37501 41252
rect 36841 41193 36854 41239
rect 36900 41193 36971 41239
rect 37017 41193 37088 41239
rect 37134 41193 37206 41239
rect 37252 41193 37324 41239
rect 37370 41193 37442 41239
rect 37488 41193 37501 41239
rect 36841 41164 37501 41193
rect 44799 41326 45323 41355
rect 44799 41280 44812 41326
rect 44858 41280 44925 41326
rect 44971 41280 45038 41326
rect 45084 41280 45151 41326
rect 45197 41280 45264 41326
rect 45310 41280 45323 41326
rect 54750 41550 55849 41583
rect 54750 41504 54793 41550
rect 54839 41504 54956 41550
rect 55002 41504 55118 41550
rect 55164 41504 55279 41550
rect 55325 41504 55439 41550
rect 55485 41504 55599 41550
rect 55645 41504 55760 41550
rect 55806 41504 55849 41550
rect 54750 41471 55849 41504
rect 44799 41251 45323 41280
rect 31336 40878 33336 40907
rect 31336 40832 31349 40878
rect 33323 40832 33336 40878
rect 35260 41015 36360 41044
rect 35260 40969 35273 41015
rect 35523 40969 35580 41015
rect 35626 40969 35683 41015
rect 35729 40969 35786 41015
rect 35832 40969 35889 41015
rect 35935 40969 35992 41015
rect 36038 40969 36095 41015
rect 36141 40969 36198 41015
rect 36244 40969 36301 41015
rect 36347 40969 36360 41015
rect 35260 40940 36360 40969
rect 31336 40819 33336 40832
rect 48765 41239 49865 41252
rect 48765 41193 48778 41239
rect 48824 41193 48881 41239
rect 48927 41193 48984 41239
rect 49030 41193 49087 41239
rect 49133 41193 49190 41239
rect 49236 41193 49293 41239
rect 49339 41193 49396 41239
rect 49442 41193 49499 41239
rect 49545 41193 49602 41239
rect 49852 41193 49865 41239
rect 48765 41164 49865 41193
rect 36841 41015 37501 41044
rect 36841 40969 36854 41015
rect 36900 40969 36971 41015
rect 37017 40969 37088 41015
rect 37134 40969 37206 41015
rect 37252 40969 37324 41015
rect 37370 40969 37442 41015
rect 37488 40969 37501 41015
rect 36841 40940 37501 40969
rect 39008 41015 39326 41028
rect 39008 40969 39021 41015
rect 39067 40969 39144 41015
rect 39190 40969 39267 41015
rect 39313 40969 39326 41015
rect 39008 40940 39326 40969
rect 44799 41102 45323 41131
rect 44799 41056 44812 41102
rect 44858 41056 44925 41102
rect 44971 41056 45038 41102
rect 45084 41056 45151 41102
rect 45197 41056 45264 41102
rect 45310 41056 45323 41102
rect 44799 41027 45323 41056
rect 48765 41015 49865 41044
rect 48765 40969 48778 41015
rect 48824 40969 48881 41015
rect 48927 40969 48984 41015
rect 49030 40969 49087 41015
rect 49133 40969 49190 41015
rect 49236 40969 49293 41015
rect 49339 40969 49396 41015
rect 49442 40969 49499 41015
rect 49545 40969 49602 41015
rect 49852 40969 49865 41015
rect 48765 40940 49865 40969
rect 35260 40791 36360 40820
rect 35260 40745 35273 40791
rect 35523 40745 35580 40791
rect 35626 40745 35683 40791
rect 35729 40745 35786 40791
rect 35832 40745 35889 40791
rect 35935 40745 35992 40791
rect 36038 40745 36095 40791
rect 36141 40745 36198 40791
rect 36244 40745 36301 40791
rect 36347 40745 36360 40791
rect 35260 40732 36360 40745
rect 36841 40791 37501 40820
rect 36841 40745 36854 40791
rect 36900 40745 36971 40791
rect 37017 40745 37088 40791
rect 37134 40745 37206 40791
rect 37252 40745 37324 40791
rect 37370 40745 37442 40791
rect 37488 40745 37501 40791
rect 36841 40732 37501 40745
rect 39008 40791 39326 40820
rect 39008 40745 39021 40791
rect 39067 40745 39144 40791
rect 39190 40745 39267 40791
rect 39313 40745 39326 40791
rect 39008 40732 39326 40745
rect 44799 40878 45323 40907
rect 44799 40832 44812 40878
rect 44858 40832 44925 40878
rect 44971 40832 45038 40878
rect 45084 40832 45151 40878
rect 45197 40832 45264 40878
rect 45310 40832 45323 40878
rect 44799 40819 45323 40832
rect 51789 41326 53789 41355
rect 51789 41280 51802 41326
rect 53776 41280 53789 41326
rect 51789 41251 53789 41280
rect 51789 41102 53789 41131
rect 51789 41056 51802 41102
rect 53776 41056 53789 41102
rect 51789 41027 53789 41056
rect 51789 40878 53789 40907
rect 48765 40791 49865 40820
rect 48765 40745 48778 40791
rect 48824 40745 48881 40791
rect 48927 40745 48984 40791
rect 49030 40745 49087 40791
rect 49133 40745 49190 40791
rect 49236 40745 49293 40791
rect 49339 40745 49396 40791
rect 49442 40745 49499 40791
rect 49545 40745 49602 40791
rect 49852 40745 49865 40791
rect 51789 40832 51802 40878
rect 53776 40832 53789 40878
rect 51789 40819 53789 40832
rect 48765 40732 49865 40745
rect 29274 40650 30373 40683
rect 29274 40604 29317 40650
rect 29363 40604 29478 40650
rect 29524 40604 29638 40650
rect 29684 40604 29798 40650
rect 29844 40604 29959 40650
rect 30005 40604 30121 40650
rect 30167 40604 30284 40650
rect 30330 40604 30373 40650
rect 29274 40571 30373 40604
rect 54750 40650 55849 40683
rect 54750 40604 54793 40650
rect 54839 40604 54956 40650
rect 55002 40604 55118 40650
rect 55164 40604 55279 40650
rect 55325 40604 55439 40650
rect 55485 40604 55599 40650
rect 55645 40604 55760 40650
rect 55806 40604 55849 40650
rect 54750 40571 55849 40604
rect 35260 40509 36360 40522
rect 31336 40422 33336 40435
rect 31336 40376 31349 40422
rect 33323 40376 33336 40422
rect 35260 40463 35273 40509
rect 35523 40463 35580 40509
rect 35626 40463 35683 40509
rect 35729 40463 35786 40509
rect 35832 40463 35889 40509
rect 35935 40463 35992 40509
rect 36038 40463 36095 40509
rect 36141 40463 36198 40509
rect 36244 40463 36301 40509
rect 36347 40463 36360 40509
rect 35260 40434 36360 40463
rect 36841 40509 37501 40522
rect 36841 40463 36854 40509
rect 36900 40463 36971 40509
rect 37017 40463 37088 40509
rect 37134 40463 37206 40509
rect 37252 40463 37324 40509
rect 37370 40463 37442 40509
rect 37488 40463 37501 40509
rect 36841 40434 37501 40463
rect 39008 40509 39326 40522
rect 39008 40463 39021 40509
rect 39067 40463 39144 40509
rect 39190 40463 39267 40509
rect 39313 40463 39326 40509
rect 39008 40434 39326 40463
rect 48765 40509 49865 40522
rect 31336 40347 33336 40376
rect 31336 40198 33336 40227
rect 31336 40152 31349 40198
rect 33323 40152 33336 40198
rect 31336 40123 33336 40152
rect 31336 39974 33336 40003
rect 31336 39928 31349 39974
rect 33323 39928 33336 39974
rect 31336 39899 33336 39928
rect 29274 39750 30373 39783
rect 29274 39704 29317 39750
rect 29363 39704 29478 39750
rect 29524 39704 29638 39750
rect 29684 39704 29798 39750
rect 29844 39704 29959 39750
rect 30005 39704 30121 39750
rect 30167 39704 30284 39750
rect 30330 39704 30373 39750
rect 29274 39671 30373 39704
rect 35260 40285 36360 40314
rect 35260 40239 35273 40285
rect 35523 40239 35580 40285
rect 35626 40239 35683 40285
rect 35729 40239 35786 40285
rect 35832 40239 35889 40285
rect 35935 40239 35992 40285
rect 36038 40239 36095 40285
rect 36141 40239 36198 40285
rect 36244 40239 36301 40285
rect 36347 40239 36360 40285
rect 35260 40210 36360 40239
rect 36841 40285 37501 40314
rect 36841 40239 36854 40285
rect 36900 40239 36971 40285
rect 37017 40239 37088 40285
rect 37134 40239 37206 40285
rect 37252 40239 37324 40285
rect 37370 40239 37442 40285
rect 37488 40239 37501 40285
rect 36841 40210 37501 40239
rect 48765 40463 48778 40509
rect 48824 40463 48881 40509
rect 48927 40463 48984 40509
rect 49030 40463 49087 40509
rect 49133 40463 49190 40509
rect 49236 40463 49293 40509
rect 49339 40463 49396 40509
rect 49442 40463 49499 40509
rect 49545 40463 49602 40509
rect 49852 40463 49865 40509
rect 44799 40422 45323 40435
rect 48765 40434 49865 40463
rect 44799 40376 44812 40422
rect 44858 40376 44925 40422
rect 44971 40376 45038 40422
rect 45084 40376 45151 40422
rect 45197 40376 45264 40422
rect 45310 40376 45323 40422
rect 44799 40347 45323 40376
rect 39008 40285 39326 40314
rect 39008 40239 39021 40285
rect 39067 40239 39144 40285
rect 39190 40239 39267 40285
rect 39313 40239 39326 40285
rect 39008 40226 39326 40239
rect 51789 40422 53789 40435
rect 44799 40198 45323 40227
rect 44799 40152 44812 40198
rect 44858 40152 44925 40198
rect 44971 40152 45038 40198
rect 45084 40152 45151 40198
rect 45197 40152 45264 40198
rect 45310 40152 45323 40198
rect 44799 40123 45323 40152
rect 48765 40285 49865 40314
rect 48765 40239 48778 40285
rect 48824 40239 48881 40285
rect 48927 40239 48984 40285
rect 49030 40239 49087 40285
rect 49133 40239 49190 40285
rect 49236 40239 49293 40285
rect 49339 40239 49396 40285
rect 49442 40239 49499 40285
rect 49545 40239 49602 40285
rect 49852 40239 49865 40285
rect 48765 40210 49865 40239
rect 51789 40376 51802 40422
rect 53776 40376 53789 40422
rect 51789 40347 53789 40376
rect 35260 40061 36360 40090
rect 35260 40015 35273 40061
rect 35523 40015 35580 40061
rect 35626 40015 35683 40061
rect 35729 40015 35786 40061
rect 35832 40015 35889 40061
rect 35935 40015 35992 40061
rect 36038 40015 36095 40061
rect 36141 40015 36198 40061
rect 36244 40015 36301 40061
rect 36347 40015 36360 40061
rect 35260 40002 36360 40015
rect 36841 40061 37501 40090
rect 36841 40015 36854 40061
rect 36900 40015 36971 40061
rect 37017 40015 37088 40061
rect 37134 40015 37206 40061
rect 37252 40015 37324 40061
rect 37370 40015 37442 40061
rect 37488 40015 37501 40061
rect 36841 40002 37501 40015
rect 48765 40061 49865 40090
rect 48765 40015 48778 40061
rect 48824 40015 48881 40061
rect 48927 40015 48984 40061
rect 49030 40015 49087 40061
rect 49133 40015 49190 40061
rect 49236 40015 49293 40061
rect 49339 40015 49396 40061
rect 49442 40015 49499 40061
rect 49545 40015 49602 40061
rect 49852 40015 49865 40061
rect 44799 39974 45323 40003
rect 48765 40002 49865 40015
rect 44799 39928 44812 39974
rect 44858 39928 44925 39974
rect 44971 39928 45038 39974
rect 45084 39928 45151 39974
rect 45197 39928 45264 39974
rect 45310 39928 45323 39974
rect 31336 39750 33336 39779
rect 31336 39704 31349 39750
rect 33323 39704 33336 39750
rect 31336 39675 33336 39704
rect 31336 39526 33336 39555
rect 31336 39480 31349 39526
rect 33323 39480 33336 39526
rect 31336 39451 33336 39480
rect 31336 39302 33336 39331
rect 31336 39256 31349 39302
rect 33323 39256 33336 39302
rect 31336 39227 33336 39256
rect 44799 39899 45323 39928
rect 51789 40198 53789 40227
rect 51789 40152 51802 40198
rect 53776 40152 53789 40198
rect 51789 40123 53789 40152
rect 51789 39974 53789 40003
rect 51789 39928 51802 39974
rect 53776 39928 53789 39974
rect 51789 39899 53789 39928
rect 44799 39750 45323 39779
rect 44799 39704 44812 39750
rect 44858 39704 44925 39750
rect 44971 39704 45038 39750
rect 45084 39704 45151 39750
rect 45197 39704 45264 39750
rect 45310 39704 45323 39750
rect 44799 39675 45323 39704
rect 51789 39750 53789 39779
rect 51789 39704 51802 39750
rect 53776 39704 53789 39750
rect 51789 39675 53789 39704
rect 35260 39439 36360 39452
rect 35260 39393 35273 39439
rect 35523 39393 35580 39439
rect 35626 39393 35683 39439
rect 35729 39393 35786 39439
rect 35832 39393 35889 39439
rect 35935 39393 35992 39439
rect 36038 39393 36095 39439
rect 36141 39393 36198 39439
rect 36244 39393 36301 39439
rect 36347 39393 36360 39439
rect 35260 39364 36360 39393
rect 36841 39439 37501 39452
rect 36841 39393 36854 39439
rect 36900 39393 36971 39439
rect 37017 39393 37088 39439
rect 37134 39393 37206 39439
rect 37252 39393 37324 39439
rect 37370 39393 37442 39439
rect 37488 39393 37501 39439
rect 36841 39364 37501 39393
rect 44799 39526 45323 39555
rect 44799 39480 44812 39526
rect 44858 39480 44925 39526
rect 44971 39480 45038 39526
rect 45084 39480 45151 39526
rect 45197 39480 45264 39526
rect 45310 39480 45323 39526
rect 54750 39750 55849 39783
rect 54750 39704 54793 39750
rect 54839 39704 54956 39750
rect 55002 39704 55118 39750
rect 55164 39704 55279 39750
rect 55325 39704 55439 39750
rect 55485 39704 55599 39750
rect 55645 39704 55760 39750
rect 55806 39704 55849 39750
rect 54750 39671 55849 39704
rect 44799 39451 45323 39480
rect 31336 39078 33336 39107
rect 31336 39032 31349 39078
rect 33323 39032 33336 39078
rect 35260 39215 36360 39244
rect 35260 39169 35273 39215
rect 35523 39169 35580 39215
rect 35626 39169 35683 39215
rect 35729 39169 35786 39215
rect 35832 39169 35889 39215
rect 35935 39169 35992 39215
rect 36038 39169 36095 39215
rect 36141 39169 36198 39215
rect 36244 39169 36301 39215
rect 36347 39169 36360 39215
rect 35260 39140 36360 39169
rect 31336 39019 33336 39032
rect 48765 39439 49865 39452
rect 48765 39393 48778 39439
rect 48824 39393 48881 39439
rect 48927 39393 48984 39439
rect 49030 39393 49087 39439
rect 49133 39393 49190 39439
rect 49236 39393 49293 39439
rect 49339 39393 49396 39439
rect 49442 39393 49499 39439
rect 49545 39393 49602 39439
rect 49852 39393 49865 39439
rect 48765 39364 49865 39393
rect 36841 39215 37501 39244
rect 36841 39169 36854 39215
rect 36900 39169 36971 39215
rect 37017 39169 37088 39215
rect 37134 39169 37206 39215
rect 37252 39169 37324 39215
rect 37370 39169 37442 39215
rect 37488 39169 37501 39215
rect 36841 39140 37501 39169
rect 39008 39215 39326 39228
rect 39008 39169 39021 39215
rect 39067 39169 39144 39215
rect 39190 39169 39267 39215
rect 39313 39169 39326 39215
rect 39008 39140 39326 39169
rect 44799 39302 45323 39331
rect 44799 39256 44812 39302
rect 44858 39256 44925 39302
rect 44971 39256 45038 39302
rect 45084 39256 45151 39302
rect 45197 39256 45264 39302
rect 45310 39256 45323 39302
rect 44799 39227 45323 39256
rect 48765 39215 49865 39244
rect 48765 39169 48778 39215
rect 48824 39169 48881 39215
rect 48927 39169 48984 39215
rect 49030 39169 49087 39215
rect 49133 39169 49190 39215
rect 49236 39169 49293 39215
rect 49339 39169 49396 39215
rect 49442 39169 49499 39215
rect 49545 39169 49602 39215
rect 49852 39169 49865 39215
rect 48765 39140 49865 39169
rect 35260 38991 36360 39020
rect 35260 38945 35273 38991
rect 35523 38945 35580 38991
rect 35626 38945 35683 38991
rect 35729 38945 35786 38991
rect 35832 38945 35889 38991
rect 35935 38945 35992 38991
rect 36038 38945 36095 38991
rect 36141 38945 36198 38991
rect 36244 38945 36301 38991
rect 36347 38945 36360 38991
rect 35260 38932 36360 38945
rect 36841 38991 37501 39020
rect 36841 38945 36854 38991
rect 36900 38945 36971 38991
rect 37017 38945 37088 38991
rect 37134 38945 37206 38991
rect 37252 38945 37324 38991
rect 37370 38945 37442 38991
rect 37488 38945 37501 38991
rect 36841 38932 37501 38945
rect 39008 38991 39326 39020
rect 39008 38945 39021 38991
rect 39067 38945 39144 38991
rect 39190 38945 39267 38991
rect 39313 38945 39326 38991
rect 39008 38932 39326 38945
rect 44799 39078 45323 39107
rect 44799 39032 44812 39078
rect 44858 39032 44925 39078
rect 44971 39032 45038 39078
rect 45084 39032 45151 39078
rect 45197 39032 45264 39078
rect 45310 39032 45323 39078
rect 44799 39019 45323 39032
rect 51789 39526 53789 39555
rect 51789 39480 51802 39526
rect 53776 39480 53789 39526
rect 51789 39451 53789 39480
rect 51789 39302 53789 39331
rect 51789 39256 51802 39302
rect 53776 39256 53789 39302
rect 51789 39227 53789 39256
rect 51789 39078 53789 39107
rect 48765 38991 49865 39020
rect 48765 38945 48778 38991
rect 48824 38945 48881 38991
rect 48927 38945 48984 38991
rect 49030 38945 49087 38991
rect 49133 38945 49190 38991
rect 49236 38945 49293 38991
rect 49339 38945 49396 38991
rect 49442 38945 49499 38991
rect 49545 38945 49602 38991
rect 49852 38945 49865 38991
rect 51789 39032 51802 39078
rect 53776 39032 53789 39078
rect 51789 39019 53789 39032
rect 48765 38932 49865 38945
rect 29274 38850 30373 38883
rect 29274 38804 29317 38850
rect 29363 38804 29478 38850
rect 29524 38804 29638 38850
rect 29684 38804 29798 38850
rect 29844 38804 29959 38850
rect 30005 38804 30121 38850
rect 30167 38804 30284 38850
rect 30330 38804 30373 38850
rect 29274 38771 30373 38804
rect 54750 38850 55849 38883
rect 54750 38804 54793 38850
rect 54839 38804 54956 38850
rect 55002 38804 55118 38850
rect 55164 38804 55279 38850
rect 55325 38804 55439 38850
rect 55485 38804 55599 38850
rect 55645 38804 55760 38850
rect 55806 38804 55849 38850
rect 54750 38771 55849 38804
rect 35260 38709 36360 38722
rect 31336 38622 33336 38635
rect 31336 38576 31349 38622
rect 33323 38576 33336 38622
rect 35260 38663 35273 38709
rect 35523 38663 35580 38709
rect 35626 38663 35683 38709
rect 35729 38663 35786 38709
rect 35832 38663 35889 38709
rect 35935 38663 35992 38709
rect 36038 38663 36095 38709
rect 36141 38663 36198 38709
rect 36244 38663 36301 38709
rect 36347 38663 36360 38709
rect 35260 38634 36360 38663
rect 36841 38709 37501 38722
rect 36841 38663 36854 38709
rect 36900 38663 36971 38709
rect 37017 38663 37088 38709
rect 37134 38663 37206 38709
rect 37252 38663 37324 38709
rect 37370 38663 37442 38709
rect 37488 38663 37501 38709
rect 36841 38634 37501 38663
rect 39008 38709 39326 38722
rect 39008 38663 39021 38709
rect 39067 38663 39144 38709
rect 39190 38663 39267 38709
rect 39313 38663 39326 38709
rect 39008 38634 39326 38663
rect 48765 38709 49865 38722
rect 31336 38547 33336 38576
rect 31336 38398 33336 38427
rect 31336 38352 31349 38398
rect 33323 38352 33336 38398
rect 31336 38323 33336 38352
rect 31336 38174 33336 38203
rect 31336 38128 31349 38174
rect 33323 38128 33336 38174
rect 31336 38099 33336 38128
rect 29274 37950 30373 37983
rect 29274 37904 29317 37950
rect 29363 37904 29478 37950
rect 29524 37904 29638 37950
rect 29684 37904 29798 37950
rect 29844 37904 29959 37950
rect 30005 37904 30121 37950
rect 30167 37904 30284 37950
rect 30330 37904 30373 37950
rect 29274 37871 30373 37904
rect 35260 38485 36360 38514
rect 35260 38439 35273 38485
rect 35523 38439 35580 38485
rect 35626 38439 35683 38485
rect 35729 38439 35786 38485
rect 35832 38439 35889 38485
rect 35935 38439 35992 38485
rect 36038 38439 36095 38485
rect 36141 38439 36198 38485
rect 36244 38439 36301 38485
rect 36347 38439 36360 38485
rect 35260 38410 36360 38439
rect 36841 38485 37501 38514
rect 36841 38439 36854 38485
rect 36900 38439 36971 38485
rect 37017 38439 37088 38485
rect 37134 38439 37206 38485
rect 37252 38439 37324 38485
rect 37370 38439 37442 38485
rect 37488 38439 37501 38485
rect 36841 38410 37501 38439
rect 48765 38663 48778 38709
rect 48824 38663 48881 38709
rect 48927 38663 48984 38709
rect 49030 38663 49087 38709
rect 49133 38663 49190 38709
rect 49236 38663 49293 38709
rect 49339 38663 49396 38709
rect 49442 38663 49499 38709
rect 49545 38663 49602 38709
rect 49852 38663 49865 38709
rect 44799 38622 45323 38635
rect 48765 38634 49865 38663
rect 44799 38576 44812 38622
rect 44858 38576 44925 38622
rect 44971 38576 45038 38622
rect 45084 38576 45151 38622
rect 45197 38576 45264 38622
rect 45310 38576 45323 38622
rect 44799 38547 45323 38576
rect 39008 38485 39326 38514
rect 39008 38439 39021 38485
rect 39067 38439 39144 38485
rect 39190 38439 39267 38485
rect 39313 38439 39326 38485
rect 39008 38426 39326 38439
rect 51789 38622 53789 38635
rect 44799 38398 45323 38427
rect 44799 38352 44812 38398
rect 44858 38352 44925 38398
rect 44971 38352 45038 38398
rect 45084 38352 45151 38398
rect 45197 38352 45264 38398
rect 45310 38352 45323 38398
rect 44799 38323 45323 38352
rect 48765 38485 49865 38514
rect 48765 38439 48778 38485
rect 48824 38439 48881 38485
rect 48927 38439 48984 38485
rect 49030 38439 49087 38485
rect 49133 38439 49190 38485
rect 49236 38439 49293 38485
rect 49339 38439 49396 38485
rect 49442 38439 49499 38485
rect 49545 38439 49602 38485
rect 49852 38439 49865 38485
rect 48765 38410 49865 38439
rect 51789 38576 51802 38622
rect 53776 38576 53789 38622
rect 51789 38547 53789 38576
rect 35260 38261 36360 38290
rect 35260 38215 35273 38261
rect 35523 38215 35580 38261
rect 35626 38215 35683 38261
rect 35729 38215 35786 38261
rect 35832 38215 35889 38261
rect 35935 38215 35992 38261
rect 36038 38215 36095 38261
rect 36141 38215 36198 38261
rect 36244 38215 36301 38261
rect 36347 38215 36360 38261
rect 35260 38202 36360 38215
rect 36841 38261 37501 38290
rect 36841 38215 36854 38261
rect 36900 38215 36971 38261
rect 37017 38215 37088 38261
rect 37134 38215 37206 38261
rect 37252 38215 37324 38261
rect 37370 38215 37442 38261
rect 37488 38215 37501 38261
rect 36841 38202 37501 38215
rect 48765 38261 49865 38290
rect 48765 38215 48778 38261
rect 48824 38215 48881 38261
rect 48927 38215 48984 38261
rect 49030 38215 49087 38261
rect 49133 38215 49190 38261
rect 49236 38215 49293 38261
rect 49339 38215 49396 38261
rect 49442 38215 49499 38261
rect 49545 38215 49602 38261
rect 49852 38215 49865 38261
rect 44799 38174 45323 38203
rect 48765 38202 49865 38215
rect 44799 38128 44812 38174
rect 44858 38128 44925 38174
rect 44971 38128 45038 38174
rect 45084 38128 45151 38174
rect 45197 38128 45264 38174
rect 45310 38128 45323 38174
rect 31336 37950 33336 37979
rect 31336 37904 31349 37950
rect 33323 37904 33336 37950
rect 31336 37875 33336 37904
rect 31336 37726 33336 37755
rect 31336 37680 31349 37726
rect 33323 37680 33336 37726
rect 31336 37651 33336 37680
rect 31336 37502 33336 37531
rect 31336 37456 31349 37502
rect 33323 37456 33336 37502
rect 31336 37427 33336 37456
rect 44799 38099 45323 38128
rect 51789 38398 53789 38427
rect 51789 38352 51802 38398
rect 53776 38352 53789 38398
rect 51789 38323 53789 38352
rect 51789 38174 53789 38203
rect 51789 38128 51802 38174
rect 53776 38128 53789 38174
rect 51789 38099 53789 38128
rect 44799 37950 45323 37979
rect 44799 37904 44812 37950
rect 44858 37904 44925 37950
rect 44971 37904 45038 37950
rect 45084 37904 45151 37950
rect 45197 37904 45264 37950
rect 45310 37904 45323 37950
rect 44799 37875 45323 37904
rect 51789 37950 53789 37979
rect 51789 37904 51802 37950
rect 53776 37904 53789 37950
rect 51789 37875 53789 37904
rect 35260 37639 36360 37652
rect 35260 37593 35273 37639
rect 35523 37593 35580 37639
rect 35626 37593 35683 37639
rect 35729 37593 35786 37639
rect 35832 37593 35889 37639
rect 35935 37593 35992 37639
rect 36038 37593 36095 37639
rect 36141 37593 36198 37639
rect 36244 37593 36301 37639
rect 36347 37593 36360 37639
rect 35260 37564 36360 37593
rect 36841 37639 37501 37652
rect 36841 37593 36854 37639
rect 36900 37593 36971 37639
rect 37017 37593 37088 37639
rect 37134 37593 37206 37639
rect 37252 37593 37324 37639
rect 37370 37593 37442 37639
rect 37488 37593 37501 37639
rect 36841 37564 37501 37593
rect 44799 37726 45323 37755
rect 44799 37680 44812 37726
rect 44858 37680 44925 37726
rect 44971 37680 45038 37726
rect 45084 37680 45151 37726
rect 45197 37680 45264 37726
rect 45310 37680 45323 37726
rect 54750 37950 55849 37983
rect 54750 37904 54793 37950
rect 54839 37904 54956 37950
rect 55002 37904 55118 37950
rect 55164 37904 55279 37950
rect 55325 37904 55439 37950
rect 55485 37904 55599 37950
rect 55645 37904 55760 37950
rect 55806 37904 55849 37950
rect 54750 37871 55849 37904
rect 44799 37651 45323 37680
rect 31336 37278 33336 37307
rect 31336 37232 31349 37278
rect 33323 37232 33336 37278
rect 35260 37415 36360 37444
rect 35260 37369 35273 37415
rect 35523 37369 35580 37415
rect 35626 37369 35683 37415
rect 35729 37369 35786 37415
rect 35832 37369 35889 37415
rect 35935 37369 35992 37415
rect 36038 37369 36095 37415
rect 36141 37369 36198 37415
rect 36244 37369 36301 37415
rect 36347 37369 36360 37415
rect 35260 37340 36360 37369
rect 31336 37219 33336 37232
rect 48765 37639 49865 37652
rect 48765 37593 48778 37639
rect 48824 37593 48881 37639
rect 48927 37593 48984 37639
rect 49030 37593 49087 37639
rect 49133 37593 49190 37639
rect 49236 37593 49293 37639
rect 49339 37593 49396 37639
rect 49442 37593 49499 37639
rect 49545 37593 49602 37639
rect 49852 37593 49865 37639
rect 48765 37564 49865 37593
rect 36841 37415 37501 37444
rect 36841 37369 36854 37415
rect 36900 37369 36971 37415
rect 37017 37369 37088 37415
rect 37134 37369 37206 37415
rect 37252 37369 37324 37415
rect 37370 37369 37442 37415
rect 37488 37369 37501 37415
rect 36841 37340 37501 37369
rect 39008 37415 39326 37428
rect 39008 37369 39021 37415
rect 39067 37369 39144 37415
rect 39190 37369 39267 37415
rect 39313 37369 39326 37415
rect 39008 37340 39326 37369
rect 44799 37502 45323 37531
rect 44799 37456 44812 37502
rect 44858 37456 44925 37502
rect 44971 37456 45038 37502
rect 45084 37456 45151 37502
rect 45197 37456 45264 37502
rect 45310 37456 45323 37502
rect 44799 37427 45323 37456
rect 48765 37415 49865 37444
rect 48765 37369 48778 37415
rect 48824 37369 48881 37415
rect 48927 37369 48984 37415
rect 49030 37369 49087 37415
rect 49133 37369 49190 37415
rect 49236 37369 49293 37415
rect 49339 37369 49396 37415
rect 49442 37369 49499 37415
rect 49545 37369 49602 37415
rect 49852 37369 49865 37415
rect 48765 37340 49865 37369
rect 35260 37191 36360 37220
rect 35260 37145 35273 37191
rect 35523 37145 35580 37191
rect 35626 37145 35683 37191
rect 35729 37145 35786 37191
rect 35832 37145 35889 37191
rect 35935 37145 35992 37191
rect 36038 37145 36095 37191
rect 36141 37145 36198 37191
rect 36244 37145 36301 37191
rect 36347 37145 36360 37191
rect 35260 37132 36360 37145
rect 36841 37191 37501 37220
rect 36841 37145 36854 37191
rect 36900 37145 36971 37191
rect 37017 37145 37088 37191
rect 37134 37145 37206 37191
rect 37252 37145 37324 37191
rect 37370 37145 37442 37191
rect 37488 37145 37501 37191
rect 36841 37132 37501 37145
rect 39008 37191 39326 37220
rect 39008 37145 39021 37191
rect 39067 37145 39144 37191
rect 39190 37145 39267 37191
rect 39313 37145 39326 37191
rect 39008 37132 39326 37145
rect 44799 37278 45323 37307
rect 44799 37232 44812 37278
rect 44858 37232 44925 37278
rect 44971 37232 45038 37278
rect 45084 37232 45151 37278
rect 45197 37232 45264 37278
rect 45310 37232 45323 37278
rect 44799 37219 45323 37232
rect 51789 37726 53789 37755
rect 51789 37680 51802 37726
rect 53776 37680 53789 37726
rect 51789 37651 53789 37680
rect 51789 37502 53789 37531
rect 51789 37456 51802 37502
rect 53776 37456 53789 37502
rect 51789 37427 53789 37456
rect 51789 37278 53789 37307
rect 48765 37191 49865 37220
rect 48765 37145 48778 37191
rect 48824 37145 48881 37191
rect 48927 37145 48984 37191
rect 49030 37145 49087 37191
rect 49133 37145 49190 37191
rect 49236 37145 49293 37191
rect 49339 37145 49396 37191
rect 49442 37145 49499 37191
rect 49545 37145 49602 37191
rect 49852 37145 49865 37191
rect 51789 37232 51802 37278
rect 53776 37232 53789 37278
rect 51789 37219 53789 37232
rect 48765 37132 49865 37145
rect 29274 37050 30373 37083
rect 29274 37004 29317 37050
rect 29363 37004 29478 37050
rect 29524 37004 29638 37050
rect 29684 37004 29798 37050
rect 29844 37004 29959 37050
rect 30005 37004 30121 37050
rect 30167 37004 30284 37050
rect 30330 37004 30373 37050
rect 29274 36971 30373 37004
rect 54750 37050 55849 37083
rect 54750 37004 54793 37050
rect 54839 37004 54956 37050
rect 55002 37004 55118 37050
rect 55164 37004 55279 37050
rect 55325 37004 55439 37050
rect 55485 37004 55599 37050
rect 55645 37004 55760 37050
rect 55806 37004 55849 37050
rect 54750 36971 55849 37004
rect 35260 36909 36360 36922
rect 31336 36822 33336 36835
rect 31336 36776 31349 36822
rect 33323 36776 33336 36822
rect 35260 36863 35273 36909
rect 35523 36863 35580 36909
rect 35626 36863 35683 36909
rect 35729 36863 35786 36909
rect 35832 36863 35889 36909
rect 35935 36863 35992 36909
rect 36038 36863 36095 36909
rect 36141 36863 36198 36909
rect 36244 36863 36301 36909
rect 36347 36863 36360 36909
rect 35260 36834 36360 36863
rect 36841 36909 37501 36922
rect 36841 36863 36854 36909
rect 36900 36863 36971 36909
rect 37017 36863 37088 36909
rect 37134 36863 37206 36909
rect 37252 36863 37324 36909
rect 37370 36863 37442 36909
rect 37488 36863 37501 36909
rect 36841 36834 37501 36863
rect 39008 36909 39326 36922
rect 39008 36863 39021 36909
rect 39067 36863 39144 36909
rect 39190 36863 39267 36909
rect 39313 36863 39326 36909
rect 39008 36834 39326 36863
rect 48765 36909 49865 36922
rect 31336 36747 33336 36776
rect 31336 36598 33336 36627
rect 31336 36552 31349 36598
rect 33323 36552 33336 36598
rect 31336 36523 33336 36552
rect 31336 36374 33336 36403
rect 31336 36328 31349 36374
rect 33323 36328 33336 36374
rect 31336 36299 33336 36328
rect 29274 36150 30373 36183
rect 29274 36104 29317 36150
rect 29363 36104 29478 36150
rect 29524 36104 29638 36150
rect 29684 36104 29798 36150
rect 29844 36104 29959 36150
rect 30005 36104 30121 36150
rect 30167 36104 30284 36150
rect 30330 36104 30373 36150
rect 29274 36058 30373 36104
rect 35260 36685 36360 36714
rect 35260 36639 35273 36685
rect 35523 36639 35580 36685
rect 35626 36639 35683 36685
rect 35729 36639 35786 36685
rect 35832 36639 35889 36685
rect 35935 36639 35992 36685
rect 36038 36639 36095 36685
rect 36141 36639 36198 36685
rect 36244 36639 36301 36685
rect 36347 36639 36360 36685
rect 35260 36610 36360 36639
rect 36841 36685 37501 36714
rect 36841 36639 36854 36685
rect 36900 36639 36971 36685
rect 37017 36639 37088 36685
rect 37134 36639 37206 36685
rect 37252 36639 37324 36685
rect 37370 36639 37442 36685
rect 37488 36639 37501 36685
rect 36841 36610 37501 36639
rect 48765 36863 48778 36909
rect 48824 36863 48881 36909
rect 48927 36863 48984 36909
rect 49030 36863 49087 36909
rect 49133 36863 49190 36909
rect 49236 36863 49293 36909
rect 49339 36863 49396 36909
rect 49442 36863 49499 36909
rect 49545 36863 49602 36909
rect 49852 36863 49865 36909
rect 44799 36822 45323 36835
rect 48765 36834 49865 36863
rect 44799 36776 44812 36822
rect 44858 36776 44925 36822
rect 44971 36776 45038 36822
rect 45084 36776 45151 36822
rect 45197 36776 45264 36822
rect 45310 36776 45323 36822
rect 44799 36747 45323 36776
rect 39008 36685 39326 36714
rect 39008 36639 39021 36685
rect 39067 36639 39144 36685
rect 39190 36639 39267 36685
rect 39313 36639 39326 36685
rect 39008 36626 39326 36639
rect 51789 36822 53789 36835
rect 44799 36598 45323 36627
rect 44799 36552 44812 36598
rect 44858 36552 44925 36598
rect 44971 36552 45038 36598
rect 45084 36552 45151 36598
rect 45197 36552 45264 36598
rect 45310 36552 45323 36598
rect 44799 36523 45323 36552
rect 48765 36685 49865 36714
rect 48765 36639 48778 36685
rect 48824 36639 48881 36685
rect 48927 36639 48984 36685
rect 49030 36639 49087 36685
rect 49133 36639 49190 36685
rect 49236 36639 49293 36685
rect 49339 36639 49396 36685
rect 49442 36639 49499 36685
rect 49545 36639 49602 36685
rect 49852 36639 49865 36685
rect 48765 36610 49865 36639
rect 51789 36776 51802 36822
rect 53776 36776 53789 36822
rect 51789 36747 53789 36776
rect 35260 36461 36360 36490
rect 35260 36415 35273 36461
rect 35523 36415 35580 36461
rect 35626 36415 35683 36461
rect 35729 36415 35786 36461
rect 35832 36415 35889 36461
rect 35935 36415 35992 36461
rect 36038 36415 36095 36461
rect 36141 36415 36198 36461
rect 36244 36415 36301 36461
rect 36347 36415 36360 36461
rect 35260 36402 36360 36415
rect 36841 36461 37501 36490
rect 36841 36415 36854 36461
rect 36900 36415 36971 36461
rect 37017 36415 37088 36461
rect 37134 36415 37206 36461
rect 37252 36415 37324 36461
rect 37370 36415 37442 36461
rect 37488 36415 37501 36461
rect 36841 36402 37501 36415
rect 48765 36461 49865 36490
rect 48765 36415 48778 36461
rect 48824 36415 48881 36461
rect 48927 36415 48984 36461
rect 49030 36415 49087 36461
rect 49133 36415 49190 36461
rect 49236 36415 49293 36461
rect 49339 36415 49396 36461
rect 49442 36415 49499 36461
rect 49545 36415 49602 36461
rect 49852 36415 49865 36461
rect 44799 36374 45323 36403
rect 48765 36402 49865 36415
rect 44799 36328 44812 36374
rect 44858 36328 44925 36374
rect 44971 36328 45038 36374
rect 45084 36328 45151 36374
rect 45197 36328 45264 36374
rect 45310 36328 45323 36374
rect 31336 36150 33336 36179
rect 31336 36104 31349 36150
rect 33323 36104 33336 36150
rect 31336 36091 33336 36104
rect 44799 36299 45323 36328
rect 51789 36598 53789 36627
rect 51789 36552 51802 36598
rect 53776 36552 53789 36598
rect 51789 36523 53789 36552
rect 51789 36374 53789 36403
rect 51789 36328 51802 36374
rect 53776 36328 53789 36374
rect 51789 36299 53789 36328
rect 44799 36150 45323 36179
rect 44799 36104 44812 36150
rect 44858 36104 44925 36150
rect 44971 36104 45038 36150
rect 45084 36104 45151 36150
rect 45197 36104 45264 36150
rect 45310 36104 45323 36150
rect 44799 36091 45323 36104
rect 51789 36150 53789 36179
rect 51789 36104 51802 36150
rect 53776 36104 53789 36150
rect 51789 36091 53789 36104
rect 54750 36150 55849 36183
rect 54750 36104 54793 36150
rect 54839 36104 54956 36150
rect 55002 36104 55118 36150
rect 55164 36104 55279 36150
rect 55325 36104 55439 36150
rect 55485 36104 55599 36150
rect 55645 36104 55760 36150
rect 55806 36104 55849 36150
rect 54750 36058 55849 36104
<< mvndiffc >>
rect 33014 65548 33774 65594
rect 33831 65548 33877 65594
rect 33934 65548 33980 65594
rect 34037 65548 34083 65594
rect 34140 65548 34186 65594
rect 34243 65548 34289 65594
rect 34346 65548 34392 65594
rect 34449 65548 34495 65594
rect 34552 65548 34598 65594
rect 34655 65548 34701 65594
rect 34758 65548 34804 65594
rect 34861 65548 34907 65594
rect 34964 65548 35010 65594
rect 40075 65548 40121 65594
rect 40189 65548 40235 65594
rect 40303 65548 40349 65594
rect 40417 65548 40463 65594
rect 40531 65548 40577 65594
rect 40976 65549 41022 65595
rect 41079 65549 41125 65595
rect 41182 65549 41228 65595
rect 41286 65549 41332 65595
rect 41390 65549 41436 65595
rect 41494 65549 41540 65595
rect 41598 65549 41644 65595
rect 41702 65549 41748 65595
rect 41806 65549 41852 65595
rect 41910 65549 41956 65595
rect 42014 65549 42060 65595
rect 42118 65549 42164 65595
rect 42222 65549 42268 65595
rect 33014 65324 33774 65370
rect 33831 65324 33877 65370
rect 33934 65324 33980 65370
rect 34037 65324 34083 65370
rect 34140 65324 34186 65370
rect 34243 65324 34289 65370
rect 34346 65324 34392 65370
rect 34449 65324 34495 65370
rect 34552 65324 34598 65370
rect 34655 65324 34701 65370
rect 34758 65324 34804 65370
rect 34861 65324 34907 65370
rect 34964 65324 35010 65370
rect 40075 65324 40121 65370
rect 40189 65324 40235 65370
rect 40303 65324 40349 65370
rect 40417 65324 40463 65370
rect 40531 65324 40577 65370
rect 44445 65548 44491 65594
rect 44559 65548 44605 65594
rect 44673 65548 44719 65594
rect 44787 65548 44833 65594
rect 44901 65548 44947 65594
rect 50014 65548 50774 65594
rect 50831 65548 50877 65594
rect 50934 65548 50980 65594
rect 51037 65548 51083 65594
rect 51140 65548 51186 65594
rect 51243 65548 51289 65594
rect 51346 65548 51392 65594
rect 51449 65548 51495 65594
rect 51552 65548 51598 65594
rect 51655 65548 51701 65594
rect 51758 65548 51804 65594
rect 51861 65548 51907 65594
rect 51964 65548 52010 65594
rect 40976 65325 41022 65371
rect 41079 65325 41125 65371
rect 41182 65325 41228 65371
rect 41286 65325 41332 65371
rect 41390 65325 41436 65371
rect 41494 65325 41540 65371
rect 41598 65325 41644 65371
rect 41702 65325 41748 65371
rect 41806 65325 41852 65371
rect 41910 65325 41956 65371
rect 42014 65325 42060 65371
rect 42118 65325 42164 65371
rect 42222 65325 42268 65371
rect 44445 65324 44491 65370
rect 44559 65324 44605 65370
rect 44673 65324 44719 65370
rect 44787 65324 44833 65370
rect 44901 65324 44947 65370
rect 50014 65324 50774 65370
rect 50831 65324 50877 65370
rect 50934 65324 50980 65370
rect 51037 65324 51083 65370
rect 51140 65324 51186 65370
rect 51243 65324 51289 65370
rect 51346 65324 51392 65370
rect 51449 65324 51495 65370
rect 51552 65324 51598 65370
rect 51655 65324 51701 65370
rect 51758 65324 51804 65370
rect 51861 65324 51907 65370
rect 51964 65324 52010 65370
rect 33684 64904 33730 64950
rect 33787 64904 33833 64950
rect 33890 64904 33936 64950
rect 33993 64904 34039 64950
rect 34096 64904 34142 64950
rect 34199 64904 34245 64950
rect 34302 64904 34348 64950
rect 34405 64904 34451 64950
rect 34508 64904 34554 64950
rect 34612 64904 34658 64950
rect 39740 64904 39786 64950
rect 39862 64904 39908 64950
rect 39985 64904 40031 64950
rect 40108 64904 40154 64950
rect 43739 64904 43785 64950
rect 43906 64904 43952 64950
rect 44071 64904 44117 64950
rect 44236 64904 44282 64950
rect 33684 64680 33730 64726
rect 33787 64680 33833 64726
rect 33890 64680 33936 64726
rect 33993 64680 34039 64726
rect 34096 64680 34142 64726
rect 34199 64680 34245 64726
rect 34302 64680 34348 64726
rect 34405 64680 34451 64726
rect 34508 64680 34554 64726
rect 34612 64680 34658 64726
rect 39740 64680 39786 64726
rect 39862 64680 39908 64726
rect 39985 64680 40031 64726
rect 40108 64680 40154 64726
rect 50467 64904 50513 64950
rect 50571 64904 50617 64950
rect 50674 64904 50720 64950
rect 50777 64904 50823 64950
rect 50880 64904 50926 64950
rect 50983 64904 51029 64950
rect 51086 64904 51132 64950
rect 51189 64904 51235 64950
rect 51292 64904 51338 64950
rect 51395 64904 51441 64950
rect 50467 64680 50513 64726
rect 50571 64680 50617 64726
rect 50674 64680 50720 64726
rect 50777 64680 50823 64726
rect 50880 64680 50926 64726
rect 50983 64680 51029 64726
rect 51086 64680 51132 64726
rect 51189 64680 51235 64726
rect 51292 64680 51338 64726
rect 51395 64680 51441 64726
rect 37909 64593 37955 64639
rect 38026 64593 38072 64639
rect 38143 64593 38189 64639
rect 38261 64593 38307 64639
rect 38379 64593 38425 64639
rect 38497 64593 38543 64639
rect 33684 64456 33730 64502
rect 33787 64456 33833 64502
rect 33890 64456 33936 64502
rect 33993 64456 34039 64502
rect 34096 64456 34142 64502
rect 34199 64456 34245 64502
rect 34302 64456 34348 64502
rect 34405 64456 34451 64502
rect 34508 64456 34554 64502
rect 34612 64456 34658 64502
rect 33816 64197 33862 64243
rect 34002 64197 34048 64243
rect 34189 64197 34235 64243
rect 34376 64197 34422 64243
rect 34562 64197 34608 64243
rect 37909 64369 37955 64415
rect 38026 64369 38072 64415
rect 38143 64369 38189 64415
rect 38261 64369 38307 64415
rect 38379 64369 38425 64415
rect 38497 64369 38543 64415
rect 39641 64369 39687 64415
rect 50467 64456 50513 64502
rect 50571 64456 50617 64502
rect 50674 64456 50720 64502
rect 50777 64456 50823 64502
rect 50880 64456 50926 64502
rect 50983 64456 51029 64502
rect 51086 64456 51132 64502
rect 51189 64456 51235 64502
rect 51292 64456 51338 64502
rect 51395 64456 51441 64502
rect 37909 64145 37955 64191
rect 38026 64145 38072 64191
rect 38143 64145 38189 64191
rect 38261 64145 38307 64191
rect 38379 64145 38425 64191
rect 38497 64145 38543 64191
rect 39641 64145 39687 64191
rect 43739 64211 43785 64257
rect 43906 64211 43952 64257
rect 44071 64211 44117 64257
rect 44236 64211 44282 64257
rect 50516 64197 50562 64243
rect 50703 64197 50749 64243
rect 50890 64197 50936 64243
rect 51076 64197 51122 64243
rect 51263 64197 51309 64243
rect 33816 63811 33862 63857
rect 34002 63811 34048 63857
rect 34189 63811 34235 63857
rect 34376 63811 34422 63857
rect 34562 63811 34608 63857
rect 37909 63863 37955 63909
rect 38026 63863 38072 63909
rect 38143 63863 38189 63909
rect 38261 63863 38307 63909
rect 38379 63863 38425 63909
rect 38497 63863 38543 63909
rect 39641 63863 39687 63909
rect 33684 63552 33730 63598
rect 33787 63552 33833 63598
rect 33890 63552 33936 63598
rect 33993 63552 34039 63598
rect 34096 63552 34142 63598
rect 34199 63552 34245 63598
rect 34302 63552 34348 63598
rect 34405 63552 34451 63598
rect 34508 63552 34554 63598
rect 34612 63552 34658 63598
rect 37909 63639 37955 63685
rect 38026 63639 38072 63685
rect 38143 63639 38189 63685
rect 38261 63639 38307 63685
rect 38379 63639 38425 63685
rect 38497 63639 38543 63685
rect 43739 63797 43785 63843
rect 43906 63797 43952 63843
rect 44071 63797 44117 63843
rect 44236 63797 44282 63843
rect 39641 63639 39687 63685
rect 50516 63811 50562 63857
rect 50703 63811 50749 63857
rect 50890 63811 50936 63857
rect 51076 63811 51122 63857
rect 51263 63811 51309 63857
rect 37909 63415 37955 63461
rect 38026 63415 38072 63461
rect 38143 63415 38189 63461
rect 38261 63415 38307 63461
rect 38379 63415 38425 63461
rect 38497 63415 38543 63461
rect 50467 63552 50513 63598
rect 50571 63552 50617 63598
rect 50674 63552 50720 63598
rect 50777 63552 50823 63598
rect 50880 63552 50926 63598
rect 50983 63552 51029 63598
rect 51086 63552 51132 63598
rect 51189 63552 51235 63598
rect 51292 63552 51338 63598
rect 51395 63552 51441 63598
rect 33684 63328 33730 63374
rect 33787 63328 33833 63374
rect 33890 63328 33936 63374
rect 33993 63328 34039 63374
rect 34096 63328 34142 63374
rect 34199 63328 34245 63374
rect 34302 63328 34348 63374
rect 34405 63328 34451 63374
rect 34508 63328 34554 63374
rect 34612 63328 34658 63374
rect 39740 63328 39786 63374
rect 39862 63328 39908 63374
rect 39985 63328 40031 63374
rect 40108 63328 40154 63374
rect 33684 63104 33730 63150
rect 33787 63104 33833 63150
rect 33890 63104 33936 63150
rect 33993 63104 34039 63150
rect 34096 63104 34142 63150
rect 34199 63104 34245 63150
rect 34302 63104 34348 63150
rect 34405 63104 34451 63150
rect 34508 63104 34554 63150
rect 34612 63104 34658 63150
rect 39740 63104 39786 63150
rect 39862 63104 39908 63150
rect 39985 63104 40031 63150
rect 40108 63104 40154 63150
rect 50467 63328 50513 63374
rect 50571 63328 50617 63374
rect 50674 63328 50720 63374
rect 50777 63328 50823 63374
rect 50880 63328 50926 63374
rect 50983 63328 51029 63374
rect 51086 63328 51132 63374
rect 51189 63328 51235 63374
rect 51292 63328 51338 63374
rect 51395 63328 51441 63374
rect 43739 63104 43785 63150
rect 43906 63104 43952 63150
rect 44071 63104 44117 63150
rect 44236 63104 44282 63150
rect 33684 62880 33730 62926
rect 33787 62880 33833 62926
rect 33890 62880 33936 62926
rect 33993 62880 34039 62926
rect 34096 62880 34142 62926
rect 34199 62880 34245 62926
rect 34302 62880 34348 62926
rect 34405 62880 34451 62926
rect 34508 62880 34554 62926
rect 34612 62880 34658 62926
rect 39740 62880 39786 62926
rect 39862 62880 39908 62926
rect 39985 62880 40031 62926
rect 40108 62880 40154 62926
rect 50467 63104 50513 63150
rect 50571 63104 50617 63150
rect 50674 63104 50720 63150
rect 50777 63104 50823 63150
rect 50880 63104 50926 63150
rect 50983 63104 51029 63150
rect 51086 63104 51132 63150
rect 51189 63104 51235 63150
rect 51292 63104 51338 63150
rect 51395 63104 51441 63150
rect 50467 62880 50513 62926
rect 50571 62880 50617 62926
rect 50674 62880 50720 62926
rect 50777 62880 50823 62926
rect 50880 62880 50926 62926
rect 50983 62880 51029 62926
rect 51086 62880 51132 62926
rect 51189 62880 51235 62926
rect 51292 62880 51338 62926
rect 51395 62880 51441 62926
rect 37909 62793 37955 62839
rect 38026 62793 38072 62839
rect 38143 62793 38189 62839
rect 38261 62793 38307 62839
rect 38379 62793 38425 62839
rect 38497 62793 38543 62839
rect 33684 62656 33730 62702
rect 33787 62656 33833 62702
rect 33890 62656 33936 62702
rect 33993 62656 34039 62702
rect 34096 62656 34142 62702
rect 34199 62656 34245 62702
rect 34302 62656 34348 62702
rect 34405 62656 34451 62702
rect 34508 62656 34554 62702
rect 34612 62656 34658 62702
rect 33816 62397 33862 62443
rect 34002 62397 34048 62443
rect 34189 62397 34235 62443
rect 34376 62397 34422 62443
rect 34562 62397 34608 62443
rect 37909 62569 37955 62615
rect 38026 62569 38072 62615
rect 38143 62569 38189 62615
rect 38261 62569 38307 62615
rect 38379 62569 38425 62615
rect 38497 62569 38543 62615
rect 39641 62569 39687 62615
rect 50467 62656 50513 62702
rect 50571 62656 50617 62702
rect 50674 62656 50720 62702
rect 50777 62656 50823 62702
rect 50880 62656 50926 62702
rect 50983 62656 51029 62702
rect 51086 62656 51132 62702
rect 51189 62656 51235 62702
rect 51292 62656 51338 62702
rect 51395 62656 51441 62702
rect 37909 62345 37955 62391
rect 38026 62345 38072 62391
rect 38143 62345 38189 62391
rect 38261 62345 38307 62391
rect 38379 62345 38425 62391
rect 38497 62345 38543 62391
rect 39641 62345 39687 62391
rect 43739 62411 43785 62457
rect 43906 62411 43952 62457
rect 44071 62411 44117 62457
rect 44236 62411 44282 62457
rect 50516 62397 50562 62443
rect 50703 62397 50749 62443
rect 50890 62397 50936 62443
rect 51076 62397 51122 62443
rect 51263 62397 51309 62443
rect 33816 62011 33862 62057
rect 34002 62011 34048 62057
rect 34189 62011 34235 62057
rect 34376 62011 34422 62057
rect 34562 62011 34608 62057
rect 37909 62063 37955 62109
rect 38026 62063 38072 62109
rect 38143 62063 38189 62109
rect 38261 62063 38307 62109
rect 38379 62063 38425 62109
rect 38497 62063 38543 62109
rect 39641 62063 39687 62109
rect 33684 61752 33730 61798
rect 33787 61752 33833 61798
rect 33890 61752 33936 61798
rect 33993 61752 34039 61798
rect 34096 61752 34142 61798
rect 34199 61752 34245 61798
rect 34302 61752 34348 61798
rect 34405 61752 34451 61798
rect 34508 61752 34554 61798
rect 34612 61752 34658 61798
rect 37909 61839 37955 61885
rect 38026 61839 38072 61885
rect 38143 61839 38189 61885
rect 38261 61839 38307 61885
rect 38379 61839 38425 61885
rect 38497 61839 38543 61885
rect 43739 61997 43785 62043
rect 43906 61997 43952 62043
rect 44071 61997 44117 62043
rect 44236 61997 44282 62043
rect 39641 61839 39687 61885
rect 50516 62011 50562 62057
rect 50703 62011 50749 62057
rect 50890 62011 50936 62057
rect 51076 62011 51122 62057
rect 51263 62011 51309 62057
rect 37909 61615 37955 61661
rect 38026 61615 38072 61661
rect 38143 61615 38189 61661
rect 38261 61615 38307 61661
rect 38379 61615 38425 61661
rect 38497 61615 38543 61661
rect 50467 61752 50513 61798
rect 50571 61752 50617 61798
rect 50674 61752 50720 61798
rect 50777 61752 50823 61798
rect 50880 61752 50926 61798
rect 50983 61752 51029 61798
rect 51086 61752 51132 61798
rect 51189 61752 51235 61798
rect 51292 61752 51338 61798
rect 51395 61752 51441 61798
rect 33684 61528 33730 61574
rect 33787 61528 33833 61574
rect 33890 61528 33936 61574
rect 33993 61528 34039 61574
rect 34096 61528 34142 61574
rect 34199 61528 34245 61574
rect 34302 61528 34348 61574
rect 34405 61528 34451 61574
rect 34508 61528 34554 61574
rect 34612 61528 34658 61574
rect 39740 61528 39786 61574
rect 39862 61528 39908 61574
rect 39985 61528 40031 61574
rect 40108 61528 40154 61574
rect 33684 61304 33730 61350
rect 33787 61304 33833 61350
rect 33890 61304 33936 61350
rect 33993 61304 34039 61350
rect 34096 61304 34142 61350
rect 34199 61304 34245 61350
rect 34302 61304 34348 61350
rect 34405 61304 34451 61350
rect 34508 61304 34554 61350
rect 34612 61304 34658 61350
rect 39740 61304 39786 61350
rect 39862 61304 39908 61350
rect 39985 61304 40031 61350
rect 40108 61304 40154 61350
rect 50467 61528 50513 61574
rect 50571 61528 50617 61574
rect 50674 61528 50720 61574
rect 50777 61528 50823 61574
rect 50880 61528 50926 61574
rect 50983 61528 51029 61574
rect 51086 61528 51132 61574
rect 51189 61528 51235 61574
rect 51292 61528 51338 61574
rect 51395 61528 51441 61574
rect 43739 61304 43785 61350
rect 43906 61304 43952 61350
rect 44071 61304 44117 61350
rect 44236 61304 44282 61350
rect 33684 61080 33730 61126
rect 33787 61080 33833 61126
rect 33890 61080 33936 61126
rect 33993 61080 34039 61126
rect 34096 61080 34142 61126
rect 34199 61080 34245 61126
rect 34302 61080 34348 61126
rect 34405 61080 34451 61126
rect 34508 61080 34554 61126
rect 34612 61080 34658 61126
rect 39740 61080 39786 61126
rect 39862 61080 39908 61126
rect 39985 61080 40031 61126
rect 40108 61080 40154 61126
rect 50467 61304 50513 61350
rect 50571 61304 50617 61350
rect 50674 61304 50720 61350
rect 50777 61304 50823 61350
rect 50880 61304 50926 61350
rect 50983 61304 51029 61350
rect 51086 61304 51132 61350
rect 51189 61304 51235 61350
rect 51292 61304 51338 61350
rect 51395 61304 51441 61350
rect 50467 61080 50513 61126
rect 50571 61080 50617 61126
rect 50674 61080 50720 61126
rect 50777 61080 50823 61126
rect 50880 61080 50926 61126
rect 50983 61080 51029 61126
rect 51086 61080 51132 61126
rect 51189 61080 51235 61126
rect 51292 61080 51338 61126
rect 51395 61080 51441 61126
rect 37909 60993 37955 61039
rect 38026 60993 38072 61039
rect 38143 60993 38189 61039
rect 38261 60993 38307 61039
rect 38379 60993 38425 61039
rect 38497 60993 38543 61039
rect 33684 60856 33730 60902
rect 33787 60856 33833 60902
rect 33890 60856 33936 60902
rect 33993 60856 34039 60902
rect 34096 60856 34142 60902
rect 34199 60856 34245 60902
rect 34302 60856 34348 60902
rect 34405 60856 34451 60902
rect 34508 60856 34554 60902
rect 34612 60856 34658 60902
rect 33816 60597 33862 60643
rect 34002 60597 34048 60643
rect 34189 60597 34235 60643
rect 34376 60597 34422 60643
rect 34562 60597 34608 60643
rect 37909 60769 37955 60815
rect 38026 60769 38072 60815
rect 38143 60769 38189 60815
rect 38261 60769 38307 60815
rect 38379 60769 38425 60815
rect 38497 60769 38543 60815
rect 39641 60769 39687 60815
rect 50467 60856 50513 60902
rect 50571 60856 50617 60902
rect 50674 60856 50720 60902
rect 50777 60856 50823 60902
rect 50880 60856 50926 60902
rect 50983 60856 51029 60902
rect 51086 60856 51132 60902
rect 51189 60856 51235 60902
rect 51292 60856 51338 60902
rect 51395 60856 51441 60902
rect 37909 60545 37955 60591
rect 38026 60545 38072 60591
rect 38143 60545 38189 60591
rect 38261 60545 38307 60591
rect 38379 60545 38425 60591
rect 38497 60545 38543 60591
rect 39641 60545 39687 60591
rect 43739 60611 43785 60657
rect 43906 60611 43952 60657
rect 44071 60611 44117 60657
rect 44236 60611 44282 60657
rect 50516 60597 50562 60643
rect 50703 60597 50749 60643
rect 50890 60597 50936 60643
rect 51076 60597 51122 60643
rect 51263 60597 51309 60643
rect 33816 60211 33862 60257
rect 34002 60211 34048 60257
rect 34189 60211 34235 60257
rect 34376 60211 34422 60257
rect 34562 60211 34608 60257
rect 37909 60263 37955 60309
rect 38026 60263 38072 60309
rect 38143 60263 38189 60309
rect 38261 60263 38307 60309
rect 38379 60263 38425 60309
rect 38497 60263 38543 60309
rect 39641 60263 39687 60309
rect 33684 59952 33730 59998
rect 33787 59952 33833 59998
rect 33890 59952 33936 59998
rect 33993 59952 34039 59998
rect 34096 59952 34142 59998
rect 34199 59952 34245 59998
rect 34302 59952 34348 59998
rect 34405 59952 34451 59998
rect 34508 59952 34554 59998
rect 34612 59952 34658 59998
rect 37909 60039 37955 60085
rect 38026 60039 38072 60085
rect 38143 60039 38189 60085
rect 38261 60039 38307 60085
rect 38379 60039 38425 60085
rect 38497 60039 38543 60085
rect 43739 60197 43785 60243
rect 43906 60197 43952 60243
rect 44071 60197 44117 60243
rect 44236 60197 44282 60243
rect 39641 60039 39687 60085
rect 50516 60211 50562 60257
rect 50703 60211 50749 60257
rect 50890 60211 50936 60257
rect 51076 60211 51122 60257
rect 51263 60211 51309 60257
rect 37909 59815 37955 59861
rect 38026 59815 38072 59861
rect 38143 59815 38189 59861
rect 38261 59815 38307 59861
rect 38379 59815 38425 59861
rect 38497 59815 38543 59861
rect 50467 59952 50513 59998
rect 50571 59952 50617 59998
rect 50674 59952 50720 59998
rect 50777 59952 50823 59998
rect 50880 59952 50926 59998
rect 50983 59952 51029 59998
rect 51086 59952 51132 59998
rect 51189 59952 51235 59998
rect 51292 59952 51338 59998
rect 51395 59952 51441 59998
rect 33684 59728 33730 59774
rect 33787 59728 33833 59774
rect 33890 59728 33936 59774
rect 33993 59728 34039 59774
rect 34096 59728 34142 59774
rect 34199 59728 34245 59774
rect 34302 59728 34348 59774
rect 34405 59728 34451 59774
rect 34508 59728 34554 59774
rect 34612 59728 34658 59774
rect 39740 59728 39786 59774
rect 39862 59728 39908 59774
rect 39985 59728 40031 59774
rect 40108 59728 40154 59774
rect 33684 59504 33730 59550
rect 33787 59504 33833 59550
rect 33890 59504 33936 59550
rect 33993 59504 34039 59550
rect 34096 59504 34142 59550
rect 34199 59504 34245 59550
rect 34302 59504 34348 59550
rect 34405 59504 34451 59550
rect 34508 59504 34554 59550
rect 34612 59504 34658 59550
rect 39740 59504 39786 59550
rect 39862 59504 39908 59550
rect 39985 59504 40031 59550
rect 40108 59504 40154 59550
rect 50467 59728 50513 59774
rect 50571 59728 50617 59774
rect 50674 59728 50720 59774
rect 50777 59728 50823 59774
rect 50880 59728 50926 59774
rect 50983 59728 51029 59774
rect 51086 59728 51132 59774
rect 51189 59728 51235 59774
rect 51292 59728 51338 59774
rect 51395 59728 51441 59774
rect 43739 59504 43785 59550
rect 43906 59504 43952 59550
rect 44071 59504 44117 59550
rect 44236 59504 44282 59550
rect 33684 59280 33730 59326
rect 33787 59280 33833 59326
rect 33890 59280 33936 59326
rect 33993 59280 34039 59326
rect 34096 59280 34142 59326
rect 34199 59280 34245 59326
rect 34302 59280 34348 59326
rect 34405 59280 34451 59326
rect 34508 59280 34554 59326
rect 34612 59280 34658 59326
rect 39740 59280 39786 59326
rect 39862 59280 39908 59326
rect 39985 59280 40031 59326
rect 40108 59280 40154 59326
rect 50467 59504 50513 59550
rect 50571 59504 50617 59550
rect 50674 59504 50720 59550
rect 50777 59504 50823 59550
rect 50880 59504 50926 59550
rect 50983 59504 51029 59550
rect 51086 59504 51132 59550
rect 51189 59504 51235 59550
rect 51292 59504 51338 59550
rect 51395 59504 51441 59550
rect 50467 59280 50513 59326
rect 50571 59280 50617 59326
rect 50674 59280 50720 59326
rect 50777 59280 50823 59326
rect 50880 59280 50926 59326
rect 50983 59280 51029 59326
rect 51086 59280 51132 59326
rect 51189 59280 51235 59326
rect 51292 59280 51338 59326
rect 51395 59280 51441 59326
rect 37909 59193 37955 59239
rect 38026 59193 38072 59239
rect 38143 59193 38189 59239
rect 38261 59193 38307 59239
rect 38379 59193 38425 59239
rect 38497 59193 38543 59239
rect 33684 59056 33730 59102
rect 33787 59056 33833 59102
rect 33890 59056 33936 59102
rect 33993 59056 34039 59102
rect 34096 59056 34142 59102
rect 34199 59056 34245 59102
rect 34302 59056 34348 59102
rect 34405 59056 34451 59102
rect 34508 59056 34554 59102
rect 34612 59056 34658 59102
rect 33816 58797 33862 58843
rect 34002 58797 34048 58843
rect 34189 58797 34235 58843
rect 34376 58797 34422 58843
rect 34562 58797 34608 58843
rect 37909 58969 37955 59015
rect 38026 58969 38072 59015
rect 38143 58969 38189 59015
rect 38261 58969 38307 59015
rect 38379 58969 38425 59015
rect 38497 58969 38543 59015
rect 39641 58969 39687 59015
rect 50467 59056 50513 59102
rect 50571 59056 50617 59102
rect 50674 59056 50720 59102
rect 50777 59056 50823 59102
rect 50880 59056 50926 59102
rect 50983 59056 51029 59102
rect 51086 59056 51132 59102
rect 51189 59056 51235 59102
rect 51292 59056 51338 59102
rect 51395 59056 51441 59102
rect 37909 58745 37955 58791
rect 38026 58745 38072 58791
rect 38143 58745 38189 58791
rect 38261 58745 38307 58791
rect 38379 58745 38425 58791
rect 38497 58745 38543 58791
rect 39641 58745 39687 58791
rect 43739 58811 43785 58857
rect 43906 58811 43952 58857
rect 44071 58811 44117 58857
rect 44236 58811 44282 58857
rect 50516 58797 50562 58843
rect 50703 58797 50749 58843
rect 50890 58797 50936 58843
rect 51076 58797 51122 58843
rect 51263 58797 51309 58843
rect 33816 58411 33862 58457
rect 34002 58411 34048 58457
rect 34189 58411 34235 58457
rect 34376 58411 34422 58457
rect 34562 58411 34608 58457
rect 37909 58463 37955 58509
rect 38026 58463 38072 58509
rect 38143 58463 38189 58509
rect 38261 58463 38307 58509
rect 38379 58463 38425 58509
rect 38497 58463 38543 58509
rect 39641 58463 39687 58509
rect 33684 58152 33730 58198
rect 33787 58152 33833 58198
rect 33890 58152 33936 58198
rect 33993 58152 34039 58198
rect 34096 58152 34142 58198
rect 34199 58152 34245 58198
rect 34302 58152 34348 58198
rect 34405 58152 34451 58198
rect 34508 58152 34554 58198
rect 34612 58152 34658 58198
rect 37909 58239 37955 58285
rect 38026 58239 38072 58285
rect 38143 58239 38189 58285
rect 38261 58239 38307 58285
rect 38379 58239 38425 58285
rect 38497 58239 38543 58285
rect 43739 58397 43785 58443
rect 43906 58397 43952 58443
rect 44071 58397 44117 58443
rect 44236 58397 44282 58443
rect 39641 58239 39687 58285
rect 50516 58411 50562 58457
rect 50703 58411 50749 58457
rect 50890 58411 50936 58457
rect 51076 58411 51122 58457
rect 51263 58411 51309 58457
rect 37909 58015 37955 58061
rect 38026 58015 38072 58061
rect 38143 58015 38189 58061
rect 38261 58015 38307 58061
rect 38379 58015 38425 58061
rect 38497 58015 38543 58061
rect 50467 58152 50513 58198
rect 50571 58152 50617 58198
rect 50674 58152 50720 58198
rect 50777 58152 50823 58198
rect 50880 58152 50926 58198
rect 50983 58152 51029 58198
rect 51086 58152 51132 58198
rect 51189 58152 51235 58198
rect 51292 58152 51338 58198
rect 51395 58152 51441 58198
rect 33684 57928 33730 57974
rect 33787 57928 33833 57974
rect 33890 57928 33936 57974
rect 33993 57928 34039 57974
rect 34096 57928 34142 57974
rect 34199 57928 34245 57974
rect 34302 57928 34348 57974
rect 34405 57928 34451 57974
rect 34508 57928 34554 57974
rect 34612 57928 34658 57974
rect 39740 57928 39786 57974
rect 39862 57928 39908 57974
rect 39985 57928 40031 57974
rect 40108 57928 40154 57974
rect 33684 57704 33730 57750
rect 33787 57704 33833 57750
rect 33890 57704 33936 57750
rect 33993 57704 34039 57750
rect 34096 57704 34142 57750
rect 34199 57704 34245 57750
rect 34302 57704 34348 57750
rect 34405 57704 34451 57750
rect 34508 57704 34554 57750
rect 34612 57704 34658 57750
rect 39740 57704 39786 57750
rect 39862 57704 39908 57750
rect 39985 57704 40031 57750
rect 40108 57704 40154 57750
rect 50467 57928 50513 57974
rect 50571 57928 50617 57974
rect 50674 57928 50720 57974
rect 50777 57928 50823 57974
rect 50880 57928 50926 57974
rect 50983 57928 51029 57974
rect 51086 57928 51132 57974
rect 51189 57928 51235 57974
rect 51292 57928 51338 57974
rect 51395 57928 51441 57974
rect 43739 57704 43785 57750
rect 43906 57704 43952 57750
rect 44071 57704 44117 57750
rect 44236 57704 44282 57750
rect 33684 57480 33730 57526
rect 33787 57480 33833 57526
rect 33890 57480 33936 57526
rect 33993 57480 34039 57526
rect 34096 57480 34142 57526
rect 34199 57480 34245 57526
rect 34302 57480 34348 57526
rect 34405 57480 34451 57526
rect 34508 57480 34554 57526
rect 34612 57480 34658 57526
rect 39740 57480 39786 57526
rect 39862 57480 39908 57526
rect 39985 57480 40031 57526
rect 40108 57480 40154 57526
rect 50467 57704 50513 57750
rect 50571 57704 50617 57750
rect 50674 57704 50720 57750
rect 50777 57704 50823 57750
rect 50880 57704 50926 57750
rect 50983 57704 51029 57750
rect 51086 57704 51132 57750
rect 51189 57704 51235 57750
rect 51292 57704 51338 57750
rect 51395 57704 51441 57750
rect 50467 57480 50513 57526
rect 50571 57480 50617 57526
rect 50674 57480 50720 57526
rect 50777 57480 50823 57526
rect 50880 57480 50926 57526
rect 50983 57480 51029 57526
rect 51086 57480 51132 57526
rect 51189 57480 51235 57526
rect 51292 57480 51338 57526
rect 51395 57480 51441 57526
rect 37909 57393 37955 57439
rect 38026 57393 38072 57439
rect 38143 57393 38189 57439
rect 38261 57393 38307 57439
rect 38379 57393 38425 57439
rect 38497 57393 38543 57439
rect 33684 57256 33730 57302
rect 33787 57256 33833 57302
rect 33890 57256 33936 57302
rect 33993 57256 34039 57302
rect 34096 57256 34142 57302
rect 34199 57256 34245 57302
rect 34302 57256 34348 57302
rect 34405 57256 34451 57302
rect 34508 57256 34554 57302
rect 34612 57256 34658 57302
rect 33816 56997 33862 57043
rect 34002 56997 34048 57043
rect 34189 56997 34235 57043
rect 34376 56997 34422 57043
rect 34562 56997 34608 57043
rect 37909 57169 37955 57215
rect 38026 57169 38072 57215
rect 38143 57169 38189 57215
rect 38261 57169 38307 57215
rect 38379 57169 38425 57215
rect 38497 57169 38543 57215
rect 39641 57169 39687 57215
rect 50467 57256 50513 57302
rect 50571 57256 50617 57302
rect 50674 57256 50720 57302
rect 50777 57256 50823 57302
rect 50880 57256 50926 57302
rect 50983 57256 51029 57302
rect 51086 57256 51132 57302
rect 51189 57256 51235 57302
rect 51292 57256 51338 57302
rect 51395 57256 51441 57302
rect 37909 56945 37955 56991
rect 38026 56945 38072 56991
rect 38143 56945 38189 56991
rect 38261 56945 38307 56991
rect 38379 56945 38425 56991
rect 38497 56945 38543 56991
rect 39641 56945 39687 56991
rect 43739 57011 43785 57057
rect 43906 57011 43952 57057
rect 44071 57011 44117 57057
rect 44236 57011 44282 57057
rect 50516 56997 50562 57043
rect 50703 56997 50749 57043
rect 50890 56997 50936 57043
rect 51076 56997 51122 57043
rect 51263 56997 51309 57043
rect 33816 56611 33862 56657
rect 34002 56611 34048 56657
rect 34189 56611 34235 56657
rect 34376 56611 34422 56657
rect 34562 56611 34608 56657
rect 37909 56663 37955 56709
rect 38026 56663 38072 56709
rect 38143 56663 38189 56709
rect 38261 56663 38307 56709
rect 38379 56663 38425 56709
rect 38497 56663 38543 56709
rect 39641 56663 39687 56709
rect 33684 56352 33730 56398
rect 33787 56352 33833 56398
rect 33890 56352 33936 56398
rect 33993 56352 34039 56398
rect 34096 56352 34142 56398
rect 34199 56352 34245 56398
rect 34302 56352 34348 56398
rect 34405 56352 34451 56398
rect 34508 56352 34554 56398
rect 34612 56352 34658 56398
rect 37909 56439 37955 56485
rect 38026 56439 38072 56485
rect 38143 56439 38189 56485
rect 38261 56439 38307 56485
rect 38379 56439 38425 56485
rect 38497 56439 38543 56485
rect 43739 56597 43785 56643
rect 43906 56597 43952 56643
rect 44071 56597 44117 56643
rect 44236 56597 44282 56643
rect 39641 56439 39687 56485
rect 50516 56611 50562 56657
rect 50703 56611 50749 56657
rect 50890 56611 50936 56657
rect 51076 56611 51122 56657
rect 51263 56611 51309 56657
rect 37909 56215 37955 56261
rect 38026 56215 38072 56261
rect 38143 56215 38189 56261
rect 38261 56215 38307 56261
rect 38379 56215 38425 56261
rect 38497 56215 38543 56261
rect 50467 56352 50513 56398
rect 50571 56352 50617 56398
rect 50674 56352 50720 56398
rect 50777 56352 50823 56398
rect 50880 56352 50926 56398
rect 50983 56352 51029 56398
rect 51086 56352 51132 56398
rect 51189 56352 51235 56398
rect 51292 56352 51338 56398
rect 51395 56352 51441 56398
rect 33684 56128 33730 56174
rect 33787 56128 33833 56174
rect 33890 56128 33936 56174
rect 33993 56128 34039 56174
rect 34096 56128 34142 56174
rect 34199 56128 34245 56174
rect 34302 56128 34348 56174
rect 34405 56128 34451 56174
rect 34508 56128 34554 56174
rect 34612 56128 34658 56174
rect 39740 56128 39786 56174
rect 39862 56128 39908 56174
rect 39985 56128 40031 56174
rect 40108 56128 40154 56174
rect 33684 55904 33730 55950
rect 33787 55904 33833 55950
rect 33890 55904 33936 55950
rect 33993 55904 34039 55950
rect 34096 55904 34142 55950
rect 34199 55904 34245 55950
rect 34302 55904 34348 55950
rect 34405 55904 34451 55950
rect 34508 55904 34554 55950
rect 34612 55904 34658 55950
rect 39740 55904 39786 55950
rect 39862 55904 39908 55950
rect 39985 55904 40031 55950
rect 40108 55904 40154 55950
rect 50467 56128 50513 56174
rect 50571 56128 50617 56174
rect 50674 56128 50720 56174
rect 50777 56128 50823 56174
rect 50880 56128 50926 56174
rect 50983 56128 51029 56174
rect 51086 56128 51132 56174
rect 51189 56128 51235 56174
rect 51292 56128 51338 56174
rect 51395 56128 51441 56174
rect 43739 55904 43785 55950
rect 43906 55904 43952 55950
rect 44071 55904 44117 55950
rect 44236 55904 44282 55950
rect 33684 55680 33730 55726
rect 33787 55680 33833 55726
rect 33890 55680 33936 55726
rect 33993 55680 34039 55726
rect 34096 55680 34142 55726
rect 34199 55680 34245 55726
rect 34302 55680 34348 55726
rect 34405 55680 34451 55726
rect 34508 55680 34554 55726
rect 34612 55680 34658 55726
rect 39740 55680 39786 55726
rect 39862 55680 39908 55726
rect 39985 55680 40031 55726
rect 40108 55680 40154 55726
rect 50467 55904 50513 55950
rect 50571 55904 50617 55950
rect 50674 55904 50720 55950
rect 50777 55904 50823 55950
rect 50880 55904 50926 55950
rect 50983 55904 51029 55950
rect 51086 55904 51132 55950
rect 51189 55904 51235 55950
rect 51292 55904 51338 55950
rect 51395 55904 51441 55950
rect 50467 55680 50513 55726
rect 50571 55680 50617 55726
rect 50674 55680 50720 55726
rect 50777 55680 50823 55726
rect 50880 55680 50926 55726
rect 50983 55680 51029 55726
rect 51086 55680 51132 55726
rect 51189 55680 51235 55726
rect 51292 55680 51338 55726
rect 51395 55680 51441 55726
rect 37909 55593 37955 55639
rect 38026 55593 38072 55639
rect 38143 55593 38189 55639
rect 38261 55593 38307 55639
rect 38379 55593 38425 55639
rect 38497 55593 38543 55639
rect 33684 55456 33730 55502
rect 33787 55456 33833 55502
rect 33890 55456 33936 55502
rect 33993 55456 34039 55502
rect 34096 55456 34142 55502
rect 34199 55456 34245 55502
rect 34302 55456 34348 55502
rect 34405 55456 34451 55502
rect 34508 55456 34554 55502
rect 34612 55456 34658 55502
rect 33816 55197 33862 55243
rect 34002 55197 34048 55243
rect 34189 55197 34235 55243
rect 34376 55197 34422 55243
rect 34562 55197 34608 55243
rect 37909 55369 37955 55415
rect 38026 55369 38072 55415
rect 38143 55369 38189 55415
rect 38261 55369 38307 55415
rect 38379 55369 38425 55415
rect 38497 55369 38543 55415
rect 39641 55369 39687 55415
rect 50467 55456 50513 55502
rect 50571 55456 50617 55502
rect 50674 55456 50720 55502
rect 50777 55456 50823 55502
rect 50880 55456 50926 55502
rect 50983 55456 51029 55502
rect 51086 55456 51132 55502
rect 51189 55456 51235 55502
rect 51292 55456 51338 55502
rect 51395 55456 51441 55502
rect 37909 55145 37955 55191
rect 38026 55145 38072 55191
rect 38143 55145 38189 55191
rect 38261 55145 38307 55191
rect 38379 55145 38425 55191
rect 38497 55145 38543 55191
rect 39641 55145 39687 55191
rect 43739 55211 43785 55257
rect 43906 55211 43952 55257
rect 44071 55211 44117 55257
rect 44236 55211 44282 55257
rect 50516 55197 50562 55243
rect 50703 55197 50749 55243
rect 50890 55197 50936 55243
rect 51076 55197 51122 55243
rect 51263 55197 51309 55243
rect 33816 54811 33862 54857
rect 34002 54811 34048 54857
rect 34189 54811 34235 54857
rect 34376 54811 34422 54857
rect 34562 54811 34608 54857
rect 37909 54863 37955 54909
rect 38026 54863 38072 54909
rect 38143 54863 38189 54909
rect 38261 54863 38307 54909
rect 38379 54863 38425 54909
rect 38497 54863 38543 54909
rect 39641 54863 39687 54909
rect 33684 54552 33730 54598
rect 33787 54552 33833 54598
rect 33890 54552 33936 54598
rect 33993 54552 34039 54598
rect 34096 54552 34142 54598
rect 34199 54552 34245 54598
rect 34302 54552 34348 54598
rect 34405 54552 34451 54598
rect 34508 54552 34554 54598
rect 34612 54552 34658 54598
rect 37909 54639 37955 54685
rect 38026 54639 38072 54685
rect 38143 54639 38189 54685
rect 38261 54639 38307 54685
rect 38379 54639 38425 54685
rect 38497 54639 38543 54685
rect 43739 54797 43785 54843
rect 43906 54797 43952 54843
rect 44071 54797 44117 54843
rect 44236 54797 44282 54843
rect 39641 54639 39687 54685
rect 50516 54811 50562 54857
rect 50703 54811 50749 54857
rect 50890 54811 50936 54857
rect 51076 54811 51122 54857
rect 51263 54811 51309 54857
rect 37909 54415 37955 54461
rect 38026 54415 38072 54461
rect 38143 54415 38189 54461
rect 38261 54415 38307 54461
rect 38379 54415 38425 54461
rect 38497 54415 38543 54461
rect 50467 54552 50513 54598
rect 50571 54552 50617 54598
rect 50674 54552 50720 54598
rect 50777 54552 50823 54598
rect 50880 54552 50926 54598
rect 50983 54552 51029 54598
rect 51086 54552 51132 54598
rect 51189 54552 51235 54598
rect 51292 54552 51338 54598
rect 51395 54552 51441 54598
rect 33684 54328 33730 54374
rect 33787 54328 33833 54374
rect 33890 54328 33936 54374
rect 33993 54328 34039 54374
rect 34096 54328 34142 54374
rect 34199 54328 34245 54374
rect 34302 54328 34348 54374
rect 34405 54328 34451 54374
rect 34508 54328 34554 54374
rect 34612 54328 34658 54374
rect 39740 54328 39786 54374
rect 39862 54328 39908 54374
rect 39985 54328 40031 54374
rect 40108 54328 40154 54374
rect 33684 54104 33730 54150
rect 33787 54104 33833 54150
rect 33890 54104 33936 54150
rect 33993 54104 34039 54150
rect 34096 54104 34142 54150
rect 34199 54104 34245 54150
rect 34302 54104 34348 54150
rect 34405 54104 34451 54150
rect 34508 54104 34554 54150
rect 34612 54104 34658 54150
rect 39740 54104 39786 54150
rect 39862 54104 39908 54150
rect 39985 54104 40031 54150
rect 40108 54104 40154 54150
rect 50467 54328 50513 54374
rect 50571 54328 50617 54374
rect 50674 54328 50720 54374
rect 50777 54328 50823 54374
rect 50880 54328 50926 54374
rect 50983 54328 51029 54374
rect 51086 54328 51132 54374
rect 51189 54328 51235 54374
rect 51292 54328 51338 54374
rect 51395 54328 51441 54374
rect 43739 54104 43785 54150
rect 43906 54104 43952 54150
rect 44071 54104 44117 54150
rect 44236 54104 44282 54150
rect 33684 53880 33730 53926
rect 33787 53880 33833 53926
rect 33890 53880 33936 53926
rect 33993 53880 34039 53926
rect 34096 53880 34142 53926
rect 34199 53880 34245 53926
rect 34302 53880 34348 53926
rect 34405 53880 34451 53926
rect 34508 53880 34554 53926
rect 34612 53880 34658 53926
rect 39740 53880 39786 53926
rect 39862 53880 39908 53926
rect 39985 53880 40031 53926
rect 40108 53880 40154 53926
rect 50467 54104 50513 54150
rect 50571 54104 50617 54150
rect 50674 54104 50720 54150
rect 50777 54104 50823 54150
rect 50880 54104 50926 54150
rect 50983 54104 51029 54150
rect 51086 54104 51132 54150
rect 51189 54104 51235 54150
rect 51292 54104 51338 54150
rect 51395 54104 51441 54150
rect 50467 53880 50513 53926
rect 50571 53880 50617 53926
rect 50674 53880 50720 53926
rect 50777 53880 50823 53926
rect 50880 53880 50926 53926
rect 50983 53880 51029 53926
rect 51086 53880 51132 53926
rect 51189 53880 51235 53926
rect 51292 53880 51338 53926
rect 51395 53880 51441 53926
rect 37909 53793 37955 53839
rect 38026 53793 38072 53839
rect 38143 53793 38189 53839
rect 38261 53793 38307 53839
rect 38379 53793 38425 53839
rect 38497 53793 38543 53839
rect 33684 53656 33730 53702
rect 33787 53656 33833 53702
rect 33890 53656 33936 53702
rect 33993 53656 34039 53702
rect 34096 53656 34142 53702
rect 34199 53656 34245 53702
rect 34302 53656 34348 53702
rect 34405 53656 34451 53702
rect 34508 53656 34554 53702
rect 34612 53656 34658 53702
rect 33816 53397 33862 53443
rect 34002 53397 34048 53443
rect 34189 53397 34235 53443
rect 34376 53397 34422 53443
rect 34562 53397 34608 53443
rect 37909 53569 37955 53615
rect 38026 53569 38072 53615
rect 38143 53569 38189 53615
rect 38261 53569 38307 53615
rect 38379 53569 38425 53615
rect 38497 53569 38543 53615
rect 39641 53569 39687 53615
rect 50467 53656 50513 53702
rect 50571 53656 50617 53702
rect 50674 53656 50720 53702
rect 50777 53656 50823 53702
rect 50880 53656 50926 53702
rect 50983 53656 51029 53702
rect 51086 53656 51132 53702
rect 51189 53656 51235 53702
rect 51292 53656 51338 53702
rect 51395 53656 51441 53702
rect 37909 53345 37955 53391
rect 38026 53345 38072 53391
rect 38143 53345 38189 53391
rect 38261 53345 38307 53391
rect 38379 53345 38425 53391
rect 38497 53345 38543 53391
rect 39641 53345 39687 53391
rect 43739 53411 43785 53457
rect 43906 53411 43952 53457
rect 44071 53411 44117 53457
rect 44236 53411 44282 53457
rect 50516 53397 50562 53443
rect 50703 53397 50749 53443
rect 50890 53397 50936 53443
rect 51076 53397 51122 53443
rect 51263 53397 51309 53443
rect 33816 53011 33862 53057
rect 34002 53011 34048 53057
rect 34189 53011 34235 53057
rect 34376 53011 34422 53057
rect 34562 53011 34608 53057
rect 37909 53063 37955 53109
rect 38026 53063 38072 53109
rect 38143 53063 38189 53109
rect 38261 53063 38307 53109
rect 38379 53063 38425 53109
rect 38497 53063 38543 53109
rect 39641 53063 39687 53109
rect 33684 52752 33730 52798
rect 33787 52752 33833 52798
rect 33890 52752 33936 52798
rect 33993 52752 34039 52798
rect 34096 52752 34142 52798
rect 34199 52752 34245 52798
rect 34302 52752 34348 52798
rect 34405 52752 34451 52798
rect 34508 52752 34554 52798
rect 34612 52752 34658 52798
rect 37909 52839 37955 52885
rect 38026 52839 38072 52885
rect 38143 52839 38189 52885
rect 38261 52839 38307 52885
rect 38379 52839 38425 52885
rect 38497 52839 38543 52885
rect 43739 52997 43785 53043
rect 43906 52997 43952 53043
rect 44071 52997 44117 53043
rect 44236 52997 44282 53043
rect 39641 52839 39687 52885
rect 50516 53011 50562 53057
rect 50703 53011 50749 53057
rect 50890 53011 50936 53057
rect 51076 53011 51122 53057
rect 51263 53011 51309 53057
rect 37909 52615 37955 52661
rect 38026 52615 38072 52661
rect 38143 52615 38189 52661
rect 38261 52615 38307 52661
rect 38379 52615 38425 52661
rect 38497 52615 38543 52661
rect 50467 52752 50513 52798
rect 50571 52752 50617 52798
rect 50674 52752 50720 52798
rect 50777 52752 50823 52798
rect 50880 52752 50926 52798
rect 50983 52752 51029 52798
rect 51086 52752 51132 52798
rect 51189 52752 51235 52798
rect 51292 52752 51338 52798
rect 51395 52752 51441 52798
rect 33684 52528 33730 52574
rect 33787 52528 33833 52574
rect 33890 52528 33936 52574
rect 33993 52528 34039 52574
rect 34096 52528 34142 52574
rect 34199 52528 34245 52574
rect 34302 52528 34348 52574
rect 34405 52528 34451 52574
rect 34508 52528 34554 52574
rect 34612 52528 34658 52574
rect 39740 52528 39786 52574
rect 39862 52528 39908 52574
rect 39985 52528 40031 52574
rect 40108 52528 40154 52574
rect 33684 52304 33730 52350
rect 33787 52304 33833 52350
rect 33890 52304 33936 52350
rect 33993 52304 34039 52350
rect 34096 52304 34142 52350
rect 34199 52304 34245 52350
rect 34302 52304 34348 52350
rect 34405 52304 34451 52350
rect 34508 52304 34554 52350
rect 34612 52304 34658 52350
rect 39740 52304 39786 52350
rect 39862 52304 39908 52350
rect 39985 52304 40031 52350
rect 40108 52304 40154 52350
rect 50467 52528 50513 52574
rect 50571 52528 50617 52574
rect 50674 52528 50720 52574
rect 50777 52528 50823 52574
rect 50880 52528 50926 52574
rect 50983 52528 51029 52574
rect 51086 52528 51132 52574
rect 51189 52528 51235 52574
rect 51292 52528 51338 52574
rect 51395 52528 51441 52574
rect 43739 52304 43785 52350
rect 43906 52304 43952 52350
rect 44071 52304 44117 52350
rect 44236 52304 44282 52350
rect 33684 52080 33730 52126
rect 33787 52080 33833 52126
rect 33890 52080 33936 52126
rect 33993 52080 34039 52126
rect 34096 52080 34142 52126
rect 34199 52080 34245 52126
rect 34302 52080 34348 52126
rect 34405 52080 34451 52126
rect 34508 52080 34554 52126
rect 34612 52080 34658 52126
rect 39740 52080 39786 52126
rect 39862 52080 39908 52126
rect 39985 52080 40031 52126
rect 40108 52080 40154 52126
rect 50467 52304 50513 52350
rect 50571 52304 50617 52350
rect 50674 52304 50720 52350
rect 50777 52304 50823 52350
rect 50880 52304 50926 52350
rect 50983 52304 51029 52350
rect 51086 52304 51132 52350
rect 51189 52304 51235 52350
rect 51292 52304 51338 52350
rect 51395 52304 51441 52350
rect 50467 52080 50513 52126
rect 50571 52080 50617 52126
rect 50674 52080 50720 52126
rect 50777 52080 50823 52126
rect 50880 52080 50926 52126
rect 50983 52080 51029 52126
rect 51086 52080 51132 52126
rect 51189 52080 51235 52126
rect 51292 52080 51338 52126
rect 51395 52080 51441 52126
rect 37909 51993 37955 52039
rect 38026 51993 38072 52039
rect 38143 51993 38189 52039
rect 38261 51993 38307 52039
rect 38379 51993 38425 52039
rect 38497 51993 38543 52039
rect 33684 51856 33730 51902
rect 33787 51856 33833 51902
rect 33890 51856 33936 51902
rect 33993 51856 34039 51902
rect 34096 51856 34142 51902
rect 34199 51856 34245 51902
rect 34302 51856 34348 51902
rect 34405 51856 34451 51902
rect 34508 51856 34554 51902
rect 34612 51856 34658 51902
rect 33816 51597 33862 51643
rect 34002 51597 34048 51643
rect 34189 51597 34235 51643
rect 34376 51597 34422 51643
rect 34562 51597 34608 51643
rect 37909 51769 37955 51815
rect 38026 51769 38072 51815
rect 38143 51769 38189 51815
rect 38261 51769 38307 51815
rect 38379 51769 38425 51815
rect 38497 51769 38543 51815
rect 39641 51769 39687 51815
rect 50467 51856 50513 51902
rect 50571 51856 50617 51902
rect 50674 51856 50720 51902
rect 50777 51856 50823 51902
rect 50880 51856 50926 51902
rect 50983 51856 51029 51902
rect 51086 51856 51132 51902
rect 51189 51856 51235 51902
rect 51292 51856 51338 51902
rect 51395 51856 51441 51902
rect 37909 51545 37955 51591
rect 38026 51545 38072 51591
rect 38143 51545 38189 51591
rect 38261 51545 38307 51591
rect 38379 51545 38425 51591
rect 38497 51545 38543 51591
rect 39641 51545 39687 51591
rect 43739 51611 43785 51657
rect 43906 51611 43952 51657
rect 44071 51611 44117 51657
rect 44236 51611 44282 51657
rect 50516 51597 50562 51643
rect 50703 51597 50749 51643
rect 50890 51597 50936 51643
rect 51076 51597 51122 51643
rect 51263 51597 51309 51643
rect 33816 51211 33862 51257
rect 34002 51211 34048 51257
rect 34189 51211 34235 51257
rect 34376 51211 34422 51257
rect 34562 51211 34608 51257
rect 37909 51263 37955 51309
rect 38026 51263 38072 51309
rect 38143 51263 38189 51309
rect 38261 51263 38307 51309
rect 38379 51263 38425 51309
rect 38497 51263 38543 51309
rect 39641 51263 39687 51309
rect 33684 50952 33730 50998
rect 33787 50952 33833 50998
rect 33890 50952 33936 50998
rect 33993 50952 34039 50998
rect 34096 50952 34142 50998
rect 34199 50952 34245 50998
rect 34302 50952 34348 50998
rect 34405 50952 34451 50998
rect 34508 50952 34554 50998
rect 34612 50952 34658 50998
rect 37909 51039 37955 51085
rect 38026 51039 38072 51085
rect 38143 51039 38189 51085
rect 38261 51039 38307 51085
rect 38379 51039 38425 51085
rect 38497 51039 38543 51085
rect 43739 51197 43785 51243
rect 43906 51197 43952 51243
rect 44071 51197 44117 51243
rect 44236 51197 44282 51243
rect 39641 51039 39687 51085
rect 50516 51211 50562 51257
rect 50703 51211 50749 51257
rect 50890 51211 50936 51257
rect 51076 51211 51122 51257
rect 51263 51211 51309 51257
rect 37909 50815 37955 50861
rect 38026 50815 38072 50861
rect 38143 50815 38189 50861
rect 38261 50815 38307 50861
rect 38379 50815 38425 50861
rect 38497 50815 38543 50861
rect 50467 50952 50513 50998
rect 50571 50952 50617 50998
rect 50674 50952 50720 50998
rect 50777 50952 50823 50998
rect 50880 50952 50926 50998
rect 50983 50952 51029 50998
rect 51086 50952 51132 50998
rect 51189 50952 51235 50998
rect 51292 50952 51338 50998
rect 51395 50952 51441 50998
rect 33684 50728 33730 50774
rect 33787 50728 33833 50774
rect 33890 50728 33936 50774
rect 33993 50728 34039 50774
rect 34096 50728 34142 50774
rect 34199 50728 34245 50774
rect 34302 50728 34348 50774
rect 34405 50728 34451 50774
rect 34508 50728 34554 50774
rect 34612 50728 34658 50774
rect 39740 50728 39786 50774
rect 39862 50728 39908 50774
rect 39985 50728 40031 50774
rect 40108 50728 40154 50774
rect 33684 50504 33730 50550
rect 33787 50504 33833 50550
rect 33890 50504 33936 50550
rect 33993 50504 34039 50550
rect 34096 50504 34142 50550
rect 34199 50504 34245 50550
rect 34302 50504 34348 50550
rect 34405 50504 34451 50550
rect 34508 50504 34554 50550
rect 34612 50504 34658 50550
rect 39740 50504 39786 50550
rect 39862 50504 39908 50550
rect 39985 50504 40031 50550
rect 40108 50504 40154 50550
rect 50467 50728 50513 50774
rect 50571 50728 50617 50774
rect 50674 50728 50720 50774
rect 50777 50728 50823 50774
rect 50880 50728 50926 50774
rect 50983 50728 51029 50774
rect 51086 50728 51132 50774
rect 51189 50728 51235 50774
rect 51292 50728 51338 50774
rect 51395 50728 51441 50774
rect 43739 50504 43785 50550
rect 43906 50504 43952 50550
rect 44071 50504 44117 50550
rect 44236 50504 44282 50550
rect 33684 50280 33730 50326
rect 33787 50280 33833 50326
rect 33890 50280 33936 50326
rect 33993 50280 34039 50326
rect 34096 50280 34142 50326
rect 34199 50280 34245 50326
rect 34302 50280 34348 50326
rect 34405 50280 34451 50326
rect 34508 50280 34554 50326
rect 34612 50280 34658 50326
rect 39740 50280 39786 50326
rect 39862 50280 39908 50326
rect 39985 50280 40031 50326
rect 40108 50280 40154 50326
rect 50467 50504 50513 50550
rect 50571 50504 50617 50550
rect 50674 50504 50720 50550
rect 50777 50504 50823 50550
rect 50880 50504 50926 50550
rect 50983 50504 51029 50550
rect 51086 50504 51132 50550
rect 51189 50504 51235 50550
rect 51292 50504 51338 50550
rect 51395 50504 51441 50550
rect 50467 50280 50513 50326
rect 50571 50280 50617 50326
rect 50674 50280 50720 50326
rect 50777 50280 50823 50326
rect 50880 50280 50926 50326
rect 50983 50280 51029 50326
rect 51086 50280 51132 50326
rect 51189 50280 51235 50326
rect 51292 50280 51338 50326
rect 51395 50280 51441 50326
rect 37909 50193 37955 50239
rect 38026 50193 38072 50239
rect 38143 50193 38189 50239
rect 38261 50193 38307 50239
rect 38379 50193 38425 50239
rect 38497 50193 38543 50239
rect 33684 50056 33730 50102
rect 33787 50056 33833 50102
rect 33890 50056 33936 50102
rect 33993 50056 34039 50102
rect 34096 50056 34142 50102
rect 34199 50056 34245 50102
rect 34302 50056 34348 50102
rect 34405 50056 34451 50102
rect 34508 50056 34554 50102
rect 34612 50056 34658 50102
rect 33816 49797 33862 49843
rect 34002 49797 34048 49843
rect 34189 49797 34235 49843
rect 34376 49797 34422 49843
rect 34562 49797 34608 49843
rect 37909 49969 37955 50015
rect 38026 49969 38072 50015
rect 38143 49969 38189 50015
rect 38261 49969 38307 50015
rect 38379 49969 38425 50015
rect 38497 49969 38543 50015
rect 39641 49969 39687 50015
rect 50467 50056 50513 50102
rect 50571 50056 50617 50102
rect 50674 50056 50720 50102
rect 50777 50056 50823 50102
rect 50880 50056 50926 50102
rect 50983 50056 51029 50102
rect 51086 50056 51132 50102
rect 51189 50056 51235 50102
rect 51292 50056 51338 50102
rect 51395 50056 51441 50102
rect 37909 49745 37955 49791
rect 38026 49745 38072 49791
rect 38143 49745 38189 49791
rect 38261 49745 38307 49791
rect 38379 49745 38425 49791
rect 38497 49745 38543 49791
rect 39641 49745 39687 49791
rect 43739 49811 43785 49857
rect 43906 49811 43952 49857
rect 44071 49811 44117 49857
rect 44236 49811 44282 49857
rect 50516 49797 50562 49843
rect 50703 49797 50749 49843
rect 50890 49797 50936 49843
rect 51076 49797 51122 49843
rect 51263 49797 51309 49843
rect 33816 49411 33862 49457
rect 34002 49411 34048 49457
rect 34189 49411 34235 49457
rect 34376 49411 34422 49457
rect 34562 49411 34608 49457
rect 37909 49463 37955 49509
rect 38026 49463 38072 49509
rect 38143 49463 38189 49509
rect 38261 49463 38307 49509
rect 38379 49463 38425 49509
rect 38497 49463 38543 49509
rect 39641 49463 39687 49509
rect 33684 49152 33730 49198
rect 33787 49152 33833 49198
rect 33890 49152 33936 49198
rect 33993 49152 34039 49198
rect 34096 49152 34142 49198
rect 34199 49152 34245 49198
rect 34302 49152 34348 49198
rect 34405 49152 34451 49198
rect 34508 49152 34554 49198
rect 34612 49152 34658 49198
rect 37909 49239 37955 49285
rect 38026 49239 38072 49285
rect 38143 49239 38189 49285
rect 38261 49239 38307 49285
rect 38379 49239 38425 49285
rect 38497 49239 38543 49285
rect 43739 49397 43785 49443
rect 43906 49397 43952 49443
rect 44071 49397 44117 49443
rect 44236 49397 44282 49443
rect 39641 49239 39687 49285
rect 50516 49411 50562 49457
rect 50703 49411 50749 49457
rect 50890 49411 50936 49457
rect 51076 49411 51122 49457
rect 51263 49411 51309 49457
rect 37909 49015 37955 49061
rect 38026 49015 38072 49061
rect 38143 49015 38189 49061
rect 38261 49015 38307 49061
rect 38379 49015 38425 49061
rect 38497 49015 38543 49061
rect 50467 49152 50513 49198
rect 50571 49152 50617 49198
rect 50674 49152 50720 49198
rect 50777 49152 50823 49198
rect 50880 49152 50926 49198
rect 50983 49152 51029 49198
rect 51086 49152 51132 49198
rect 51189 49152 51235 49198
rect 51292 49152 51338 49198
rect 51395 49152 51441 49198
rect 33684 48928 33730 48974
rect 33787 48928 33833 48974
rect 33890 48928 33936 48974
rect 33993 48928 34039 48974
rect 34096 48928 34142 48974
rect 34199 48928 34245 48974
rect 34302 48928 34348 48974
rect 34405 48928 34451 48974
rect 34508 48928 34554 48974
rect 34612 48928 34658 48974
rect 39740 48928 39786 48974
rect 39862 48928 39908 48974
rect 39985 48928 40031 48974
rect 40108 48928 40154 48974
rect 33684 48704 33730 48750
rect 33787 48704 33833 48750
rect 33890 48704 33936 48750
rect 33993 48704 34039 48750
rect 34096 48704 34142 48750
rect 34199 48704 34245 48750
rect 34302 48704 34348 48750
rect 34405 48704 34451 48750
rect 34508 48704 34554 48750
rect 34612 48704 34658 48750
rect 39740 48704 39786 48750
rect 39862 48704 39908 48750
rect 39985 48704 40031 48750
rect 40108 48704 40154 48750
rect 50467 48928 50513 48974
rect 50571 48928 50617 48974
rect 50674 48928 50720 48974
rect 50777 48928 50823 48974
rect 50880 48928 50926 48974
rect 50983 48928 51029 48974
rect 51086 48928 51132 48974
rect 51189 48928 51235 48974
rect 51292 48928 51338 48974
rect 51395 48928 51441 48974
rect 43739 48704 43785 48750
rect 43906 48704 43952 48750
rect 44071 48704 44117 48750
rect 44236 48704 44282 48750
rect 33684 48480 33730 48526
rect 33787 48480 33833 48526
rect 33890 48480 33936 48526
rect 33993 48480 34039 48526
rect 34096 48480 34142 48526
rect 34199 48480 34245 48526
rect 34302 48480 34348 48526
rect 34405 48480 34451 48526
rect 34508 48480 34554 48526
rect 34612 48480 34658 48526
rect 39740 48480 39786 48526
rect 39862 48480 39908 48526
rect 39985 48480 40031 48526
rect 40108 48480 40154 48526
rect 50467 48704 50513 48750
rect 50571 48704 50617 48750
rect 50674 48704 50720 48750
rect 50777 48704 50823 48750
rect 50880 48704 50926 48750
rect 50983 48704 51029 48750
rect 51086 48704 51132 48750
rect 51189 48704 51235 48750
rect 51292 48704 51338 48750
rect 51395 48704 51441 48750
rect 50467 48480 50513 48526
rect 50571 48480 50617 48526
rect 50674 48480 50720 48526
rect 50777 48480 50823 48526
rect 50880 48480 50926 48526
rect 50983 48480 51029 48526
rect 51086 48480 51132 48526
rect 51189 48480 51235 48526
rect 51292 48480 51338 48526
rect 51395 48480 51441 48526
rect 37909 48393 37955 48439
rect 38026 48393 38072 48439
rect 38143 48393 38189 48439
rect 38261 48393 38307 48439
rect 38379 48393 38425 48439
rect 38497 48393 38543 48439
rect 33684 48256 33730 48302
rect 33787 48256 33833 48302
rect 33890 48256 33936 48302
rect 33993 48256 34039 48302
rect 34096 48256 34142 48302
rect 34199 48256 34245 48302
rect 34302 48256 34348 48302
rect 34405 48256 34451 48302
rect 34508 48256 34554 48302
rect 34612 48256 34658 48302
rect 33816 47997 33862 48043
rect 34002 47997 34048 48043
rect 34189 47997 34235 48043
rect 34376 47997 34422 48043
rect 34562 47997 34608 48043
rect 37909 48169 37955 48215
rect 38026 48169 38072 48215
rect 38143 48169 38189 48215
rect 38261 48169 38307 48215
rect 38379 48169 38425 48215
rect 38497 48169 38543 48215
rect 39641 48169 39687 48215
rect 50467 48256 50513 48302
rect 50571 48256 50617 48302
rect 50674 48256 50720 48302
rect 50777 48256 50823 48302
rect 50880 48256 50926 48302
rect 50983 48256 51029 48302
rect 51086 48256 51132 48302
rect 51189 48256 51235 48302
rect 51292 48256 51338 48302
rect 51395 48256 51441 48302
rect 37909 47945 37955 47991
rect 38026 47945 38072 47991
rect 38143 47945 38189 47991
rect 38261 47945 38307 47991
rect 38379 47945 38425 47991
rect 38497 47945 38543 47991
rect 39641 47945 39687 47991
rect 43739 48011 43785 48057
rect 43906 48011 43952 48057
rect 44071 48011 44117 48057
rect 44236 48011 44282 48057
rect 50516 47997 50562 48043
rect 50703 47997 50749 48043
rect 50890 47997 50936 48043
rect 51076 47997 51122 48043
rect 51263 47997 51309 48043
rect 33816 47611 33862 47657
rect 34002 47611 34048 47657
rect 34189 47611 34235 47657
rect 34376 47611 34422 47657
rect 34562 47611 34608 47657
rect 37909 47663 37955 47709
rect 38026 47663 38072 47709
rect 38143 47663 38189 47709
rect 38261 47663 38307 47709
rect 38379 47663 38425 47709
rect 38497 47663 38543 47709
rect 39641 47663 39687 47709
rect 33684 47352 33730 47398
rect 33787 47352 33833 47398
rect 33890 47352 33936 47398
rect 33993 47352 34039 47398
rect 34096 47352 34142 47398
rect 34199 47352 34245 47398
rect 34302 47352 34348 47398
rect 34405 47352 34451 47398
rect 34508 47352 34554 47398
rect 34612 47352 34658 47398
rect 37909 47439 37955 47485
rect 38026 47439 38072 47485
rect 38143 47439 38189 47485
rect 38261 47439 38307 47485
rect 38379 47439 38425 47485
rect 38497 47439 38543 47485
rect 43739 47597 43785 47643
rect 43906 47597 43952 47643
rect 44071 47597 44117 47643
rect 44236 47597 44282 47643
rect 39641 47439 39687 47485
rect 50516 47611 50562 47657
rect 50703 47611 50749 47657
rect 50890 47611 50936 47657
rect 51076 47611 51122 47657
rect 51263 47611 51309 47657
rect 37909 47215 37955 47261
rect 38026 47215 38072 47261
rect 38143 47215 38189 47261
rect 38261 47215 38307 47261
rect 38379 47215 38425 47261
rect 38497 47215 38543 47261
rect 50467 47352 50513 47398
rect 50571 47352 50617 47398
rect 50674 47352 50720 47398
rect 50777 47352 50823 47398
rect 50880 47352 50926 47398
rect 50983 47352 51029 47398
rect 51086 47352 51132 47398
rect 51189 47352 51235 47398
rect 51292 47352 51338 47398
rect 51395 47352 51441 47398
rect 33684 47128 33730 47174
rect 33787 47128 33833 47174
rect 33890 47128 33936 47174
rect 33993 47128 34039 47174
rect 34096 47128 34142 47174
rect 34199 47128 34245 47174
rect 34302 47128 34348 47174
rect 34405 47128 34451 47174
rect 34508 47128 34554 47174
rect 34612 47128 34658 47174
rect 39740 47128 39786 47174
rect 39862 47128 39908 47174
rect 39985 47128 40031 47174
rect 40108 47128 40154 47174
rect 33684 46904 33730 46950
rect 33787 46904 33833 46950
rect 33890 46904 33936 46950
rect 33993 46904 34039 46950
rect 34096 46904 34142 46950
rect 34199 46904 34245 46950
rect 34302 46904 34348 46950
rect 34405 46904 34451 46950
rect 34508 46904 34554 46950
rect 34612 46904 34658 46950
rect 39740 46904 39786 46950
rect 39862 46904 39908 46950
rect 39985 46904 40031 46950
rect 40108 46904 40154 46950
rect 50467 47128 50513 47174
rect 50571 47128 50617 47174
rect 50674 47128 50720 47174
rect 50777 47128 50823 47174
rect 50880 47128 50926 47174
rect 50983 47128 51029 47174
rect 51086 47128 51132 47174
rect 51189 47128 51235 47174
rect 51292 47128 51338 47174
rect 51395 47128 51441 47174
rect 43739 46904 43785 46950
rect 43906 46904 43952 46950
rect 44071 46904 44117 46950
rect 44236 46904 44282 46950
rect 33684 46680 33730 46726
rect 33787 46680 33833 46726
rect 33890 46680 33936 46726
rect 33993 46680 34039 46726
rect 34096 46680 34142 46726
rect 34199 46680 34245 46726
rect 34302 46680 34348 46726
rect 34405 46680 34451 46726
rect 34508 46680 34554 46726
rect 34612 46680 34658 46726
rect 39740 46680 39786 46726
rect 39862 46680 39908 46726
rect 39985 46680 40031 46726
rect 40108 46680 40154 46726
rect 50467 46904 50513 46950
rect 50571 46904 50617 46950
rect 50674 46904 50720 46950
rect 50777 46904 50823 46950
rect 50880 46904 50926 46950
rect 50983 46904 51029 46950
rect 51086 46904 51132 46950
rect 51189 46904 51235 46950
rect 51292 46904 51338 46950
rect 51395 46904 51441 46950
rect 50467 46680 50513 46726
rect 50571 46680 50617 46726
rect 50674 46680 50720 46726
rect 50777 46680 50823 46726
rect 50880 46680 50926 46726
rect 50983 46680 51029 46726
rect 51086 46680 51132 46726
rect 51189 46680 51235 46726
rect 51292 46680 51338 46726
rect 51395 46680 51441 46726
rect 37909 46593 37955 46639
rect 38026 46593 38072 46639
rect 38143 46593 38189 46639
rect 38261 46593 38307 46639
rect 38379 46593 38425 46639
rect 38497 46593 38543 46639
rect 33684 46456 33730 46502
rect 33787 46456 33833 46502
rect 33890 46456 33936 46502
rect 33993 46456 34039 46502
rect 34096 46456 34142 46502
rect 34199 46456 34245 46502
rect 34302 46456 34348 46502
rect 34405 46456 34451 46502
rect 34508 46456 34554 46502
rect 34612 46456 34658 46502
rect 33816 46197 33862 46243
rect 34002 46197 34048 46243
rect 34189 46197 34235 46243
rect 34376 46197 34422 46243
rect 34562 46197 34608 46243
rect 37909 46369 37955 46415
rect 38026 46369 38072 46415
rect 38143 46369 38189 46415
rect 38261 46369 38307 46415
rect 38379 46369 38425 46415
rect 38497 46369 38543 46415
rect 39641 46369 39687 46415
rect 50467 46456 50513 46502
rect 50571 46456 50617 46502
rect 50674 46456 50720 46502
rect 50777 46456 50823 46502
rect 50880 46456 50926 46502
rect 50983 46456 51029 46502
rect 51086 46456 51132 46502
rect 51189 46456 51235 46502
rect 51292 46456 51338 46502
rect 51395 46456 51441 46502
rect 37909 46145 37955 46191
rect 38026 46145 38072 46191
rect 38143 46145 38189 46191
rect 38261 46145 38307 46191
rect 38379 46145 38425 46191
rect 38497 46145 38543 46191
rect 39641 46145 39687 46191
rect 43739 46211 43785 46257
rect 43906 46211 43952 46257
rect 44071 46211 44117 46257
rect 44236 46211 44282 46257
rect 50516 46197 50562 46243
rect 50703 46197 50749 46243
rect 50890 46197 50936 46243
rect 51076 46197 51122 46243
rect 51263 46197 51309 46243
rect 33816 45811 33862 45857
rect 34002 45811 34048 45857
rect 34189 45811 34235 45857
rect 34376 45811 34422 45857
rect 34562 45811 34608 45857
rect 37909 45863 37955 45909
rect 38026 45863 38072 45909
rect 38143 45863 38189 45909
rect 38261 45863 38307 45909
rect 38379 45863 38425 45909
rect 38497 45863 38543 45909
rect 39641 45863 39687 45909
rect 33684 45552 33730 45598
rect 33787 45552 33833 45598
rect 33890 45552 33936 45598
rect 33993 45552 34039 45598
rect 34096 45552 34142 45598
rect 34199 45552 34245 45598
rect 34302 45552 34348 45598
rect 34405 45552 34451 45598
rect 34508 45552 34554 45598
rect 34612 45552 34658 45598
rect 37909 45639 37955 45685
rect 38026 45639 38072 45685
rect 38143 45639 38189 45685
rect 38261 45639 38307 45685
rect 38379 45639 38425 45685
rect 38497 45639 38543 45685
rect 43739 45797 43785 45843
rect 43906 45797 43952 45843
rect 44071 45797 44117 45843
rect 44236 45797 44282 45843
rect 39641 45639 39687 45685
rect 50516 45811 50562 45857
rect 50703 45811 50749 45857
rect 50890 45811 50936 45857
rect 51076 45811 51122 45857
rect 51263 45811 51309 45857
rect 37909 45415 37955 45461
rect 38026 45415 38072 45461
rect 38143 45415 38189 45461
rect 38261 45415 38307 45461
rect 38379 45415 38425 45461
rect 38497 45415 38543 45461
rect 50467 45552 50513 45598
rect 50571 45552 50617 45598
rect 50674 45552 50720 45598
rect 50777 45552 50823 45598
rect 50880 45552 50926 45598
rect 50983 45552 51029 45598
rect 51086 45552 51132 45598
rect 51189 45552 51235 45598
rect 51292 45552 51338 45598
rect 51395 45552 51441 45598
rect 33684 45328 33730 45374
rect 33787 45328 33833 45374
rect 33890 45328 33936 45374
rect 33993 45328 34039 45374
rect 34096 45328 34142 45374
rect 34199 45328 34245 45374
rect 34302 45328 34348 45374
rect 34405 45328 34451 45374
rect 34508 45328 34554 45374
rect 34612 45328 34658 45374
rect 39740 45328 39786 45374
rect 39862 45328 39908 45374
rect 39985 45328 40031 45374
rect 40108 45328 40154 45374
rect 33684 45104 33730 45150
rect 33787 45104 33833 45150
rect 33890 45104 33936 45150
rect 33993 45104 34039 45150
rect 34096 45104 34142 45150
rect 34199 45104 34245 45150
rect 34302 45104 34348 45150
rect 34405 45104 34451 45150
rect 34508 45104 34554 45150
rect 34612 45104 34658 45150
rect 39740 45104 39786 45150
rect 39862 45104 39908 45150
rect 39985 45104 40031 45150
rect 40108 45104 40154 45150
rect 50467 45328 50513 45374
rect 50571 45328 50617 45374
rect 50674 45328 50720 45374
rect 50777 45328 50823 45374
rect 50880 45328 50926 45374
rect 50983 45328 51029 45374
rect 51086 45328 51132 45374
rect 51189 45328 51235 45374
rect 51292 45328 51338 45374
rect 51395 45328 51441 45374
rect 43739 45104 43785 45150
rect 43906 45104 43952 45150
rect 44071 45104 44117 45150
rect 44236 45104 44282 45150
rect 33684 44880 33730 44926
rect 33787 44880 33833 44926
rect 33890 44880 33936 44926
rect 33993 44880 34039 44926
rect 34096 44880 34142 44926
rect 34199 44880 34245 44926
rect 34302 44880 34348 44926
rect 34405 44880 34451 44926
rect 34508 44880 34554 44926
rect 34612 44880 34658 44926
rect 39740 44880 39786 44926
rect 39862 44880 39908 44926
rect 39985 44880 40031 44926
rect 40108 44880 40154 44926
rect 50467 45104 50513 45150
rect 50571 45104 50617 45150
rect 50674 45104 50720 45150
rect 50777 45104 50823 45150
rect 50880 45104 50926 45150
rect 50983 45104 51029 45150
rect 51086 45104 51132 45150
rect 51189 45104 51235 45150
rect 51292 45104 51338 45150
rect 51395 45104 51441 45150
rect 50467 44880 50513 44926
rect 50571 44880 50617 44926
rect 50674 44880 50720 44926
rect 50777 44880 50823 44926
rect 50880 44880 50926 44926
rect 50983 44880 51029 44926
rect 51086 44880 51132 44926
rect 51189 44880 51235 44926
rect 51292 44880 51338 44926
rect 51395 44880 51441 44926
rect 37909 44793 37955 44839
rect 38026 44793 38072 44839
rect 38143 44793 38189 44839
rect 38261 44793 38307 44839
rect 38379 44793 38425 44839
rect 38497 44793 38543 44839
rect 33684 44656 33730 44702
rect 33787 44656 33833 44702
rect 33890 44656 33936 44702
rect 33993 44656 34039 44702
rect 34096 44656 34142 44702
rect 34199 44656 34245 44702
rect 34302 44656 34348 44702
rect 34405 44656 34451 44702
rect 34508 44656 34554 44702
rect 34612 44656 34658 44702
rect 33816 44397 33862 44443
rect 34002 44397 34048 44443
rect 34189 44397 34235 44443
rect 34376 44397 34422 44443
rect 34562 44397 34608 44443
rect 37909 44569 37955 44615
rect 38026 44569 38072 44615
rect 38143 44569 38189 44615
rect 38261 44569 38307 44615
rect 38379 44569 38425 44615
rect 38497 44569 38543 44615
rect 39641 44569 39687 44615
rect 50467 44656 50513 44702
rect 50571 44656 50617 44702
rect 50674 44656 50720 44702
rect 50777 44656 50823 44702
rect 50880 44656 50926 44702
rect 50983 44656 51029 44702
rect 51086 44656 51132 44702
rect 51189 44656 51235 44702
rect 51292 44656 51338 44702
rect 51395 44656 51441 44702
rect 37909 44345 37955 44391
rect 38026 44345 38072 44391
rect 38143 44345 38189 44391
rect 38261 44345 38307 44391
rect 38379 44345 38425 44391
rect 38497 44345 38543 44391
rect 39641 44345 39687 44391
rect 43739 44411 43785 44457
rect 43906 44411 43952 44457
rect 44071 44411 44117 44457
rect 44236 44411 44282 44457
rect 50516 44397 50562 44443
rect 50703 44397 50749 44443
rect 50890 44397 50936 44443
rect 51076 44397 51122 44443
rect 51263 44397 51309 44443
rect 33816 44011 33862 44057
rect 34002 44011 34048 44057
rect 34189 44011 34235 44057
rect 34376 44011 34422 44057
rect 34562 44011 34608 44057
rect 37909 44063 37955 44109
rect 38026 44063 38072 44109
rect 38143 44063 38189 44109
rect 38261 44063 38307 44109
rect 38379 44063 38425 44109
rect 38497 44063 38543 44109
rect 39641 44063 39687 44109
rect 33684 43752 33730 43798
rect 33787 43752 33833 43798
rect 33890 43752 33936 43798
rect 33993 43752 34039 43798
rect 34096 43752 34142 43798
rect 34199 43752 34245 43798
rect 34302 43752 34348 43798
rect 34405 43752 34451 43798
rect 34508 43752 34554 43798
rect 34612 43752 34658 43798
rect 37909 43839 37955 43885
rect 38026 43839 38072 43885
rect 38143 43839 38189 43885
rect 38261 43839 38307 43885
rect 38379 43839 38425 43885
rect 38497 43839 38543 43885
rect 43739 43997 43785 44043
rect 43906 43997 43952 44043
rect 44071 43997 44117 44043
rect 44236 43997 44282 44043
rect 39641 43839 39687 43885
rect 50516 44011 50562 44057
rect 50703 44011 50749 44057
rect 50890 44011 50936 44057
rect 51076 44011 51122 44057
rect 51263 44011 51309 44057
rect 37909 43615 37955 43661
rect 38026 43615 38072 43661
rect 38143 43615 38189 43661
rect 38261 43615 38307 43661
rect 38379 43615 38425 43661
rect 38497 43615 38543 43661
rect 50467 43752 50513 43798
rect 50571 43752 50617 43798
rect 50674 43752 50720 43798
rect 50777 43752 50823 43798
rect 50880 43752 50926 43798
rect 50983 43752 51029 43798
rect 51086 43752 51132 43798
rect 51189 43752 51235 43798
rect 51292 43752 51338 43798
rect 51395 43752 51441 43798
rect 33684 43528 33730 43574
rect 33787 43528 33833 43574
rect 33890 43528 33936 43574
rect 33993 43528 34039 43574
rect 34096 43528 34142 43574
rect 34199 43528 34245 43574
rect 34302 43528 34348 43574
rect 34405 43528 34451 43574
rect 34508 43528 34554 43574
rect 34612 43528 34658 43574
rect 39740 43528 39786 43574
rect 39862 43528 39908 43574
rect 39985 43528 40031 43574
rect 40108 43528 40154 43574
rect 33684 43304 33730 43350
rect 33787 43304 33833 43350
rect 33890 43304 33936 43350
rect 33993 43304 34039 43350
rect 34096 43304 34142 43350
rect 34199 43304 34245 43350
rect 34302 43304 34348 43350
rect 34405 43304 34451 43350
rect 34508 43304 34554 43350
rect 34612 43304 34658 43350
rect 39740 43304 39786 43350
rect 39862 43304 39908 43350
rect 39985 43304 40031 43350
rect 40108 43304 40154 43350
rect 50467 43528 50513 43574
rect 50571 43528 50617 43574
rect 50674 43528 50720 43574
rect 50777 43528 50823 43574
rect 50880 43528 50926 43574
rect 50983 43528 51029 43574
rect 51086 43528 51132 43574
rect 51189 43528 51235 43574
rect 51292 43528 51338 43574
rect 51395 43528 51441 43574
rect 43739 43304 43785 43350
rect 43906 43304 43952 43350
rect 44071 43304 44117 43350
rect 44236 43304 44282 43350
rect 33684 43080 33730 43126
rect 33787 43080 33833 43126
rect 33890 43080 33936 43126
rect 33993 43080 34039 43126
rect 34096 43080 34142 43126
rect 34199 43080 34245 43126
rect 34302 43080 34348 43126
rect 34405 43080 34451 43126
rect 34508 43080 34554 43126
rect 34612 43080 34658 43126
rect 39740 43080 39786 43126
rect 39862 43080 39908 43126
rect 39985 43080 40031 43126
rect 40108 43080 40154 43126
rect 50467 43304 50513 43350
rect 50571 43304 50617 43350
rect 50674 43304 50720 43350
rect 50777 43304 50823 43350
rect 50880 43304 50926 43350
rect 50983 43304 51029 43350
rect 51086 43304 51132 43350
rect 51189 43304 51235 43350
rect 51292 43304 51338 43350
rect 51395 43304 51441 43350
rect 50467 43080 50513 43126
rect 50571 43080 50617 43126
rect 50674 43080 50720 43126
rect 50777 43080 50823 43126
rect 50880 43080 50926 43126
rect 50983 43080 51029 43126
rect 51086 43080 51132 43126
rect 51189 43080 51235 43126
rect 51292 43080 51338 43126
rect 51395 43080 51441 43126
rect 37909 42993 37955 43039
rect 38026 42993 38072 43039
rect 38143 42993 38189 43039
rect 38261 42993 38307 43039
rect 38379 42993 38425 43039
rect 38497 42993 38543 43039
rect 33684 42856 33730 42902
rect 33787 42856 33833 42902
rect 33890 42856 33936 42902
rect 33993 42856 34039 42902
rect 34096 42856 34142 42902
rect 34199 42856 34245 42902
rect 34302 42856 34348 42902
rect 34405 42856 34451 42902
rect 34508 42856 34554 42902
rect 34612 42856 34658 42902
rect 33816 42597 33862 42643
rect 34002 42597 34048 42643
rect 34189 42597 34235 42643
rect 34376 42597 34422 42643
rect 34562 42597 34608 42643
rect 37909 42769 37955 42815
rect 38026 42769 38072 42815
rect 38143 42769 38189 42815
rect 38261 42769 38307 42815
rect 38379 42769 38425 42815
rect 38497 42769 38543 42815
rect 39641 42769 39687 42815
rect 50467 42856 50513 42902
rect 50571 42856 50617 42902
rect 50674 42856 50720 42902
rect 50777 42856 50823 42902
rect 50880 42856 50926 42902
rect 50983 42856 51029 42902
rect 51086 42856 51132 42902
rect 51189 42856 51235 42902
rect 51292 42856 51338 42902
rect 51395 42856 51441 42902
rect 37909 42545 37955 42591
rect 38026 42545 38072 42591
rect 38143 42545 38189 42591
rect 38261 42545 38307 42591
rect 38379 42545 38425 42591
rect 38497 42545 38543 42591
rect 39641 42545 39687 42591
rect 43739 42611 43785 42657
rect 43906 42611 43952 42657
rect 44071 42611 44117 42657
rect 44236 42611 44282 42657
rect 50516 42597 50562 42643
rect 50703 42597 50749 42643
rect 50890 42597 50936 42643
rect 51076 42597 51122 42643
rect 51263 42597 51309 42643
rect 33816 42211 33862 42257
rect 34002 42211 34048 42257
rect 34189 42211 34235 42257
rect 34376 42211 34422 42257
rect 34562 42211 34608 42257
rect 37909 42263 37955 42309
rect 38026 42263 38072 42309
rect 38143 42263 38189 42309
rect 38261 42263 38307 42309
rect 38379 42263 38425 42309
rect 38497 42263 38543 42309
rect 39641 42263 39687 42309
rect 33684 41952 33730 41998
rect 33787 41952 33833 41998
rect 33890 41952 33936 41998
rect 33993 41952 34039 41998
rect 34096 41952 34142 41998
rect 34199 41952 34245 41998
rect 34302 41952 34348 41998
rect 34405 41952 34451 41998
rect 34508 41952 34554 41998
rect 34612 41952 34658 41998
rect 37909 42039 37955 42085
rect 38026 42039 38072 42085
rect 38143 42039 38189 42085
rect 38261 42039 38307 42085
rect 38379 42039 38425 42085
rect 38497 42039 38543 42085
rect 43739 42197 43785 42243
rect 43906 42197 43952 42243
rect 44071 42197 44117 42243
rect 44236 42197 44282 42243
rect 39641 42039 39687 42085
rect 50516 42211 50562 42257
rect 50703 42211 50749 42257
rect 50890 42211 50936 42257
rect 51076 42211 51122 42257
rect 51263 42211 51309 42257
rect 37909 41815 37955 41861
rect 38026 41815 38072 41861
rect 38143 41815 38189 41861
rect 38261 41815 38307 41861
rect 38379 41815 38425 41861
rect 38497 41815 38543 41861
rect 50467 41952 50513 41998
rect 50571 41952 50617 41998
rect 50674 41952 50720 41998
rect 50777 41952 50823 41998
rect 50880 41952 50926 41998
rect 50983 41952 51029 41998
rect 51086 41952 51132 41998
rect 51189 41952 51235 41998
rect 51292 41952 51338 41998
rect 51395 41952 51441 41998
rect 33684 41728 33730 41774
rect 33787 41728 33833 41774
rect 33890 41728 33936 41774
rect 33993 41728 34039 41774
rect 34096 41728 34142 41774
rect 34199 41728 34245 41774
rect 34302 41728 34348 41774
rect 34405 41728 34451 41774
rect 34508 41728 34554 41774
rect 34612 41728 34658 41774
rect 39740 41728 39786 41774
rect 39862 41728 39908 41774
rect 39985 41728 40031 41774
rect 40108 41728 40154 41774
rect 33684 41504 33730 41550
rect 33787 41504 33833 41550
rect 33890 41504 33936 41550
rect 33993 41504 34039 41550
rect 34096 41504 34142 41550
rect 34199 41504 34245 41550
rect 34302 41504 34348 41550
rect 34405 41504 34451 41550
rect 34508 41504 34554 41550
rect 34612 41504 34658 41550
rect 39740 41504 39786 41550
rect 39862 41504 39908 41550
rect 39985 41504 40031 41550
rect 40108 41504 40154 41550
rect 50467 41728 50513 41774
rect 50571 41728 50617 41774
rect 50674 41728 50720 41774
rect 50777 41728 50823 41774
rect 50880 41728 50926 41774
rect 50983 41728 51029 41774
rect 51086 41728 51132 41774
rect 51189 41728 51235 41774
rect 51292 41728 51338 41774
rect 51395 41728 51441 41774
rect 43739 41504 43785 41550
rect 43906 41504 43952 41550
rect 44071 41504 44117 41550
rect 44236 41504 44282 41550
rect 33684 41280 33730 41326
rect 33787 41280 33833 41326
rect 33890 41280 33936 41326
rect 33993 41280 34039 41326
rect 34096 41280 34142 41326
rect 34199 41280 34245 41326
rect 34302 41280 34348 41326
rect 34405 41280 34451 41326
rect 34508 41280 34554 41326
rect 34612 41280 34658 41326
rect 39740 41280 39786 41326
rect 39862 41280 39908 41326
rect 39985 41280 40031 41326
rect 40108 41280 40154 41326
rect 50467 41504 50513 41550
rect 50571 41504 50617 41550
rect 50674 41504 50720 41550
rect 50777 41504 50823 41550
rect 50880 41504 50926 41550
rect 50983 41504 51029 41550
rect 51086 41504 51132 41550
rect 51189 41504 51235 41550
rect 51292 41504 51338 41550
rect 51395 41504 51441 41550
rect 50467 41280 50513 41326
rect 50571 41280 50617 41326
rect 50674 41280 50720 41326
rect 50777 41280 50823 41326
rect 50880 41280 50926 41326
rect 50983 41280 51029 41326
rect 51086 41280 51132 41326
rect 51189 41280 51235 41326
rect 51292 41280 51338 41326
rect 51395 41280 51441 41326
rect 37909 41193 37955 41239
rect 38026 41193 38072 41239
rect 38143 41193 38189 41239
rect 38261 41193 38307 41239
rect 38379 41193 38425 41239
rect 38497 41193 38543 41239
rect 33684 41056 33730 41102
rect 33787 41056 33833 41102
rect 33890 41056 33936 41102
rect 33993 41056 34039 41102
rect 34096 41056 34142 41102
rect 34199 41056 34245 41102
rect 34302 41056 34348 41102
rect 34405 41056 34451 41102
rect 34508 41056 34554 41102
rect 34612 41056 34658 41102
rect 33816 40797 33862 40843
rect 34002 40797 34048 40843
rect 34189 40797 34235 40843
rect 34376 40797 34422 40843
rect 34562 40797 34608 40843
rect 37909 40969 37955 41015
rect 38026 40969 38072 41015
rect 38143 40969 38189 41015
rect 38261 40969 38307 41015
rect 38379 40969 38425 41015
rect 38497 40969 38543 41015
rect 39641 40969 39687 41015
rect 50467 41056 50513 41102
rect 50571 41056 50617 41102
rect 50674 41056 50720 41102
rect 50777 41056 50823 41102
rect 50880 41056 50926 41102
rect 50983 41056 51029 41102
rect 51086 41056 51132 41102
rect 51189 41056 51235 41102
rect 51292 41056 51338 41102
rect 51395 41056 51441 41102
rect 37909 40745 37955 40791
rect 38026 40745 38072 40791
rect 38143 40745 38189 40791
rect 38261 40745 38307 40791
rect 38379 40745 38425 40791
rect 38497 40745 38543 40791
rect 39641 40745 39687 40791
rect 43739 40811 43785 40857
rect 43906 40811 43952 40857
rect 44071 40811 44117 40857
rect 44236 40811 44282 40857
rect 50516 40797 50562 40843
rect 50703 40797 50749 40843
rect 50890 40797 50936 40843
rect 51076 40797 51122 40843
rect 51263 40797 51309 40843
rect 33816 40411 33862 40457
rect 34002 40411 34048 40457
rect 34189 40411 34235 40457
rect 34376 40411 34422 40457
rect 34562 40411 34608 40457
rect 37909 40463 37955 40509
rect 38026 40463 38072 40509
rect 38143 40463 38189 40509
rect 38261 40463 38307 40509
rect 38379 40463 38425 40509
rect 38497 40463 38543 40509
rect 39641 40463 39687 40509
rect 33684 40152 33730 40198
rect 33787 40152 33833 40198
rect 33890 40152 33936 40198
rect 33993 40152 34039 40198
rect 34096 40152 34142 40198
rect 34199 40152 34245 40198
rect 34302 40152 34348 40198
rect 34405 40152 34451 40198
rect 34508 40152 34554 40198
rect 34612 40152 34658 40198
rect 37909 40239 37955 40285
rect 38026 40239 38072 40285
rect 38143 40239 38189 40285
rect 38261 40239 38307 40285
rect 38379 40239 38425 40285
rect 38497 40239 38543 40285
rect 43739 40397 43785 40443
rect 43906 40397 43952 40443
rect 44071 40397 44117 40443
rect 44236 40397 44282 40443
rect 39641 40239 39687 40285
rect 50516 40411 50562 40457
rect 50703 40411 50749 40457
rect 50890 40411 50936 40457
rect 51076 40411 51122 40457
rect 51263 40411 51309 40457
rect 37909 40015 37955 40061
rect 38026 40015 38072 40061
rect 38143 40015 38189 40061
rect 38261 40015 38307 40061
rect 38379 40015 38425 40061
rect 38497 40015 38543 40061
rect 50467 40152 50513 40198
rect 50571 40152 50617 40198
rect 50674 40152 50720 40198
rect 50777 40152 50823 40198
rect 50880 40152 50926 40198
rect 50983 40152 51029 40198
rect 51086 40152 51132 40198
rect 51189 40152 51235 40198
rect 51292 40152 51338 40198
rect 51395 40152 51441 40198
rect 33684 39928 33730 39974
rect 33787 39928 33833 39974
rect 33890 39928 33936 39974
rect 33993 39928 34039 39974
rect 34096 39928 34142 39974
rect 34199 39928 34245 39974
rect 34302 39928 34348 39974
rect 34405 39928 34451 39974
rect 34508 39928 34554 39974
rect 34612 39928 34658 39974
rect 39740 39928 39786 39974
rect 39862 39928 39908 39974
rect 39985 39928 40031 39974
rect 40108 39928 40154 39974
rect 33684 39704 33730 39750
rect 33787 39704 33833 39750
rect 33890 39704 33936 39750
rect 33993 39704 34039 39750
rect 34096 39704 34142 39750
rect 34199 39704 34245 39750
rect 34302 39704 34348 39750
rect 34405 39704 34451 39750
rect 34508 39704 34554 39750
rect 34612 39704 34658 39750
rect 39740 39704 39786 39750
rect 39862 39704 39908 39750
rect 39985 39704 40031 39750
rect 40108 39704 40154 39750
rect 50467 39928 50513 39974
rect 50571 39928 50617 39974
rect 50674 39928 50720 39974
rect 50777 39928 50823 39974
rect 50880 39928 50926 39974
rect 50983 39928 51029 39974
rect 51086 39928 51132 39974
rect 51189 39928 51235 39974
rect 51292 39928 51338 39974
rect 51395 39928 51441 39974
rect 43739 39704 43785 39750
rect 43906 39704 43952 39750
rect 44071 39704 44117 39750
rect 44236 39704 44282 39750
rect 33684 39480 33730 39526
rect 33787 39480 33833 39526
rect 33890 39480 33936 39526
rect 33993 39480 34039 39526
rect 34096 39480 34142 39526
rect 34199 39480 34245 39526
rect 34302 39480 34348 39526
rect 34405 39480 34451 39526
rect 34508 39480 34554 39526
rect 34612 39480 34658 39526
rect 39740 39480 39786 39526
rect 39862 39480 39908 39526
rect 39985 39480 40031 39526
rect 40108 39480 40154 39526
rect 50467 39704 50513 39750
rect 50571 39704 50617 39750
rect 50674 39704 50720 39750
rect 50777 39704 50823 39750
rect 50880 39704 50926 39750
rect 50983 39704 51029 39750
rect 51086 39704 51132 39750
rect 51189 39704 51235 39750
rect 51292 39704 51338 39750
rect 51395 39704 51441 39750
rect 50467 39480 50513 39526
rect 50571 39480 50617 39526
rect 50674 39480 50720 39526
rect 50777 39480 50823 39526
rect 50880 39480 50926 39526
rect 50983 39480 51029 39526
rect 51086 39480 51132 39526
rect 51189 39480 51235 39526
rect 51292 39480 51338 39526
rect 51395 39480 51441 39526
rect 37909 39393 37955 39439
rect 38026 39393 38072 39439
rect 38143 39393 38189 39439
rect 38261 39393 38307 39439
rect 38379 39393 38425 39439
rect 38497 39393 38543 39439
rect 33684 39256 33730 39302
rect 33787 39256 33833 39302
rect 33890 39256 33936 39302
rect 33993 39256 34039 39302
rect 34096 39256 34142 39302
rect 34199 39256 34245 39302
rect 34302 39256 34348 39302
rect 34405 39256 34451 39302
rect 34508 39256 34554 39302
rect 34612 39256 34658 39302
rect 33816 38997 33862 39043
rect 34002 38997 34048 39043
rect 34189 38997 34235 39043
rect 34376 38997 34422 39043
rect 34562 38997 34608 39043
rect 37909 39169 37955 39215
rect 38026 39169 38072 39215
rect 38143 39169 38189 39215
rect 38261 39169 38307 39215
rect 38379 39169 38425 39215
rect 38497 39169 38543 39215
rect 39641 39169 39687 39215
rect 50467 39256 50513 39302
rect 50571 39256 50617 39302
rect 50674 39256 50720 39302
rect 50777 39256 50823 39302
rect 50880 39256 50926 39302
rect 50983 39256 51029 39302
rect 51086 39256 51132 39302
rect 51189 39256 51235 39302
rect 51292 39256 51338 39302
rect 51395 39256 51441 39302
rect 37909 38945 37955 38991
rect 38026 38945 38072 38991
rect 38143 38945 38189 38991
rect 38261 38945 38307 38991
rect 38379 38945 38425 38991
rect 38497 38945 38543 38991
rect 39641 38945 39687 38991
rect 43739 39011 43785 39057
rect 43906 39011 43952 39057
rect 44071 39011 44117 39057
rect 44236 39011 44282 39057
rect 50516 38997 50562 39043
rect 50703 38997 50749 39043
rect 50890 38997 50936 39043
rect 51076 38997 51122 39043
rect 51263 38997 51309 39043
rect 33816 38611 33862 38657
rect 34002 38611 34048 38657
rect 34189 38611 34235 38657
rect 34376 38611 34422 38657
rect 34562 38611 34608 38657
rect 37909 38663 37955 38709
rect 38026 38663 38072 38709
rect 38143 38663 38189 38709
rect 38261 38663 38307 38709
rect 38379 38663 38425 38709
rect 38497 38663 38543 38709
rect 39641 38663 39687 38709
rect 33684 38352 33730 38398
rect 33787 38352 33833 38398
rect 33890 38352 33936 38398
rect 33993 38352 34039 38398
rect 34096 38352 34142 38398
rect 34199 38352 34245 38398
rect 34302 38352 34348 38398
rect 34405 38352 34451 38398
rect 34508 38352 34554 38398
rect 34612 38352 34658 38398
rect 37909 38439 37955 38485
rect 38026 38439 38072 38485
rect 38143 38439 38189 38485
rect 38261 38439 38307 38485
rect 38379 38439 38425 38485
rect 38497 38439 38543 38485
rect 43739 38597 43785 38643
rect 43906 38597 43952 38643
rect 44071 38597 44117 38643
rect 44236 38597 44282 38643
rect 39641 38439 39687 38485
rect 50516 38611 50562 38657
rect 50703 38611 50749 38657
rect 50890 38611 50936 38657
rect 51076 38611 51122 38657
rect 51263 38611 51309 38657
rect 37909 38215 37955 38261
rect 38026 38215 38072 38261
rect 38143 38215 38189 38261
rect 38261 38215 38307 38261
rect 38379 38215 38425 38261
rect 38497 38215 38543 38261
rect 50467 38352 50513 38398
rect 50571 38352 50617 38398
rect 50674 38352 50720 38398
rect 50777 38352 50823 38398
rect 50880 38352 50926 38398
rect 50983 38352 51029 38398
rect 51086 38352 51132 38398
rect 51189 38352 51235 38398
rect 51292 38352 51338 38398
rect 51395 38352 51441 38398
rect 33684 38128 33730 38174
rect 33787 38128 33833 38174
rect 33890 38128 33936 38174
rect 33993 38128 34039 38174
rect 34096 38128 34142 38174
rect 34199 38128 34245 38174
rect 34302 38128 34348 38174
rect 34405 38128 34451 38174
rect 34508 38128 34554 38174
rect 34612 38128 34658 38174
rect 39740 38128 39786 38174
rect 39862 38128 39908 38174
rect 39985 38128 40031 38174
rect 40108 38128 40154 38174
rect 33684 37904 33730 37950
rect 33787 37904 33833 37950
rect 33890 37904 33936 37950
rect 33993 37904 34039 37950
rect 34096 37904 34142 37950
rect 34199 37904 34245 37950
rect 34302 37904 34348 37950
rect 34405 37904 34451 37950
rect 34508 37904 34554 37950
rect 34612 37904 34658 37950
rect 39740 37904 39786 37950
rect 39862 37904 39908 37950
rect 39985 37904 40031 37950
rect 40108 37904 40154 37950
rect 50467 38128 50513 38174
rect 50571 38128 50617 38174
rect 50674 38128 50720 38174
rect 50777 38128 50823 38174
rect 50880 38128 50926 38174
rect 50983 38128 51029 38174
rect 51086 38128 51132 38174
rect 51189 38128 51235 38174
rect 51292 38128 51338 38174
rect 51395 38128 51441 38174
rect 43739 37904 43785 37950
rect 43906 37904 43952 37950
rect 44071 37904 44117 37950
rect 44236 37904 44282 37950
rect 33684 37680 33730 37726
rect 33787 37680 33833 37726
rect 33890 37680 33936 37726
rect 33993 37680 34039 37726
rect 34096 37680 34142 37726
rect 34199 37680 34245 37726
rect 34302 37680 34348 37726
rect 34405 37680 34451 37726
rect 34508 37680 34554 37726
rect 34612 37680 34658 37726
rect 39740 37680 39786 37726
rect 39862 37680 39908 37726
rect 39985 37680 40031 37726
rect 40108 37680 40154 37726
rect 50467 37904 50513 37950
rect 50571 37904 50617 37950
rect 50674 37904 50720 37950
rect 50777 37904 50823 37950
rect 50880 37904 50926 37950
rect 50983 37904 51029 37950
rect 51086 37904 51132 37950
rect 51189 37904 51235 37950
rect 51292 37904 51338 37950
rect 51395 37904 51441 37950
rect 50467 37680 50513 37726
rect 50571 37680 50617 37726
rect 50674 37680 50720 37726
rect 50777 37680 50823 37726
rect 50880 37680 50926 37726
rect 50983 37680 51029 37726
rect 51086 37680 51132 37726
rect 51189 37680 51235 37726
rect 51292 37680 51338 37726
rect 51395 37680 51441 37726
rect 37909 37593 37955 37639
rect 38026 37593 38072 37639
rect 38143 37593 38189 37639
rect 38261 37593 38307 37639
rect 38379 37593 38425 37639
rect 38497 37593 38543 37639
rect 33684 37456 33730 37502
rect 33787 37456 33833 37502
rect 33890 37456 33936 37502
rect 33993 37456 34039 37502
rect 34096 37456 34142 37502
rect 34199 37456 34245 37502
rect 34302 37456 34348 37502
rect 34405 37456 34451 37502
rect 34508 37456 34554 37502
rect 34612 37456 34658 37502
rect 33816 37197 33862 37243
rect 34002 37197 34048 37243
rect 34189 37197 34235 37243
rect 34376 37197 34422 37243
rect 34562 37197 34608 37243
rect 37909 37369 37955 37415
rect 38026 37369 38072 37415
rect 38143 37369 38189 37415
rect 38261 37369 38307 37415
rect 38379 37369 38425 37415
rect 38497 37369 38543 37415
rect 39641 37369 39687 37415
rect 50467 37456 50513 37502
rect 50571 37456 50617 37502
rect 50674 37456 50720 37502
rect 50777 37456 50823 37502
rect 50880 37456 50926 37502
rect 50983 37456 51029 37502
rect 51086 37456 51132 37502
rect 51189 37456 51235 37502
rect 51292 37456 51338 37502
rect 51395 37456 51441 37502
rect 37909 37145 37955 37191
rect 38026 37145 38072 37191
rect 38143 37145 38189 37191
rect 38261 37145 38307 37191
rect 38379 37145 38425 37191
rect 38497 37145 38543 37191
rect 39641 37145 39687 37191
rect 43739 37211 43785 37257
rect 43906 37211 43952 37257
rect 44071 37211 44117 37257
rect 44236 37211 44282 37257
rect 50516 37197 50562 37243
rect 50703 37197 50749 37243
rect 50890 37197 50936 37243
rect 51076 37197 51122 37243
rect 51263 37197 51309 37243
rect 33816 36811 33862 36857
rect 34002 36811 34048 36857
rect 34189 36811 34235 36857
rect 34376 36811 34422 36857
rect 34562 36811 34608 36857
rect 37909 36863 37955 36909
rect 38026 36863 38072 36909
rect 38143 36863 38189 36909
rect 38261 36863 38307 36909
rect 38379 36863 38425 36909
rect 38497 36863 38543 36909
rect 39641 36863 39687 36909
rect 33684 36552 33730 36598
rect 33787 36552 33833 36598
rect 33890 36552 33936 36598
rect 33993 36552 34039 36598
rect 34096 36552 34142 36598
rect 34199 36552 34245 36598
rect 34302 36552 34348 36598
rect 34405 36552 34451 36598
rect 34508 36552 34554 36598
rect 34612 36552 34658 36598
rect 37909 36639 37955 36685
rect 38026 36639 38072 36685
rect 38143 36639 38189 36685
rect 38261 36639 38307 36685
rect 38379 36639 38425 36685
rect 38497 36639 38543 36685
rect 43739 36797 43785 36843
rect 43906 36797 43952 36843
rect 44071 36797 44117 36843
rect 44236 36797 44282 36843
rect 39641 36639 39687 36685
rect 50516 36811 50562 36857
rect 50703 36811 50749 36857
rect 50890 36811 50936 36857
rect 51076 36811 51122 36857
rect 51263 36811 51309 36857
rect 37909 36415 37955 36461
rect 38026 36415 38072 36461
rect 38143 36415 38189 36461
rect 38261 36415 38307 36461
rect 38379 36415 38425 36461
rect 38497 36415 38543 36461
rect 50467 36552 50513 36598
rect 50571 36552 50617 36598
rect 50674 36552 50720 36598
rect 50777 36552 50823 36598
rect 50880 36552 50926 36598
rect 50983 36552 51029 36598
rect 51086 36552 51132 36598
rect 51189 36552 51235 36598
rect 51292 36552 51338 36598
rect 51395 36552 51441 36598
rect 33684 36328 33730 36374
rect 33787 36328 33833 36374
rect 33890 36328 33936 36374
rect 33993 36328 34039 36374
rect 34096 36328 34142 36374
rect 34199 36328 34245 36374
rect 34302 36328 34348 36374
rect 34405 36328 34451 36374
rect 34508 36328 34554 36374
rect 34612 36328 34658 36374
rect 39740 36328 39786 36374
rect 39862 36328 39908 36374
rect 39985 36328 40031 36374
rect 40108 36328 40154 36374
rect 33684 36104 33730 36150
rect 33787 36104 33833 36150
rect 33890 36104 33936 36150
rect 33993 36104 34039 36150
rect 34096 36104 34142 36150
rect 34199 36104 34245 36150
rect 34302 36104 34348 36150
rect 34405 36104 34451 36150
rect 34508 36104 34554 36150
rect 34612 36104 34658 36150
rect 39740 36104 39786 36150
rect 39862 36104 39908 36150
rect 39985 36104 40031 36150
rect 40108 36104 40154 36150
rect 50467 36328 50513 36374
rect 50571 36328 50617 36374
rect 50674 36328 50720 36374
rect 50777 36328 50823 36374
rect 50880 36328 50926 36374
rect 50983 36328 51029 36374
rect 51086 36328 51132 36374
rect 51189 36328 51235 36374
rect 51292 36328 51338 36374
rect 51395 36328 51441 36374
rect 43739 36104 43785 36150
rect 43906 36104 43952 36150
rect 44071 36104 44117 36150
rect 44236 36104 44282 36150
rect 50467 36104 50513 36150
rect 50571 36104 50617 36150
rect 50674 36104 50720 36150
rect 50777 36104 50823 36150
rect 50880 36104 50926 36150
rect 50983 36104 51029 36150
rect 51086 36104 51132 36150
rect 51189 36104 51235 36150
rect 51292 36104 51338 36150
rect 51395 36104 51441 36150
<< mvpdiffc >>
rect 29317 65804 29363 65850
rect 29478 65804 29524 65850
rect 29638 65804 29684 65850
rect 29798 65804 29844 65850
rect 29959 65804 30005 65850
rect 30121 65804 30167 65850
rect 30284 65804 30330 65850
rect 35409 65772 37291 65818
rect 37348 65772 37394 65818
rect 37451 65772 37497 65818
rect 37554 65772 37600 65818
rect 37657 65772 37703 65818
rect 37760 65772 37806 65818
rect 37863 65772 37909 65818
rect 35409 65548 37291 65594
rect 37348 65548 37394 65594
rect 37451 65548 37497 65594
rect 37554 65548 37600 65594
rect 37657 65548 37703 65594
rect 37760 65548 37806 65594
rect 37863 65548 37909 65594
rect 38376 65548 38422 65594
rect 38479 65548 38525 65594
rect 38582 65548 38628 65594
rect 38686 65548 38732 65594
rect 38790 65548 38836 65594
rect 38894 65548 38940 65594
rect 38998 65548 39044 65594
rect 39102 65548 39148 65594
rect 39206 65548 39252 65594
rect 39310 65548 39356 65594
rect 39414 65548 39460 65594
rect 39518 65548 39564 65594
rect 39622 65548 39668 65594
rect 42676 65548 42722 65594
rect 42779 65548 42825 65594
rect 42882 65548 42928 65594
rect 42986 65548 43032 65594
rect 43090 65548 43136 65594
rect 43194 65548 43240 65594
rect 43298 65548 43344 65594
rect 43402 65548 43448 65594
rect 43506 65548 43552 65594
rect 43610 65548 43656 65594
rect 43714 65548 43760 65594
rect 43818 65548 43864 65594
rect 43922 65548 43968 65594
rect 47114 65772 48996 65818
rect 49053 65772 49099 65818
rect 49156 65772 49202 65818
rect 49259 65772 49305 65818
rect 49362 65772 49408 65818
rect 49465 65772 49511 65818
rect 49568 65772 49614 65818
rect 35409 65324 37291 65370
rect 37348 65324 37394 65370
rect 37451 65324 37497 65370
rect 37554 65324 37600 65370
rect 37657 65324 37703 65370
rect 37760 65324 37806 65370
rect 37863 65324 37909 65370
rect 38376 65324 38422 65370
rect 38479 65324 38525 65370
rect 38582 65324 38628 65370
rect 38686 65324 38732 65370
rect 38790 65324 38836 65370
rect 38894 65324 38940 65370
rect 38998 65324 39044 65370
rect 39102 65324 39148 65370
rect 39206 65324 39252 65370
rect 39310 65324 39356 65370
rect 39414 65324 39460 65370
rect 39518 65324 39564 65370
rect 39622 65324 39668 65370
rect 45346 65548 45392 65594
rect 45449 65548 45495 65594
rect 45552 65548 45598 65594
rect 45656 65548 45702 65594
rect 45760 65548 45806 65594
rect 45864 65548 45910 65594
rect 45968 65548 46014 65594
rect 46072 65548 46118 65594
rect 46176 65548 46222 65594
rect 46280 65548 46326 65594
rect 46384 65548 46430 65594
rect 46488 65548 46534 65594
rect 46592 65548 46638 65594
rect 47114 65548 48996 65594
rect 49053 65548 49099 65594
rect 49156 65548 49202 65594
rect 49259 65548 49305 65594
rect 49362 65548 49408 65594
rect 49465 65548 49511 65594
rect 49568 65548 49614 65594
rect 54793 65804 54839 65850
rect 54956 65804 55002 65850
rect 55118 65804 55164 65850
rect 55279 65804 55325 65850
rect 55439 65804 55485 65850
rect 55599 65804 55645 65850
rect 55760 65804 55806 65850
rect 42676 65324 42722 65370
rect 42779 65324 42825 65370
rect 42882 65324 42928 65370
rect 42986 65324 43032 65370
rect 43090 65324 43136 65370
rect 43194 65324 43240 65370
rect 43298 65324 43344 65370
rect 43402 65324 43448 65370
rect 43506 65324 43552 65370
rect 43610 65324 43656 65370
rect 43714 65324 43760 65370
rect 43818 65324 43864 65370
rect 43922 65324 43968 65370
rect 45346 65324 45392 65370
rect 45449 65324 45495 65370
rect 45552 65324 45598 65370
rect 45656 65324 45702 65370
rect 45760 65324 45806 65370
rect 45864 65324 45910 65370
rect 45968 65324 46014 65370
rect 46072 65324 46118 65370
rect 46176 65324 46222 65370
rect 46280 65324 46326 65370
rect 46384 65324 46430 65370
rect 46488 65324 46534 65370
rect 46592 65324 46638 65370
rect 47114 65324 48996 65370
rect 49053 65324 49099 65370
rect 49156 65324 49202 65370
rect 49259 65324 49305 65370
rect 49362 65324 49408 65370
rect 49465 65324 49511 65370
rect 49568 65324 49614 65370
rect 29317 64904 29363 64950
rect 29478 64904 29524 64950
rect 29638 64904 29684 64950
rect 29798 64904 29844 64950
rect 29959 64904 30005 64950
rect 30121 64904 30167 64950
rect 30284 64904 30330 64950
rect 31349 64904 33323 64950
rect 31349 64680 33323 64726
rect 31349 64456 33323 64502
rect 44812 64904 44858 64950
rect 44925 64904 44971 64950
rect 45038 64904 45084 64950
rect 45151 64904 45197 64950
rect 45264 64904 45310 64950
rect 51802 64904 53776 64950
rect 35273 64593 35523 64639
rect 35580 64593 35626 64639
rect 35683 64593 35729 64639
rect 35786 64593 35832 64639
rect 35889 64593 35935 64639
rect 35992 64593 36038 64639
rect 36095 64593 36141 64639
rect 36198 64593 36244 64639
rect 36301 64593 36347 64639
rect 36854 64593 36900 64639
rect 36971 64593 37017 64639
rect 37088 64593 37134 64639
rect 37206 64593 37252 64639
rect 37324 64593 37370 64639
rect 37442 64593 37488 64639
rect 44812 64680 44858 64726
rect 44925 64680 44971 64726
rect 45038 64680 45084 64726
rect 45151 64680 45197 64726
rect 45264 64680 45310 64726
rect 54793 64904 54839 64950
rect 54956 64904 55002 64950
rect 55118 64904 55164 64950
rect 55279 64904 55325 64950
rect 55439 64904 55485 64950
rect 55599 64904 55645 64950
rect 55760 64904 55806 64950
rect 31349 64232 33323 64278
rect 35273 64369 35523 64415
rect 35580 64369 35626 64415
rect 35683 64369 35729 64415
rect 35786 64369 35832 64415
rect 35889 64369 35935 64415
rect 35992 64369 36038 64415
rect 36095 64369 36141 64415
rect 36198 64369 36244 64415
rect 36301 64369 36347 64415
rect 48778 64593 48824 64639
rect 48881 64593 48927 64639
rect 48984 64593 49030 64639
rect 49087 64593 49133 64639
rect 49190 64593 49236 64639
rect 49293 64593 49339 64639
rect 49396 64593 49442 64639
rect 49499 64593 49545 64639
rect 49602 64593 49852 64639
rect 36854 64369 36900 64415
rect 36971 64369 37017 64415
rect 37088 64369 37134 64415
rect 37206 64369 37252 64415
rect 37324 64369 37370 64415
rect 37442 64369 37488 64415
rect 39021 64369 39067 64415
rect 39144 64369 39190 64415
rect 39267 64369 39313 64415
rect 44812 64456 44858 64502
rect 44925 64456 44971 64502
rect 45038 64456 45084 64502
rect 45151 64456 45197 64502
rect 45264 64456 45310 64502
rect 48778 64369 48824 64415
rect 48881 64369 48927 64415
rect 48984 64369 49030 64415
rect 49087 64369 49133 64415
rect 49190 64369 49236 64415
rect 49293 64369 49339 64415
rect 49396 64369 49442 64415
rect 49499 64369 49545 64415
rect 49602 64369 49852 64415
rect 35273 64145 35523 64191
rect 35580 64145 35626 64191
rect 35683 64145 35729 64191
rect 35786 64145 35832 64191
rect 35889 64145 35935 64191
rect 35992 64145 36038 64191
rect 36095 64145 36141 64191
rect 36198 64145 36244 64191
rect 36301 64145 36347 64191
rect 36854 64145 36900 64191
rect 36971 64145 37017 64191
rect 37088 64145 37134 64191
rect 37206 64145 37252 64191
rect 37324 64145 37370 64191
rect 37442 64145 37488 64191
rect 39021 64145 39067 64191
rect 39144 64145 39190 64191
rect 39267 64145 39313 64191
rect 44812 64232 44858 64278
rect 44925 64232 44971 64278
rect 45038 64232 45084 64278
rect 45151 64232 45197 64278
rect 45264 64232 45310 64278
rect 51802 64680 53776 64726
rect 51802 64456 53776 64502
rect 48778 64145 48824 64191
rect 48881 64145 48927 64191
rect 48984 64145 49030 64191
rect 49087 64145 49133 64191
rect 49190 64145 49236 64191
rect 49293 64145 49339 64191
rect 49396 64145 49442 64191
rect 49499 64145 49545 64191
rect 49602 64145 49852 64191
rect 51802 64232 53776 64278
rect 29317 64004 29363 64050
rect 29478 64004 29524 64050
rect 29638 64004 29684 64050
rect 29798 64004 29844 64050
rect 29959 64004 30005 64050
rect 30121 64004 30167 64050
rect 30284 64004 30330 64050
rect 54793 64004 54839 64050
rect 54956 64004 55002 64050
rect 55118 64004 55164 64050
rect 55279 64004 55325 64050
rect 55439 64004 55485 64050
rect 55599 64004 55645 64050
rect 55760 64004 55806 64050
rect 31349 63776 33323 63822
rect 35273 63863 35523 63909
rect 35580 63863 35626 63909
rect 35683 63863 35729 63909
rect 35786 63863 35832 63909
rect 35889 63863 35935 63909
rect 35992 63863 36038 63909
rect 36095 63863 36141 63909
rect 36198 63863 36244 63909
rect 36301 63863 36347 63909
rect 36854 63863 36900 63909
rect 36971 63863 37017 63909
rect 37088 63863 37134 63909
rect 37206 63863 37252 63909
rect 37324 63863 37370 63909
rect 37442 63863 37488 63909
rect 39021 63863 39067 63909
rect 39144 63863 39190 63909
rect 39267 63863 39313 63909
rect 31349 63552 33323 63598
rect 31349 63328 33323 63374
rect 29317 63104 29363 63150
rect 29478 63104 29524 63150
rect 29638 63104 29684 63150
rect 29798 63104 29844 63150
rect 29959 63104 30005 63150
rect 30121 63104 30167 63150
rect 30284 63104 30330 63150
rect 35273 63639 35523 63685
rect 35580 63639 35626 63685
rect 35683 63639 35729 63685
rect 35786 63639 35832 63685
rect 35889 63639 35935 63685
rect 35992 63639 36038 63685
rect 36095 63639 36141 63685
rect 36198 63639 36244 63685
rect 36301 63639 36347 63685
rect 36854 63639 36900 63685
rect 36971 63639 37017 63685
rect 37088 63639 37134 63685
rect 37206 63639 37252 63685
rect 37324 63639 37370 63685
rect 37442 63639 37488 63685
rect 48778 63863 48824 63909
rect 48881 63863 48927 63909
rect 48984 63863 49030 63909
rect 49087 63863 49133 63909
rect 49190 63863 49236 63909
rect 49293 63863 49339 63909
rect 49396 63863 49442 63909
rect 49499 63863 49545 63909
rect 49602 63863 49852 63909
rect 44812 63776 44858 63822
rect 44925 63776 44971 63822
rect 45038 63776 45084 63822
rect 45151 63776 45197 63822
rect 45264 63776 45310 63822
rect 39021 63639 39067 63685
rect 39144 63639 39190 63685
rect 39267 63639 39313 63685
rect 44812 63552 44858 63598
rect 44925 63552 44971 63598
rect 45038 63552 45084 63598
rect 45151 63552 45197 63598
rect 45264 63552 45310 63598
rect 48778 63639 48824 63685
rect 48881 63639 48927 63685
rect 48984 63639 49030 63685
rect 49087 63639 49133 63685
rect 49190 63639 49236 63685
rect 49293 63639 49339 63685
rect 49396 63639 49442 63685
rect 49499 63639 49545 63685
rect 49602 63639 49852 63685
rect 51802 63776 53776 63822
rect 35273 63415 35523 63461
rect 35580 63415 35626 63461
rect 35683 63415 35729 63461
rect 35786 63415 35832 63461
rect 35889 63415 35935 63461
rect 35992 63415 36038 63461
rect 36095 63415 36141 63461
rect 36198 63415 36244 63461
rect 36301 63415 36347 63461
rect 36854 63415 36900 63461
rect 36971 63415 37017 63461
rect 37088 63415 37134 63461
rect 37206 63415 37252 63461
rect 37324 63415 37370 63461
rect 37442 63415 37488 63461
rect 48778 63415 48824 63461
rect 48881 63415 48927 63461
rect 48984 63415 49030 63461
rect 49087 63415 49133 63461
rect 49190 63415 49236 63461
rect 49293 63415 49339 63461
rect 49396 63415 49442 63461
rect 49499 63415 49545 63461
rect 49602 63415 49852 63461
rect 44812 63328 44858 63374
rect 44925 63328 44971 63374
rect 45038 63328 45084 63374
rect 45151 63328 45197 63374
rect 45264 63328 45310 63374
rect 31349 63104 33323 63150
rect 31349 62880 33323 62926
rect 31349 62656 33323 62702
rect 51802 63552 53776 63598
rect 51802 63328 53776 63374
rect 44812 63104 44858 63150
rect 44925 63104 44971 63150
rect 45038 63104 45084 63150
rect 45151 63104 45197 63150
rect 45264 63104 45310 63150
rect 51802 63104 53776 63150
rect 35273 62793 35523 62839
rect 35580 62793 35626 62839
rect 35683 62793 35729 62839
rect 35786 62793 35832 62839
rect 35889 62793 35935 62839
rect 35992 62793 36038 62839
rect 36095 62793 36141 62839
rect 36198 62793 36244 62839
rect 36301 62793 36347 62839
rect 36854 62793 36900 62839
rect 36971 62793 37017 62839
rect 37088 62793 37134 62839
rect 37206 62793 37252 62839
rect 37324 62793 37370 62839
rect 37442 62793 37488 62839
rect 44812 62880 44858 62926
rect 44925 62880 44971 62926
rect 45038 62880 45084 62926
rect 45151 62880 45197 62926
rect 45264 62880 45310 62926
rect 54793 63104 54839 63150
rect 54956 63104 55002 63150
rect 55118 63104 55164 63150
rect 55279 63104 55325 63150
rect 55439 63104 55485 63150
rect 55599 63104 55645 63150
rect 55760 63104 55806 63150
rect 31349 62432 33323 62478
rect 35273 62569 35523 62615
rect 35580 62569 35626 62615
rect 35683 62569 35729 62615
rect 35786 62569 35832 62615
rect 35889 62569 35935 62615
rect 35992 62569 36038 62615
rect 36095 62569 36141 62615
rect 36198 62569 36244 62615
rect 36301 62569 36347 62615
rect 48778 62793 48824 62839
rect 48881 62793 48927 62839
rect 48984 62793 49030 62839
rect 49087 62793 49133 62839
rect 49190 62793 49236 62839
rect 49293 62793 49339 62839
rect 49396 62793 49442 62839
rect 49499 62793 49545 62839
rect 49602 62793 49852 62839
rect 36854 62569 36900 62615
rect 36971 62569 37017 62615
rect 37088 62569 37134 62615
rect 37206 62569 37252 62615
rect 37324 62569 37370 62615
rect 37442 62569 37488 62615
rect 39021 62569 39067 62615
rect 39144 62569 39190 62615
rect 39267 62569 39313 62615
rect 44812 62656 44858 62702
rect 44925 62656 44971 62702
rect 45038 62656 45084 62702
rect 45151 62656 45197 62702
rect 45264 62656 45310 62702
rect 48778 62569 48824 62615
rect 48881 62569 48927 62615
rect 48984 62569 49030 62615
rect 49087 62569 49133 62615
rect 49190 62569 49236 62615
rect 49293 62569 49339 62615
rect 49396 62569 49442 62615
rect 49499 62569 49545 62615
rect 49602 62569 49852 62615
rect 35273 62345 35523 62391
rect 35580 62345 35626 62391
rect 35683 62345 35729 62391
rect 35786 62345 35832 62391
rect 35889 62345 35935 62391
rect 35992 62345 36038 62391
rect 36095 62345 36141 62391
rect 36198 62345 36244 62391
rect 36301 62345 36347 62391
rect 36854 62345 36900 62391
rect 36971 62345 37017 62391
rect 37088 62345 37134 62391
rect 37206 62345 37252 62391
rect 37324 62345 37370 62391
rect 37442 62345 37488 62391
rect 39021 62345 39067 62391
rect 39144 62345 39190 62391
rect 39267 62345 39313 62391
rect 44812 62432 44858 62478
rect 44925 62432 44971 62478
rect 45038 62432 45084 62478
rect 45151 62432 45197 62478
rect 45264 62432 45310 62478
rect 51802 62880 53776 62926
rect 51802 62656 53776 62702
rect 48778 62345 48824 62391
rect 48881 62345 48927 62391
rect 48984 62345 49030 62391
rect 49087 62345 49133 62391
rect 49190 62345 49236 62391
rect 49293 62345 49339 62391
rect 49396 62345 49442 62391
rect 49499 62345 49545 62391
rect 49602 62345 49852 62391
rect 51802 62432 53776 62478
rect 29317 62204 29363 62250
rect 29478 62204 29524 62250
rect 29638 62204 29684 62250
rect 29798 62204 29844 62250
rect 29959 62204 30005 62250
rect 30121 62204 30167 62250
rect 30284 62204 30330 62250
rect 54793 62204 54839 62250
rect 54956 62204 55002 62250
rect 55118 62204 55164 62250
rect 55279 62204 55325 62250
rect 55439 62204 55485 62250
rect 55599 62204 55645 62250
rect 55760 62204 55806 62250
rect 31349 61976 33323 62022
rect 35273 62063 35523 62109
rect 35580 62063 35626 62109
rect 35683 62063 35729 62109
rect 35786 62063 35832 62109
rect 35889 62063 35935 62109
rect 35992 62063 36038 62109
rect 36095 62063 36141 62109
rect 36198 62063 36244 62109
rect 36301 62063 36347 62109
rect 36854 62063 36900 62109
rect 36971 62063 37017 62109
rect 37088 62063 37134 62109
rect 37206 62063 37252 62109
rect 37324 62063 37370 62109
rect 37442 62063 37488 62109
rect 39021 62063 39067 62109
rect 39144 62063 39190 62109
rect 39267 62063 39313 62109
rect 31349 61752 33323 61798
rect 31349 61528 33323 61574
rect 29317 61304 29363 61350
rect 29478 61304 29524 61350
rect 29638 61304 29684 61350
rect 29798 61304 29844 61350
rect 29959 61304 30005 61350
rect 30121 61304 30167 61350
rect 30284 61304 30330 61350
rect 35273 61839 35523 61885
rect 35580 61839 35626 61885
rect 35683 61839 35729 61885
rect 35786 61839 35832 61885
rect 35889 61839 35935 61885
rect 35992 61839 36038 61885
rect 36095 61839 36141 61885
rect 36198 61839 36244 61885
rect 36301 61839 36347 61885
rect 36854 61839 36900 61885
rect 36971 61839 37017 61885
rect 37088 61839 37134 61885
rect 37206 61839 37252 61885
rect 37324 61839 37370 61885
rect 37442 61839 37488 61885
rect 48778 62063 48824 62109
rect 48881 62063 48927 62109
rect 48984 62063 49030 62109
rect 49087 62063 49133 62109
rect 49190 62063 49236 62109
rect 49293 62063 49339 62109
rect 49396 62063 49442 62109
rect 49499 62063 49545 62109
rect 49602 62063 49852 62109
rect 44812 61976 44858 62022
rect 44925 61976 44971 62022
rect 45038 61976 45084 62022
rect 45151 61976 45197 62022
rect 45264 61976 45310 62022
rect 39021 61839 39067 61885
rect 39144 61839 39190 61885
rect 39267 61839 39313 61885
rect 44812 61752 44858 61798
rect 44925 61752 44971 61798
rect 45038 61752 45084 61798
rect 45151 61752 45197 61798
rect 45264 61752 45310 61798
rect 48778 61839 48824 61885
rect 48881 61839 48927 61885
rect 48984 61839 49030 61885
rect 49087 61839 49133 61885
rect 49190 61839 49236 61885
rect 49293 61839 49339 61885
rect 49396 61839 49442 61885
rect 49499 61839 49545 61885
rect 49602 61839 49852 61885
rect 51802 61976 53776 62022
rect 35273 61615 35523 61661
rect 35580 61615 35626 61661
rect 35683 61615 35729 61661
rect 35786 61615 35832 61661
rect 35889 61615 35935 61661
rect 35992 61615 36038 61661
rect 36095 61615 36141 61661
rect 36198 61615 36244 61661
rect 36301 61615 36347 61661
rect 36854 61615 36900 61661
rect 36971 61615 37017 61661
rect 37088 61615 37134 61661
rect 37206 61615 37252 61661
rect 37324 61615 37370 61661
rect 37442 61615 37488 61661
rect 48778 61615 48824 61661
rect 48881 61615 48927 61661
rect 48984 61615 49030 61661
rect 49087 61615 49133 61661
rect 49190 61615 49236 61661
rect 49293 61615 49339 61661
rect 49396 61615 49442 61661
rect 49499 61615 49545 61661
rect 49602 61615 49852 61661
rect 44812 61528 44858 61574
rect 44925 61528 44971 61574
rect 45038 61528 45084 61574
rect 45151 61528 45197 61574
rect 45264 61528 45310 61574
rect 31349 61304 33323 61350
rect 31349 61080 33323 61126
rect 31349 60856 33323 60902
rect 51802 61752 53776 61798
rect 51802 61528 53776 61574
rect 44812 61304 44858 61350
rect 44925 61304 44971 61350
rect 45038 61304 45084 61350
rect 45151 61304 45197 61350
rect 45264 61304 45310 61350
rect 51802 61304 53776 61350
rect 35273 60993 35523 61039
rect 35580 60993 35626 61039
rect 35683 60993 35729 61039
rect 35786 60993 35832 61039
rect 35889 60993 35935 61039
rect 35992 60993 36038 61039
rect 36095 60993 36141 61039
rect 36198 60993 36244 61039
rect 36301 60993 36347 61039
rect 36854 60993 36900 61039
rect 36971 60993 37017 61039
rect 37088 60993 37134 61039
rect 37206 60993 37252 61039
rect 37324 60993 37370 61039
rect 37442 60993 37488 61039
rect 44812 61080 44858 61126
rect 44925 61080 44971 61126
rect 45038 61080 45084 61126
rect 45151 61080 45197 61126
rect 45264 61080 45310 61126
rect 54793 61304 54839 61350
rect 54956 61304 55002 61350
rect 55118 61304 55164 61350
rect 55279 61304 55325 61350
rect 55439 61304 55485 61350
rect 55599 61304 55645 61350
rect 55760 61304 55806 61350
rect 31349 60632 33323 60678
rect 35273 60769 35523 60815
rect 35580 60769 35626 60815
rect 35683 60769 35729 60815
rect 35786 60769 35832 60815
rect 35889 60769 35935 60815
rect 35992 60769 36038 60815
rect 36095 60769 36141 60815
rect 36198 60769 36244 60815
rect 36301 60769 36347 60815
rect 48778 60993 48824 61039
rect 48881 60993 48927 61039
rect 48984 60993 49030 61039
rect 49087 60993 49133 61039
rect 49190 60993 49236 61039
rect 49293 60993 49339 61039
rect 49396 60993 49442 61039
rect 49499 60993 49545 61039
rect 49602 60993 49852 61039
rect 36854 60769 36900 60815
rect 36971 60769 37017 60815
rect 37088 60769 37134 60815
rect 37206 60769 37252 60815
rect 37324 60769 37370 60815
rect 37442 60769 37488 60815
rect 39021 60769 39067 60815
rect 39144 60769 39190 60815
rect 39267 60769 39313 60815
rect 44812 60856 44858 60902
rect 44925 60856 44971 60902
rect 45038 60856 45084 60902
rect 45151 60856 45197 60902
rect 45264 60856 45310 60902
rect 48778 60769 48824 60815
rect 48881 60769 48927 60815
rect 48984 60769 49030 60815
rect 49087 60769 49133 60815
rect 49190 60769 49236 60815
rect 49293 60769 49339 60815
rect 49396 60769 49442 60815
rect 49499 60769 49545 60815
rect 49602 60769 49852 60815
rect 35273 60545 35523 60591
rect 35580 60545 35626 60591
rect 35683 60545 35729 60591
rect 35786 60545 35832 60591
rect 35889 60545 35935 60591
rect 35992 60545 36038 60591
rect 36095 60545 36141 60591
rect 36198 60545 36244 60591
rect 36301 60545 36347 60591
rect 36854 60545 36900 60591
rect 36971 60545 37017 60591
rect 37088 60545 37134 60591
rect 37206 60545 37252 60591
rect 37324 60545 37370 60591
rect 37442 60545 37488 60591
rect 39021 60545 39067 60591
rect 39144 60545 39190 60591
rect 39267 60545 39313 60591
rect 44812 60632 44858 60678
rect 44925 60632 44971 60678
rect 45038 60632 45084 60678
rect 45151 60632 45197 60678
rect 45264 60632 45310 60678
rect 51802 61080 53776 61126
rect 51802 60856 53776 60902
rect 48778 60545 48824 60591
rect 48881 60545 48927 60591
rect 48984 60545 49030 60591
rect 49087 60545 49133 60591
rect 49190 60545 49236 60591
rect 49293 60545 49339 60591
rect 49396 60545 49442 60591
rect 49499 60545 49545 60591
rect 49602 60545 49852 60591
rect 51802 60632 53776 60678
rect 29317 60404 29363 60450
rect 29478 60404 29524 60450
rect 29638 60404 29684 60450
rect 29798 60404 29844 60450
rect 29959 60404 30005 60450
rect 30121 60404 30167 60450
rect 30284 60404 30330 60450
rect 54793 60404 54839 60450
rect 54956 60404 55002 60450
rect 55118 60404 55164 60450
rect 55279 60404 55325 60450
rect 55439 60404 55485 60450
rect 55599 60404 55645 60450
rect 55760 60404 55806 60450
rect 31349 60176 33323 60222
rect 35273 60263 35523 60309
rect 35580 60263 35626 60309
rect 35683 60263 35729 60309
rect 35786 60263 35832 60309
rect 35889 60263 35935 60309
rect 35992 60263 36038 60309
rect 36095 60263 36141 60309
rect 36198 60263 36244 60309
rect 36301 60263 36347 60309
rect 36854 60263 36900 60309
rect 36971 60263 37017 60309
rect 37088 60263 37134 60309
rect 37206 60263 37252 60309
rect 37324 60263 37370 60309
rect 37442 60263 37488 60309
rect 39021 60263 39067 60309
rect 39144 60263 39190 60309
rect 39267 60263 39313 60309
rect 31349 59952 33323 59998
rect 31349 59728 33323 59774
rect 29317 59504 29363 59550
rect 29478 59504 29524 59550
rect 29638 59504 29684 59550
rect 29798 59504 29844 59550
rect 29959 59504 30005 59550
rect 30121 59504 30167 59550
rect 30284 59504 30330 59550
rect 35273 60039 35523 60085
rect 35580 60039 35626 60085
rect 35683 60039 35729 60085
rect 35786 60039 35832 60085
rect 35889 60039 35935 60085
rect 35992 60039 36038 60085
rect 36095 60039 36141 60085
rect 36198 60039 36244 60085
rect 36301 60039 36347 60085
rect 36854 60039 36900 60085
rect 36971 60039 37017 60085
rect 37088 60039 37134 60085
rect 37206 60039 37252 60085
rect 37324 60039 37370 60085
rect 37442 60039 37488 60085
rect 48778 60263 48824 60309
rect 48881 60263 48927 60309
rect 48984 60263 49030 60309
rect 49087 60263 49133 60309
rect 49190 60263 49236 60309
rect 49293 60263 49339 60309
rect 49396 60263 49442 60309
rect 49499 60263 49545 60309
rect 49602 60263 49852 60309
rect 44812 60176 44858 60222
rect 44925 60176 44971 60222
rect 45038 60176 45084 60222
rect 45151 60176 45197 60222
rect 45264 60176 45310 60222
rect 39021 60039 39067 60085
rect 39144 60039 39190 60085
rect 39267 60039 39313 60085
rect 44812 59952 44858 59998
rect 44925 59952 44971 59998
rect 45038 59952 45084 59998
rect 45151 59952 45197 59998
rect 45264 59952 45310 59998
rect 48778 60039 48824 60085
rect 48881 60039 48927 60085
rect 48984 60039 49030 60085
rect 49087 60039 49133 60085
rect 49190 60039 49236 60085
rect 49293 60039 49339 60085
rect 49396 60039 49442 60085
rect 49499 60039 49545 60085
rect 49602 60039 49852 60085
rect 51802 60176 53776 60222
rect 35273 59815 35523 59861
rect 35580 59815 35626 59861
rect 35683 59815 35729 59861
rect 35786 59815 35832 59861
rect 35889 59815 35935 59861
rect 35992 59815 36038 59861
rect 36095 59815 36141 59861
rect 36198 59815 36244 59861
rect 36301 59815 36347 59861
rect 36854 59815 36900 59861
rect 36971 59815 37017 59861
rect 37088 59815 37134 59861
rect 37206 59815 37252 59861
rect 37324 59815 37370 59861
rect 37442 59815 37488 59861
rect 48778 59815 48824 59861
rect 48881 59815 48927 59861
rect 48984 59815 49030 59861
rect 49087 59815 49133 59861
rect 49190 59815 49236 59861
rect 49293 59815 49339 59861
rect 49396 59815 49442 59861
rect 49499 59815 49545 59861
rect 49602 59815 49852 59861
rect 44812 59728 44858 59774
rect 44925 59728 44971 59774
rect 45038 59728 45084 59774
rect 45151 59728 45197 59774
rect 45264 59728 45310 59774
rect 31349 59504 33323 59550
rect 31349 59280 33323 59326
rect 31349 59056 33323 59102
rect 51802 59952 53776 59998
rect 51802 59728 53776 59774
rect 44812 59504 44858 59550
rect 44925 59504 44971 59550
rect 45038 59504 45084 59550
rect 45151 59504 45197 59550
rect 45264 59504 45310 59550
rect 51802 59504 53776 59550
rect 35273 59193 35523 59239
rect 35580 59193 35626 59239
rect 35683 59193 35729 59239
rect 35786 59193 35832 59239
rect 35889 59193 35935 59239
rect 35992 59193 36038 59239
rect 36095 59193 36141 59239
rect 36198 59193 36244 59239
rect 36301 59193 36347 59239
rect 36854 59193 36900 59239
rect 36971 59193 37017 59239
rect 37088 59193 37134 59239
rect 37206 59193 37252 59239
rect 37324 59193 37370 59239
rect 37442 59193 37488 59239
rect 44812 59280 44858 59326
rect 44925 59280 44971 59326
rect 45038 59280 45084 59326
rect 45151 59280 45197 59326
rect 45264 59280 45310 59326
rect 54793 59504 54839 59550
rect 54956 59504 55002 59550
rect 55118 59504 55164 59550
rect 55279 59504 55325 59550
rect 55439 59504 55485 59550
rect 55599 59504 55645 59550
rect 55760 59504 55806 59550
rect 31349 58832 33323 58878
rect 35273 58969 35523 59015
rect 35580 58969 35626 59015
rect 35683 58969 35729 59015
rect 35786 58969 35832 59015
rect 35889 58969 35935 59015
rect 35992 58969 36038 59015
rect 36095 58969 36141 59015
rect 36198 58969 36244 59015
rect 36301 58969 36347 59015
rect 48778 59193 48824 59239
rect 48881 59193 48927 59239
rect 48984 59193 49030 59239
rect 49087 59193 49133 59239
rect 49190 59193 49236 59239
rect 49293 59193 49339 59239
rect 49396 59193 49442 59239
rect 49499 59193 49545 59239
rect 49602 59193 49852 59239
rect 36854 58969 36900 59015
rect 36971 58969 37017 59015
rect 37088 58969 37134 59015
rect 37206 58969 37252 59015
rect 37324 58969 37370 59015
rect 37442 58969 37488 59015
rect 39021 58969 39067 59015
rect 39144 58969 39190 59015
rect 39267 58969 39313 59015
rect 44812 59056 44858 59102
rect 44925 59056 44971 59102
rect 45038 59056 45084 59102
rect 45151 59056 45197 59102
rect 45264 59056 45310 59102
rect 48778 58969 48824 59015
rect 48881 58969 48927 59015
rect 48984 58969 49030 59015
rect 49087 58969 49133 59015
rect 49190 58969 49236 59015
rect 49293 58969 49339 59015
rect 49396 58969 49442 59015
rect 49499 58969 49545 59015
rect 49602 58969 49852 59015
rect 35273 58745 35523 58791
rect 35580 58745 35626 58791
rect 35683 58745 35729 58791
rect 35786 58745 35832 58791
rect 35889 58745 35935 58791
rect 35992 58745 36038 58791
rect 36095 58745 36141 58791
rect 36198 58745 36244 58791
rect 36301 58745 36347 58791
rect 36854 58745 36900 58791
rect 36971 58745 37017 58791
rect 37088 58745 37134 58791
rect 37206 58745 37252 58791
rect 37324 58745 37370 58791
rect 37442 58745 37488 58791
rect 39021 58745 39067 58791
rect 39144 58745 39190 58791
rect 39267 58745 39313 58791
rect 44812 58832 44858 58878
rect 44925 58832 44971 58878
rect 45038 58832 45084 58878
rect 45151 58832 45197 58878
rect 45264 58832 45310 58878
rect 51802 59280 53776 59326
rect 51802 59056 53776 59102
rect 48778 58745 48824 58791
rect 48881 58745 48927 58791
rect 48984 58745 49030 58791
rect 49087 58745 49133 58791
rect 49190 58745 49236 58791
rect 49293 58745 49339 58791
rect 49396 58745 49442 58791
rect 49499 58745 49545 58791
rect 49602 58745 49852 58791
rect 51802 58832 53776 58878
rect 29317 58604 29363 58650
rect 29478 58604 29524 58650
rect 29638 58604 29684 58650
rect 29798 58604 29844 58650
rect 29959 58604 30005 58650
rect 30121 58604 30167 58650
rect 30284 58604 30330 58650
rect 54793 58604 54839 58650
rect 54956 58604 55002 58650
rect 55118 58604 55164 58650
rect 55279 58604 55325 58650
rect 55439 58604 55485 58650
rect 55599 58604 55645 58650
rect 55760 58604 55806 58650
rect 31349 58376 33323 58422
rect 35273 58463 35523 58509
rect 35580 58463 35626 58509
rect 35683 58463 35729 58509
rect 35786 58463 35832 58509
rect 35889 58463 35935 58509
rect 35992 58463 36038 58509
rect 36095 58463 36141 58509
rect 36198 58463 36244 58509
rect 36301 58463 36347 58509
rect 36854 58463 36900 58509
rect 36971 58463 37017 58509
rect 37088 58463 37134 58509
rect 37206 58463 37252 58509
rect 37324 58463 37370 58509
rect 37442 58463 37488 58509
rect 39021 58463 39067 58509
rect 39144 58463 39190 58509
rect 39267 58463 39313 58509
rect 31349 58152 33323 58198
rect 31349 57928 33323 57974
rect 29317 57704 29363 57750
rect 29478 57704 29524 57750
rect 29638 57704 29684 57750
rect 29798 57704 29844 57750
rect 29959 57704 30005 57750
rect 30121 57704 30167 57750
rect 30284 57704 30330 57750
rect 35273 58239 35523 58285
rect 35580 58239 35626 58285
rect 35683 58239 35729 58285
rect 35786 58239 35832 58285
rect 35889 58239 35935 58285
rect 35992 58239 36038 58285
rect 36095 58239 36141 58285
rect 36198 58239 36244 58285
rect 36301 58239 36347 58285
rect 36854 58239 36900 58285
rect 36971 58239 37017 58285
rect 37088 58239 37134 58285
rect 37206 58239 37252 58285
rect 37324 58239 37370 58285
rect 37442 58239 37488 58285
rect 48778 58463 48824 58509
rect 48881 58463 48927 58509
rect 48984 58463 49030 58509
rect 49087 58463 49133 58509
rect 49190 58463 49236 58509
rect 49293 58463 49339 58509
rect 49396 58463 49442 58509
rect 49499 58463 49545 58509
rect 49602 58463 49852 58509
rect 44812 58376 44858 58422
rect 44925 58376 44971 58422
rect 45038 58376 45084 58422
rect 45151 58376 45197 58422
rect 45264 58376 45310 58422
rect 39021 58239 39067 58285
rect 39144 58239 39190 58285
rect 39267 58239 39313 58285
rect 44812 58152 44858 58198
rect 44925 58152 44971 58198
rect 45038 58152 45084 58198
rect 45151 58152 45197 58198
rect 45264 58152 45310 58198
rect 48778 58239 48824 58285
rect 48881 58239 48927 58285
rect 48984 58239 49030 58285
rect 49087 58239 49133 58285
rect 49190 58239 49236 58285
rect 49293 58239 49339 58285
rect 49396 58239 49442 58285
rect 49499 58239 49545 58285
rect 49602 58239 49852 58285
rect 51802 58376 53776 58422
rect 35273 58015 35523 58061
rect 35580 58015 35626 58061
rect 35683 58015 35729 58061
rect 35786 58015 35832 58061
rect 35889 58015 35935 58061
rect 35992 58015 36038 58061
rect 36095 58015 36141 58061
rect 36198 58015 36244 58061
rect 36301 58015 36347 58061
rect 36854 58015 36900 58061
rect 36971 58015 37017 58061
rect 37088 58015 37134 58061
rect 37206 58015 37252 58061
rect 37324 58015 37370 58061
rect 37442 58015 37488 58061
rect 48778 58015 48824 58061
rect 48881 58015 48927 58061
rect 48984 58015 49030 58061
rect 49087 58015 49133 58061
rect 49190 58015 49236 58061
rect 49293 58015 49339 58061
rect 49396 58015 49442 58061
rect 49499 58015 49545 58061
rect 49602 58015 49852 58061
rect 44812 57928 44858 57974
rect 44925 57928 44971 57974
rect 45038 57928 45084 57974
rect 45151 57928 45197 57974
rect 45264 57928 45310 57974
rect 31349 57704 33323 57750
rect 31349 57480 33323 57526
rect 31349 57256 33323 57302
rect 51802 58152 53776 58198
rect 51802 57928 53776 57974
rect 44812 57704 44858 57750
rect 44925 57704 44971 57750
rect 45038 57704 45084 57750
rect 45151 57704 45197 57750
rect 45264 57704 45310 57750
rect 51802 57704 53776 57750
rect 35273 57393 35523 57439
rect 35580 57393 35626 57439
rect 35683 57393 35729 57439
rect 35786 57393 35832 57439
rect 35889 57393 35935 57439
rect 35992 57393 36038 57439
rect 36095 57393 36141 57439
rect 36198 57393 36244 57439
rect 36301 57393 36347 57439
rect 36854 57393 36900 57439
rect 36971 57393 37017 57439
rect 37088 57393 37134 57439
rect 37206 57393 37252 57439
rect 37324 57393 37370 57439
rect 37442 57393 37488 57439
rect 44812 57480 44858 57526
rect 44925 57480 44971 57526
rect 45038 57480 45084 57526
rect 45151 57480 45197 57526
rect 45264 57480 45310 57526
rect 54793 57704 54839 57750
rect 54956 57704 55002 57750
rect 55118 57704 55164 57750
rect 55279 57704 55325 57750
rect 55439 57704 55485 57750
rect 55599 57704 55645 57750
rect 55760 57704 55806 57750
rect 31349 57032 33323 57078
rect 35273 57169 35523 57215
rect 35580 57169 35626 57215
rect 35683 57169 35729 57215
rect 35786 57169 35832 57215
rect 35889 57169 35935 57215
rect 35992 57169 36038 57215
rect 36095 57169 36141 57215
rect 36198 57169 36244 57215
rect 36301 57169 36347 57215
rect 48778 57393 48824 57439
rect 48881 57393 48927 57439
rect 48984 57393 49030 57439
rect 49087 57393 49133 57439
rect 49190 57393 49236 57439
rect 49293 57393 49339 57439
rect 49396 57393 49442 57439
rect 49499 57393 49545 57439
rect 49602 57393 49852 57439
rect 36854 57169 36900 57215
rect 36971 57169 37017 57215
rect 37088 57169 37134 57215
rect 37206 57169 37252 57215
rect 37324 57169 37370 57215
rect 37442 57169 37488 57215
rect 39021 57169 39067 57215
rect 39144 57169 39190 57215
rect 39267 57169 39313 57215
rect 44812 57256 44858 57302
rect 44925 57256 44971 57302
rect 45038 57256 45084 57302
rect 45151 57256 45197 57302
rect 45264 57256 45310 57302
rect 48778 57169 48824 57215
rect 48881 57169 48927 57215
rect 48984 57169 49030 57215
rect 49087 57169 49133 57215
rect 49190 57169 49236 57215
rect 49293 57169 49339 57215
rect 49396 57169 49442 57215
rect 49499 57169 49545 57215
rect 49602 57169 49852 57215
rect 35273 56945 35523 56991
rect 35580 56945 35626 56991
rect 35683 56945 35729 56991
rect 35786 56945 35832 56991
rect 35889 56945 35935 56991
rect 35992 56945 36038 56991
rect 36095 56945 36141 56991
rect 36198 56945 36244 56991
rect 36301 56945 36347 56991
rect 36854 56945 36900 56991
rect 36971 56945 37017 56991
rect 37088 56945 37134 56991
rect 37206 56945 37252 56991
rect 37324 56945 37370 56991
rect 37442 56945 37488 56991
rect 39021 56945 39067 56991
rect 39144 56945 39190 56991
rect 39267 56945 39313 56991
rect 44812 57032 44858 57078
rect 44925 57032 44971 57078
rect 45038 57032 45084 57078
rect 45151 57032 45197 57078
rect 45264 57032 45310 57078
rect 51802 57480 53776 57526
rect 51802 57256 53776 57302
rect 48778 56945 48824 56991
rect 48881 56945 48927 56991
rect 48984 56945 49030 56991
rect 49087 56945 49133 56991
rect 49190 56945 49236 56991
rect 49293 56945 49339 56991
rect 49396 56945 49442 56991
rect 49499 56945 49545 56991
rect 49602 56945 49852 56991
rect 51802 57032 53776 57078
rect 29317 56804 29363 56850
rect 29478 56804 29524 56850
rect 29638 56804 29684 56850
rect 29798 56804 29844 56850
rect 29959 56804 30005 56850
rect 30121 56804 30167 56850
rect 30284 56804 30330 56850
rect 54793 56804 54839 56850
rect 54956 56804 55002 56850
rect 55118 56804 55164 56850
rect 55279 56804 55325 56850
rect 55439 56804 55485 56850
rect 55599 56804 55645 56850
rect 55760 56804 55806 56850
rect 31349 56576 33323 56622
rect 35273 56663 35523 56709
rect 35580 56663 35626 56709
rect 35683 56663 35729 56709
rect 35786 56663 35832 56709
rect 35889 56663 35935 56709
rect 35992 56663 36038 56709
rect 36095 56663 36141 56709
rect 36198 56663 36244 56709
rect 36301 56663 36347 56709
rect 36854 56663 36900 56709
rect 36971 56663 37017 56709
rect 37088 56663 37134 56709
rect 37206 56663 37252 56709
rect 37324 56663 37370 56709
rect 37442 56663 37488 56709
rect 39021 56663 39067 56709
rect 39144 56663 39190 56709
rect 39267 56663 39313 56709
rect 31349 56352 33323 56398
rect 31349 56128 33323 56174
rect 29317 55904 29363 55950
rect 29478 55904 29524 55950
rect 29638 55904 29684 55950
rect 29798 55904 29844 55950
rect 29959 55904 30005 55950
rect 30121 55904 30167 55950
rect 30284 55904 30330 55950
rect 35273 56439 35523 56485
rect 35580 56439 35626 56485
rect 35683 56439 35729 56485
rect 35786 56439 35832 56485
rect 35889 56439 35935 56485
rect 35992 56439 36038 56485
rect 36095 56439 36141 56485
rect 36198 56439 36244 56485
rect 36301 56439 36347 56485
rect 36854 56439 36900 56485
rect 36971 56439 37017 56485
rect 37088 56439 37134 56485
rect 37206 56439 37252 56485
rect 37324 56439 37370 56485
rect 37442 56439 37488 56485
rect 48778 56663 48824 56709
rect 48881 56663 48927 56709
rect 48984 56663 49030 56709
rect 49087 56663 49133 56709
rect 49190 56663 49236 56709
rect 49293 56663 49339 56709
rect 49396 56663 49442 56709
rect 49499 56663 49545 56709
rect 49602 56663 49852 56709
rect 44812 56576 44858 56622
rect 44925 56576 44971 56622
rect 45038 56576 45084 56622
rect 45151 56576 45197 56622
rect 45264 56576 45310 56622
rect 39021 56439 39067 56485
rect 39144 56439 39190 56485
rect 39267 56439 39313 56485
rect 44812 56352 44858 56398
rect 44925 56352 44971 56398
rect 45038 56352 45084 56398
rect 45151 56352 45197 56398
rect 45264 56352 45310 56398
rect 48778 56439 48824 56485
rect 48881 56439 48927 56485
rect 48984 56439 49030 56485
rect 49087 56439 49133 56485
rect 49190 56439 49236 56485
rect 49293 56439 49339 56485
rect 49396 56439 49442 56485
rect 49499 56439 49545 56485
rect 49602 56439 49852 56485
rect 51802 56576 53776 56622
rect 35273 56215 35523 56261
rect 35580 56215 35626 56261
rect 35683 56215 35729 56261
rect 35786 56215 35832 56261
rect 35889 56215 35935 56261
rect 35992 56215 36038 56261
rect 36095 56215 36141 56261
rect 36198 56215 36244 56261
rect 36301 56215 36347 56261
rect 36854 56215 36900 56261
rect 36971 56215 37017 56261
rect 37088 56215 37134 56261
rect 37206 56215 37252 56261
rect 37324 56215 37370 56261
rect 37442 56215 37488 56261
rect 48778 56215 48824 56261
rect 48881 56215 48927 56261
rect 48984 56215 49030 56261
rect 49087 56215 49133 56261
rect 49190 56215 49236 56261
rect 49293 56215 49339 56261
rect 49396 56215 49442 56261
rect 49499 56215 49545 56261
rect 49602 56215 49852 56261
rect 44812 56128 44858 56174
rect 44925 56128 44971 56174
rect 45038 56128 45084 56174
rect 45151 56128 45197 56174
rect 45264 56128 45310 56174
rect 31349 55904 33323 55950
rect 31349 55680 33323 55726
rect 31349 55456 33323 55502
rect 51802 56352 53776 56398
rect 51802 56128 53776 56174
rect 44812 55904 44858 55950
rect 44925 55904 44971 55950
rect 45038 55904 45084 55950
rect 45151 55904 45197 55950
rect 45264 55904 45310 55950
rect 51802 55904 53776 55950
rect 35273 55593 35523 55639
rect 35580 55593 35626 55639
rect 35683 55593 35729 55639
rect 35786 55593 35832 55639
rect 35889 55593 35935 55639
rect 35992 55593 36038 55639
rect 36095 55593 36141 55639
rect 36198 55593 36244 55639
rect 36301 55593 36347 55639
rect 36854 55593 36900 55639
rect 36971 55593 37017 55639
rect 37088 55593 37134 55639
rect 37206 55593 37252 55639
rect 37324 55593 37370 55639
rect 37442 55593 37488 55639
rect 44812 55680 44858 55726
rect 44925 55680 44971 55726
rect 45038 55680 45084 55726
rect 45151 55680 45197 55726
rect 45264 55680 45310 55726
rect 54793 55904 54839 55950
rect 54956 55904 55002 55950
rect 55118 55904 55164 55950
rect 55279 55904 55325 55950
rect 55439 55904 55485 55950
rect 55599 55904 55645 55950
rect 55760 55904 55806 55950
rect 31349 55232 33323 55278
rect 35273 55369 35523 55415
rect 35580 55369 35626 55415
rect 35683 55369 35729 55415
rect 35786 55369 35832 55415
rect 35889 55369 35935 55415
rect 35992 55369 36038 55415
rect 36095 55369 36141 55415
rect 36198 55369 36244 55415
rect 36301 55369 36347 55415
rect 48778 55593 48824 55639
rect 48881 55593 48927 55639
rect 48984 55593 49030 55639
rect 49087 55593 49133 55639
rect 49190 55593 49236 55639
rect 49293 55593 49339 55639
rect 49396 55593 49442 55639
rect 49499 55593 49545 55639
rect 49602 55593 49852 55639
rect 36854 55369 36900 55415
rect 36971 55369 37017 55415
rect 37088 55369 37134 55415
rect 37206 55369 37252 55415
rect 37324 55369 37370 55415
rect 37442 55369 37488 55415
rect 39021 55369 39067 55415
rect 39144 55369 39190 55415
rect 39267 55369 39313 55415
rect 44812 55456 44858 55502
rect 44925 55456 44971 55502
rect 45038 55456 45084 55502
rect 45151 55456 45197 55502
rect 45264 55456 45310 55502
rect 48778 55369 48824 55415
rect 48881 55369 48927 55415
rect 48984 55369 49030 55415
rect 49087 55369 49133 55415
rect 49190 55369 49236 55415
rect 49293 55369 49339 55415
rect 49396 55369 49442 55415
rect 49499 55369 49545 55415
rect 49602 55369 49852 55415
rect 35273 55145 35523 55191
rect 35580 55145 35626 55191
rect 35683 55145 35729 55191
rect 35786 55145 35832 55191
rect 35889 55145 35935 55191
rect 35992 55145 36038 55191
rect 36095 55145 36141 55191
rect 36198 55145 36244 55191
rect 36301 55145 36347 55191
rect 36854 55145 36900 55191
rect 36971 55145 37017 55191
rect 37088 55145 37134 55191
rect 37206 55145 37252 55191
rect 37324 55145 37370 55191
rect 37442 55145 37488 55191
rect 39021 55145 39067 55191
rect 39144 55145 39190 55191
rect 39267 55145 39313 55191
rect 44812 55232 44858 55278
rect 44925 55232 44971 55278
rect 45038 55232 45084 55278
rect 45151 55232 45197 55278
rect 45264 55232 45310 55278
rect 51802 55680 53776 55726
rect 51802 55456 53776 55502
rect 48778 55145 48824 55191
rect 48881 55145 48927 55191
rect 48984 55145 49030 55191
rect 49087 55145 49133 55191
rect 49190 55145 49236 55191
rect 49293 55145 49339 55191
rect 49396 55145 49442 55191
rect 49499 55145 49545 55191
rect 49602 55145 49852 55191
rect 51802 55232 53776 55278
rect 29317 55004 29363 55050
rect 29478 55004 29524 55050
rect 29638 55004 29684 55050
rect 29798 55004 29844 55050
rect 29959 55004 30005 55050
rect 30121 55004 30167 55050
rect 30284 55004 30330 55050
rect 54793 55004 54839 55050
rect 54956 55004 55002 55050
rect 55118 55004 55164 55050
rect 55279 55004 55325 55050
rect 55439 55004 55485 55050
rect 55599 55004 55645 55050
rect 55760 55004 55806 55050
rect 31349 54776 33323 54822
rect 35273 54863 35523 54909
rect 35580 54863 35626 54909
rect 35683 54863 35729 54909
rect 35786 54863 35832 54909
rect 35889 54863 35935 54909
rect 35992 54863 36038 54909
rect 36095 54863 36141 54909
rect 36198 54863 36244 54909
rect 36301 54863 36347 54909
rect 36854 54863 36900 54909
rect 36971 54863 37017 54909
rect 37088 54863 37134 54909
rect 37206 54863 37252 54909
rect 37324 54863 37370 54909
rect 37442 54863 37488 54909
rect 39021 54863 39067 54909
rect 39144 54863 39190 54909
rect 39267 54863 39313 54909
rect 31349 54552 33323 54598
rect 31349 54328 33323 54374
rect 29317 54104 29363 54150
rect 29478 54104 29524 54150
rect 29638 54104 29684 54150
rect 29798 54104 29844 54150
rect 29959 54104 30005 54150
rect 30121 54104 30167 54150
rect 30284 54104 30330 54150
rect 35273 54639 35523 54685
rect 35580 54639 35626 54685
rect 35683 54639 35729 54685
rect 35786 54639 35832 54685
rect 35889 54639 35935 54685
rect 35992 54639 36038 54685
rect 36095 54639 36141 54685
rect 36198 54639 36244 54685
rect 36301 54639 36347 54685
rect 36854 54639 36900 54685
rect 36971 54639 37017 54685
rect 37088 54639 37134 54685
rect 37206 54639 37252 54685
rect 37324 54639 37370 54685
rect 37442 54639 37488 54685
rect 48778 54863 48824 54909
rect 48881 54863 48927 54909
rect 48984 54863 49030 54909
rect 49087 54863 49133 54909
rect 49190 54863 49236 54909
rect 49293 54863 49339 54909
rect 49396 54863 49442 54909
rect 49499 54863 49545 54909
rect 49602 54863 49852 54909
rect 44812 54776 44858 54822
rect 44925 54776 44971 54822
rect 45038 54776 45084 54822
rect 45151 54776 45197 54822
rect 45264 54776 45310 54822
rect 39021 54639 39067 54685
rect 39144 54639 39190 54685
rect 39267 54639 39313 54685
rect 44812 54552 44858 54598
rect 44925 54552 44971 54598
rect 45038 54552 45084 54598
rect 45151 54552 45197 54598
rect 45264 54552 45310 54598
rect 48778 54639 48824 54685
rect 48881 54639 48927 54685
rect 48984 54639 49030 54685
rect 49087 54639 49133 54685
rect 49190 54639 49236 54685
rect 49293 54639 49339 54685
rect 49396 54639 49442 54685
rect 49499 54639 49545 54685
rect 49602 54639 49852 54685
rect 51802 54776 53776 54822
rect 35273 54415 35523 54461
rect 35580 54415 35626 54461
rect 35683 54415 35729 54461
rect 35786 54415 35832 54461
rect 35889 54415 35935 54461
rect 35992 54415 36038 54461
rect 36095 54415 36141 54461
rect 36198 54415 36244 54461
rect 36301 54415 36347 54461
rect 36854 54415 36900 54461
rect 36971 54415 37017 54461
rect 37088 54415 37134 54461
rect 37206 54415 37252 54461
rect 37324 54415 37370 54461
rect 37442 54415 37488 54461
rect 48778 54415 48824 54461
rect 48881 54415 48927 54461
rect 48984 54415 49030 54461
rect 49087 54415 49133 54461
rect 49190 54415 49236 54461
rect 49293 54415 49339 54461
rect 49396 54415 49442 54461
rect 49499 54415 49545 54461
rect 49602 54415 49852 54461
rect 44812 54328 44858 54374
rect 44925 54328 44971 54374
rect 45038 54328 45084 54374
rect 45151 54328 45197 54374
rect 45264 54328 45310 54374
rect 31349 54104 33323 54150
rect 31349 53880 33323 53926
rect 31349 53656 33323 53702
rect 51802 54552 53776 54598
rect 51802 54328 53776 54374
rect 44812 54104 44858 54150
rect 44925 54104 44971 54150
rect 45038 54104 45084 54150
rect 45151 54104 45197 54150
rect 45264 54104 45310 54150
rect 51802 54104 53776 54150
rect 35273 53793 35523 53839
rect 35580 53793 35626 53839
rect 35683 53793 35729 53839
rect 35786 53793 35832 53839
rect 35889 53793 35935 53839
rect 35992 53793 36038 53839
rect 36095 53793 36141 53839
rect 36198 53793 36244 53839
rect 36301 53793 36347 53839
rect 36854 53793 36900 53839
rect 36971 53793 37017 53839
rect 37088 53793 37134 53839
rect 37206 53793 37252 53839
rect 37324 53793 37370 53839
rect 37442 53793 37488 53839
rect 44812 53880 44858 53926
rect 44925 53880 44971 53926
rect 45038 53880 45084 53926
rect 45151 53880 45197 53926
rect 45264 53880 45310 53926
rect 54793 54104 54839 54150
rect 54956 54104 55002 54150
rect 55118 54104 55164 54150
rect 55279 54104 55325 54150
rect 55439 54104 55485 54150
rect 55599 54104 55645 54150
rect 55760 54104 55806 54150
rect 31349 53432 33323 53478
rect 35273 53569 35523 53615
rect 35580 53569 35626 53615
rect 35683 53569 35729 53615
rect 35786 53569 35832 53615
rect 35889 53569 35935 53615
rect 35992 53569 36038 53615
rect 36095 53569 36141 53615
rect 36198 53569 36244 53615
rect 36301 53569 36347 53615
rect 48778 53793 48824 53839
rect 48881 53793 48927 53839
rect 48984 53793 49030 53839
rect 49087 53793 49133 53839
rect 49190 53793 49236 53839
rect 49293 53793 49339 53839
rect 49396 53793 49442 53839
rect 49499 53793 49545 53839
rect 49602 53793 49852 53839
rect 36854 53569 36900 53615
rect 36971 53569 37017 53615
rect 37088 53569 37134 53615
rect 37206 53569 37252 53615
rect 37324 53569 37370 53615
rect 37442 53569 37488 53615
rect 39021 53569 39067 53615
rect 39144 53569 39190 53615
rect 39267 53569 39313 53615
rect 44812 53656 44858 53702
rect 44925 53656 44971 53702
rect 45038 53656 45084 53702
rect 45151 53656 45197 53702
rect 45264 53656 45310 53702
rect 48778 53569 48824 53615
rect 48881 53569 48927 53615
rect 48984 53569 49030 53615
rect 49087 53569 49133 53615
rect 49190 53569 49236 53615
rect 49293 53569 49339 53615
rect 49396 53569 49442 53615
rect 49499 53569 49545 53615
rect 49602 53569 49852 53615
rect 35273 53345 35523 53391
rect 35580 53345 35626 53391
rect 35683 53345 35729 53391
rect 35786 53345 35832 53391
rect 35889 53345 35935 53391
rect 35992 53345 36038 53391
rect 36095 53345 36141 53391
rect 36198 53345 36244 53391
rect 36301 53345 36347 53391
rect 36854 53345 36900 53391
rect 36971 53345 37017 53391
rect 37088 53345 37134 53391
rect 37206 53345 37252 53391
rect 37324 53345 37370 53391
rect 37442 53345 37488 53391
rect 39021 53345 39067 53391
rect 39144 53345 39190 53391
rect 39267 53345 39313 53391
rect 44812 53432 44858 53478
rect 44925 53432 44971 53478
rect 45038 53432 45084 53478
rect 45151 53432 45197 53478
rect 45264 53432 45310 53478
rect 51802 53880 53776 53926
rect 51802 53656 53776 53702
rect 48778 53345 48824 53391
rect 48881 53345 48927 53391
rect 48984 53345 49030 53391
rect 49087 53345 49133 53391
rect 49190 53345 49236 53391
rect 49293 53345 49339 53391
rect 49396 53345 49442 53391
rect 49499 53345 49545 53391
rect 49602 53345 49852 53391
rect 51802 53432 53776 53478
rect 29317 53204 29363 53250
rect 29478 53204 29524 53250
rect 29638 53204 29684 53250
rect 29798 53204 29844 53250
rect 29959 53204 30005 53250
rect 30121 53204 30167 53250
rect 30284 53204 30330 53250
rect 54793 53204 54839 53250
rect 54956 53204 55002 53250
rect 55118 53204 55164 53250
rect 55279 53204 55325 53250
rect 55439 53204 55485 53250
rect 55599 53204 55645 53250
rect 55760 53204 55806 53250
rect 31349 52976 33323 53022
rect 35273 53063 35523 53109
rect 35580 53063 35626 53109
rect 35683 53063 35729 53109
rect 35786 53063 35832 53109
rect 35889 53063 35935 53109
rect 35992 53063 36038 53109
rect 36095 53063 36141 53109
rect 36198 53063 36244 53109
rect 36301 53063 36347 53109
rect 36854 53063 36900 53109
rect 36971 53063 37017 53109
rect 37088 53063 37134 53109
rect 37206 53063 37252 53109
rect 37324 53063 37370 53109
rect 37442 53063 37488 53109
rect 39021 53063 39067 53109
rect 39144 53063 39190 53109
rect 39267 53063 39313 53109
rect 31349 52752 33323 52798
rect 31349 52528 33323 52574
rect 29317 52304 29363 52350
rect 29478 52304 29524 52350
rect 29638 52304 29684 52350
rect 29798 52304 29844 52350
rect 29959 52304 30005 52350
rect 30121 52304 30167 52350
rect 30284 52304 30330 52350
rect 35273 52839 35523 52885
rect 35580 52839 35626 52885
rect 35683 52839 35729 52885
rect 35786 52839 35832 52885
rect 35889 52839 35935 52885
rect 35992 52839 36038 52885
rect 36095 52839 36141 52885
rect 36198 52839 36244 52885
rect 36301 52839 36347 52885
rect 36854 52839 36900 52885
rect 36971 52839 37017 52885
rect 37088 52839 37134 52885
rect 37206 52839 37252 52885
rect 37324 52839 37370 52885
rect 37442 52839 37488 52885
rect 48778 53063 48824 53109
rect 48881 53063 48927 53109
rect 48984 53063 49030 53109
rect 49087 53063 49133 53109
rect 49190 53063 49236 53109
rect 49293 53063 49339 53109
rect 49396 53063 49442 53109
rect 49499 53063 49545 53109
rect 49602 53063 49852 53109
rect 44812 52976 44858 53022
rect 44925 52976 44971 53022
rect 45038 52976 45084 53022
rect 45151 52976 45197 53022
rect 45264 52976 45310 53022
rect 39021 52839 39067 52885
rect 39144 52839 39190 52885
rect 39267 52839 39313 52885
rect 44812 52752 44858 52798
rect 44925 52752 44971 52798
rect 45038 52752 45084 52798
rect 45151 52752 45197 52798
rect 45264 52752 45310 52798
rect 48778 52839 48824 52885
rect 48881 52839 48927 52885
rect 48984 52839 49030 52885
rect 49087 52839 49133 52885
rect 49190 52839 49236 52885
rect 49293 52839 49339 52885
rect 49396 52839 49442 52885
rect 49499 52839 49545 52885
rect 49602 52839 49852 52885
rect 51802 52976 53776 53022
rect 35273 52615 35523 52661
rect 35580 52615 35626 52661
rect 35683 52615 35729 52661
rect 35786 52615 35832 52661
rect 35889 52615 35935 52661
rect 35992 52615 36038 52661
rect 36095 52615 36141 52661
rect 36198 52615 36244 52661
rect 36301 52615 36347 52661
rect 36854 52615 36900 52661
rect 36971 52615 37017 52661
rect 37088 52615 37134 52661
rect 37206 52615 37252 52661
rect 37324 52615 37370 52661
rect 37442 52615 37488 52661
rect 48778 52615 48824 52661
rect 48881 52615 48927 52661
rect 48984 52615 49030 52661
rect 49087 52615 49133 52661
rect 49190 52615 49236 52661
rect 49293 52615 49339 52661
rect 49396 52615 49442 52661
rect 49499 52615 49545 52661
rect 49602 52615 49852 52661
rect 44812 52528 44858 52574
rect 44925 52528 44971 52574
rect 45038 52528 45084 52574
rect 45151 52528 45197 52574
rect 45264 52528 45310 52574
rect 31349 52304 33323 52350
rect 31349 52080 33323 52126
rect 31349 51856 33323 51902
rect 51802 52752 53776 52798
rect 51802 52528 53776 52574
rect 44812 52304 44858 52350
rect 44925 52304 44971 52350
rect 45038 52304 45084 52350
rect 45151 52304 45197 52350
rect 45264 52304 45310 52350
rect 51802 52304 53776 52350
rect 35273 51993 35523 52039
rect 35580 51993 35626 52039
rect 35683 51993 35729 52039
rect 35786 51993 35832 52039
rect 35889 51993 35935 52039
rect 35992 51993 36038 52039
rect 36095 51993 36141 52039
rect 36198 51993 36244 52039
rect 36301 51993 36347 52039
rect 36854 51993 36900 52039
rect 36971 51993 37017 52039
rect 37088 51993 37134 52039
rect 37206 51993 37252 52039
rect 37324 51993 37370 52039
rect 37442 51993 37488 52039
rect 44812 52080 44858 52126
rect 44925 52080 44971 52126
rect 45038 52080 45084 52126
rect 45151 52080 45197 52126
rect 45264 52080 45310 52126
rect 54793 52304 54839 52350
rect 54956 52304 55002 52350
rect 55118 52304 55164 52350
rect 55279 52304 55325 52350
rect 55439 52304 55485 52350
rect 55599 52304 55645 52350
rect 55760 52304 55806 52350
rect 31349 51632 33323 51678
rect 35273 51769 35523 51815
rect 35580 51769 35626 51815
rect 35683 51769 35729 51815
rect 35786 51769 35832 51815
rect 35889 51769 35935 51815
rect 35992 51769 36038 51815
rect 36095 51769 36141 51815
rect 36198 51769 36244 51815
rect 36301 51769 36347 51815
rect 48778 51993 48824 52039
rect 48881 51993 48927 52039
rect 48984 51993 49030 52039
rect 49087 51993 49133 52039
rect 49190 51993 49236 52039
rect 49293 51993 49339 52039
rect 49396 51993 49442 52039
rect 49499 51993 49545 52039
rect 49602 51993 49852 52039
rect 36854 51769 36900 51815
rect 36971 51769 37017 51815
rect 37088 51769 37134 51815
rect 37206 51769 37252 51815
rect 37324 51769 37370 51815
rect 37442 51769 37488 51815
rect 39021 51769 39067 51815
rect 39144 51769 39190 51815
rect 39267 51769 39313 51815
rect 44812 51856 44858 51902
rect 44925 51856 44971 51902
rect 45038 51856 45084 51902
rect 45151 51856 45197 51902
rect 45264 51856 45310 51902
rect 48778 51769 48824 51815
rect 48881 51769 48927 51815
rect 48984 51769 49030 51815
rect 49087 51769 49133 51815
rect 49190 51769 49236 51815
rect 49293 51769 49339 51815
rect 49396 51769 49442 51815
rect 49499 51769 49545 51815
rect 49602 51769 49852 51815
rect 35273 51545 35523 51591
rect 35580 51545 35626 51591
rect 35683 51545 35729 51591
rect 35786 51545 35832 51591
rect 35889 51545 35935 51591
rect 35992 51545 36038 51591
rect 36095 51545 36141 51591
rect 36198 51545 36244 51591
rect 36301 51545 36347 51591
rect 36854 51545 36900 51591
rect 36971 51545 37017 51591
rect 37088 51545 37134 51591
rect 37206 51545 37252 51591
rect 37324 51545 37370 51591
rect 37442 51545 37488 51591
rect 39021 51545 39067 51591
rect 39144 51545 39190 51591
rect 39267 51545 39313 51591
rect 44812 51632 44858 51678
rect 44925 51632 44971 51678
rect 45038 51632 45084 51678
rect 45151 51632 45197 51678
rect 45264 51632 45310 51678
rect 51802 52080 53776 52126
rect 51802 51856 53776 51902
rect 48778 51545 48824 51591
rect 48881 51545 48927 51591
rect 48984 51545 49030 51591
rect 49087 51545 49133 51591
rect 49190 51545 49236 51591
rect 49293 51545 49339 51591
rect 49396 51545 49442 51591
rect 49499 51545 49545 51591
rect 49602 51545 49852 51591
rect 51802 51632 53776 51678
rect 29317 51404 29363 51450
rect 29478 51404 29524 51450
rect 29638 51404 29684 51450
rect 29798 51404 29844 51450
rect 29959 51404 30005 51450
rect 30121 51404 30167 51450
rect 30284 51404 30330 51450
rect 54793 51404 54839 51450
rect 54956 51404 55002 51450
rect 55118 51404 55164 51450
rect 55279 51404 55325 51450
rect 55439 51404 55485 51450
rect 55599 51404 55645 51450
rect 55760 51404 55806 51450
rect 31349 51176 33323 51222
rect 35273 51263 35523 51309
rect 35580 51263 35626 51309
rect 35683 51263 35729 51309
rect 35786 51263 35832 51309
rect 35889 51263 35935 51309
rect 35992 51263 36038 51309
rect 36095 51263 36141 51309
rect 36198 51263 36244 51309
rect 36301 51263 36347 51309
rect 36854 51263 36900 51309
rect 36971 51263 37017 51309
rect 37088 51263 37134 51309
rect 37206 51263 37252 51309
rect 37324 51263 37370 51309
rect 37442 51263 37488 51309
rect 39021 51263 39067 51309
rect 39144 51263 39190 51309
rect 39267 51263 39313 51309
rect 31349 50952 33323 50998
rect 31349 50728 33323 50774
rect 29317 50504 29363 50550
rect 29478 50504 29524 50550
rect 29638 50504 29684 50550
rect 29798 50504 29844 50550
rect 29959 50504 30005 50550
rect 30121 50504 30167 50550
rect 30284 50504 30330 50550
rect 35273 51039 35523 51085
rect 35580 51039 35626 51085
rect 35683 51039 35729 51085
rect 35786 51039 35832 51085
rect 35889 51039 35935 51085
rect 35992 51039 36038 51085
rect 36095 51039 36141 51085
rect 36198 51039 36244 51085
rect 36301 51039 36347 51085
rect 36854 51039 36900 51085
rect 36971 51039 37017 51085
rect 37088 51039 37134 51085
rect 37206 51039 37252 51085
rect 37324 51039 37370 51085
rect 37442 51039 37488 51085
rect 48778 51263 48824 51309
rect 48881 51263 48927 51309
rect 48984 51263 49030 51309
rect 49087 51263 49133 51309
rect 49190 51263 49236 51309
rect 49293 51263 49339 51309
rect 49396 51263 49442 51309
rect 49499 51263 49545 51309
rect 49602 51263 49852 51309
rect 44812 51176 44858 51222
rect 44925 51176 44971 51222
rect 45038 51176 45084 51222
rect 45151 51176 45197 51222
rect 45264 51176 45310 51222
rect 39021 51039 39067 51085
rect 39144 51039 39190 51085
rect 39267 51039 39313 51085
rect 44812 50952 44858 50998
rect 44925 50952 44971 50998
rect 45038 50952 45084 50998
rect 45151 50952 45197 50998
rect 45264 50952 45310 50998
rect 48778 51039 48824 51085
rect 48881 51039 48927 51085
rect 48984 51039 49030 51085
rect 49087 51039 49133 51085
rect 49190 51039 49236 51085
rect 49293 51039 49339 51085
rect 49396 51039 49442 51085
rect 49499 51039 49545 51085
rect 49602 51039 49852 51085
rect 51802 51176 53776 51222
rect 35273 50815 35523 50861
rect 35580 50815 35626 50861
rect 35683 50815 35729 50861
rect 35786 50815 35832 50861
rect 35889 50815 35935 50861
rect 35992 50815 36038 50861
rect 36095 50815 36141 50861
rect 36198 50815 36244 50861
rect 36301 50815 36347 50861
rect 36854 50815 36900 50861
rect 36971 50815 37017 50861
rect 37088 50815 37134 50861
rect 37206 50815 37252 50861
rect 37324 50815 37370 50861
rect 37442 50815 37488 50861
rect 48778 50815 48824 50861
rect 48881 50815 48927 50861
rect 48984 50815 49030 50861
rect 49087 50815 49133 50861
rect 49190 50815 49236 50861
rect 49293 50815 49339 50861
rect 49396 50815 49442 50861
rect 49499 50815 49545 50861
rect 49602 50815 49852 50861
rect 44812 50728 44858 50774
rect 44925 50728 44971 50774
rect 45038 50728 45084 50774
rect 45151 50728 45197 50774
rect 45264 50728 45310 50774
rect 31349 50504 33323 50550
rect 31349 50280 33323 50326
rect 31349 50056 33323 50102
rect 51802 50952 53776 50998
rect 51802 50728 53776 50774
rect 44812 50504 44858 50550
rect 44925 50504 44971 50550
rect 45038 50504 45084 50550
rect 45151 50504 45197 50550
rect 45264 50504 45310 50550
rect 51802 50504 53776 50550
rect 35273 50193 35523 50239
rect 35580 50193 35626 50239
rect 35683 50193 35729 50239
rect 35786 50193 35832 50239
rect 35889 50193 35935 50239
rect 35992 50193 36038 50239
rect 36095 50193 36141 50239
rect 36198 50193 36244 50239
rect 36301 50193 36347 50239
rect 36854 50193 36900 50239
rect 36971 50193 37017 50239
rect 37088 50193 37134 50239
rect 37206 50193 37252 50239
rect 37324 50193 37370 50239
rect 37442 50193 37488 50239
rect 44812 50280 44858 50326
rect 44925 50280 44971 50326
rect 45038 50280 45084 50326
rect 45151 50280 45197 50326
rect 45264 50280 45310 50326
rect 54793 50504 54839 50550
rect 54956 50504 55002 50550
rect 55118 50504 55164 50550
rect 55279 50504 55325 50550
rect 55439 50504 55485 50550
rect 55599 50504 55645 50550
rect 55760 50504 55806 50550
rect 31349 49832 33323 49878
rect 35273 49969 35523 50015
rect 35580 49969 35626 50015
rect 35683 49969 35729 50015
rect 35786 49969 35832 50015
rect 35889 49969 35935 50015
rect 35992 49969 36038 50015
rect 36095 49969 36141 50015
rect 36198 49969 36244 50015
rect 36301 49969 36347 50015
rect 48778 50193 48824 50239
rect 48881 50193 48927 50239
rect 48984 50193 49030 50239
rect 49087 50193 49133 50239
rect 49190 50193 49236 50239
rect 49293 50193 49339 50239
rect 49396 50193 49442 50239
rect 49499 50193 49545 50239
rect 49602 50193 49852 50239
rect 36854 49969 36900 50015
rect 36971 49969 37017 50015
rect 37088 49969 37134 50015
rect 37206 49969 37252 50015
rect 37324 49969 37370 50015
rect 37442 49969 37488 50015
rect 39021 49969 39067 50015
rect 39144 49969 39190 50015
rect 39267 49969 39313 50015
rect 44812 50056 44858 50102
rect 44925 50056 44971 50102
rect 45038 50056 45084 50102
rect 45151 50056 45197 50102
rect 45264 50056 45310 50102
rect 48778 49969 48824 50015
rect 48881 49969 48927 50015
rect 48984 49969 49030 50015
rect 49087 49969 49133 50015
rect 49190 49969 49236 50015
rect 49293 49969 49339 50015
rect 49396 49969 49442 50015
rect 49499 49969 49545 50015
rect 49602 49969 49852 50015
rect 35273 49745 35523 49791
rect 35580 49745 35626 49791
rect 35683 49745 35729 49791
rect 35786 49745 35832 49791
rect 35889 49745 35935 49791
rect 35992 49745 36038 49791
rect 36095 49745 36141 49791
rect 36198 49745 36244 49791
rect 36301 49745 36347 49791
rect 36854 49745 36900 49791
rect 36971 49745 37017 49791
rect 37088 49745 37134 49791
rect 37206 49745 37252 49791
rect 37324 49745 37370 49791
rect 37442 49745 37488 49791
rect 39021 49745 39067 49791
rect 39144 49745 39190 49791
rect 39267 49745 39313 49791
rect 44812 49832 44858 49878
rect 44925 49832 44971 49878
rect 45038 49832 45084 49878
rect 45151 49832 45197 49878
rect 45264 49832 45310 49878
rect 51802 50280 53776 50326
rect 51802 50056 53776 50102
rect 48778 49745 48824 49791
rect 48881 49745 48927 49791
rect 48984 49745 49030 49791
rect 49087 49745 49133 49791
rect 49190 49745 49236 49791
rect 49293 49745 49339 49791
rect 49396 49745 49442 49791
rect 49499 49745 49545 49791
rect 49602 49745 49852 49791
rect 51802 49832 53776 49878
rect 29317 49604 29363 49650
rect 29478 49604 29524 49650
rect 29638 49604 29684 49650
rect 29798 49604 29844 49650
rect 29959 49604 30005 49650
rect 30121 49604 30167 49650
rect 30284 49604 30330 49650
rect 54793 49604 54839 49650
rect 54956 49604 55002 49650
rect 55118 49604 55164 49650
rect 55279 49604 55325 49650
rect 55439 49604 55485 49650
rect 55599 49604 55645 49650
rect 55760 49604 55806 49650
rect 31349 49376 33323 49422
rect 35273 49463 35523 49509
rect 35580 49463 35626 49509
rect 35683 49463 35729 49509
rect 35786 49463 35832 49509
rect 35889 49463 35935 49509
rect 35992 49463 36038 49509
rect 36095 49463 36141 49509
rect 36198 49463 36244 49509
rect 36301 49463 36347 49509
rect 36854 49463 36900 49509
rect 36971 49463 37017 49509
rect 37088 49463 37134 49509
rect 37206 49463 37252 49509
rect 37324 49463 37370 49509
rect 37442 49463 37488 49509
rect 39021 49463 39067 49509
rect 39144 49463 39190 49509
rect 39267 49463 39313 49509
rect 31349 49152 33323 49198
rect 31349 48928 33323 48974
rect 29317 48704 29363 48750
rect 29478 48704 29524 48750
rect 29638 48704 29684 48750
rect 29798 48704 29844 48750
rect 29959 48704 30005 48750
rect 30121 48704 30167 48750
rect 30284 48704 30330 48750
rect 35273 49239 35523 49285
rect 35580 49239 35626 49285
rect 35683 49239 35729 49285
rect 35786 49239 35832 49285
rect 35889 49239 35935 49285
rect 35992 49239 36038 49285
rect 36095 49239 36141 49285
rect 36198 49239 36244 49285
rect 36301 49239 36347 49285
rect 36854 49239 36900 49285
rect 36971 49239 37017 49285
rect 37088 49239 37134 49285
rect 37206 49239 37252 49285
rect 37324 49239 37370 49285
rect 37442 49239 37488 49285
rect 48778 49463 48824 49509
rect 48881 49463 48927 49509
rect 48984 49463 49030 49509
rect 49087 49463 49133 49509
rect 49190 49463 49236 49509
rect 49293 49463 49339 49509
rect 49396 49463 49442 49509
rect 49499 49463 49545 49509
rect 49602 49463 49852 49509
rect 44812 49376 44858 49422
rect 44925 49376 44971 49422
rect 45038 49376 45084 49422
rect 45151 49376 45197 49422
rect 45264 49376 45310 49422
rect 39021 49239 39067 49285
rect 39144 49239 39190 49285
rect 39267 49239 39313 49285
rect 44812 49152 44858 49198
rect 44925 49152 44971 49198
rect 45038 49152 45084 49198
rect 45151 49152 45197 49198
rect 45264 49152 45310 49198
rect 48778 49239 48824 49285
rect 48881 49239 48927 49285
rect 48984 49239 49030 49285
rect 49087 49239 49133 49285
rect 49190 49239 49236 49285
rect 49293 49239 49339 49285
rect 49396 49239 49442 49285
rect 49499 49239 49545 49285
rect 49602 49239 49852 49285
rect 51802 49376 53776 49422
rect 35273 49015 35523 49061
rect 35580 49015 35626 49061
rect 35683 49015 35729 49061
rect 35786 49015 35832 49061
rect 35889 49015 35935 49061
rect 35992 49015 36038 49061
rect 36095 49015 36141 49061
rect 36198 49015 36244 49061
rect 36301 49015 36347 49061
rect 36854 49015 36900 49061
rect 36971 49015 37017 49061
rect 37088 49015 37134 49061
rect 37206 49015 37252 49061
rect 37324 49015 37370 49061
rect 37442 49015 37488 49061
rect 48778 49015 48824 49061
rect 48881 49015 48927 49061
rect 48984 49015 49030 49061
rect 49087 49015 49133 49061
rect 49190 49015 49236 49061
rect 49293 49015 49339 49061
rect 49396 49015 49442 49061
rect 49499 49015 49545 49061
rect 49602 49015 49852 49061
rect 44812 48928 44858 48974
rect 44925 48928 44971 48974
rect 45038 48928 45084 48974
rect 45151 48928 45197 48974
rect 45264 48928 45310 48974
rect 31349 48704 33323 48750
rect 31349 48480 33323 48526
rect 31349 48256 33323 48302
rect 51802 49152 53776 49198
rect 51802 48928 53776 48974
rect 44812 48704 44858 48750
rect 44925 48704 44971 48750
rect 45038 48704 45084 48750
rect 45151 48704 45197 48750
rect 45264 48704 45310 48750
rect 51802 48704 53776 48750
rect 35273 48393 35523 48439
rect 35580 48393 35626 48439
rect 35683 48393 35729 48439
rect 35786 48393 35832 48439
rect 35889 48393 35935 48439
rect 35992 48393 36038 48439
rect 36095 48393 36141 48439
rect 36198 48393 36244 48439
rect 36301 48393 36347 48439
rect 36854 48393 36900 48439
rect 36971 48393 37017 48439
rect 37088 48393 37134 48439
rect 37206 48393 37252 48439
rect 37324 48393 37370 48439
rect 37442 48393 37488 48439
rect 44812 48480 44858 48526
rect 44925 48480 44971 48526
rect 45038 48480 45084 48526
rect 45151 48480 45197 48526
rect 45264 48480 45310 48526
rect 54793 48704 54839 48750
rect 54956 48704 55002 48750
rect 55118 48704 55164 48750
rect 55279 48704 55325 48750
rect 55439 48704 55485 48750
rect 55599 48704 55645 48750
rect 55760 48704 55806 48750
rect 31349 48032 33323 48078
rect 35273 48169 35523 48215
rect 35580 48169 35626 48215
rect 35683 48169 35729 48215
rect 35786 48169 35832 48215
rect 35889 48169 35935 48215
rect 35992 48169 36038 48215
rect 36095 48169 36141 48215
rect 36198 48169 36244 48215
rect 36301 48169 36347 48215
rect 48778 48393 48824 48439
rect 48881 48393 48927 48439
rect 48984 48393 49030 48439
rect 49087 48393 49133 48439
rect 49190 48393 49236 48439
rect 49293 48393 49339 48439
rect 49396 48393 49442 48439
rect 49499 48393 49545 48439
rect 49602 48393 49852 48439
rect 36854 48169 36900 48215
rect 36971 48169 37017 48215
rect 37088 48169 37134 48215
rect 37206 48169 37252 48215
rect 37324 48169 37370 48215
rect 37442 48169 37488 48215
rect 39021 48169 39067 48215
rect 39144 48169 39190 48215
rect 39267 48169 39313 48215
rect 44812 48256 44858 48302
rect 44925 48256 44971 48302
rect 45038 48256 45084 48302
rect 45151 48256 45197 48302
rect 45264 48256 45310 48302
rect 48778 48169 48824 48215
rect 48881 48169 48927 48215
rect 48984 48169 49030 48215
rect 49087 48169 49133 48215
rect 49190 48169 49236 48215
rect 49293 48169 49339 48215
rect 49396 48169 49442 48215
rect 49499 48169 49545 48215
rect 49602 48169 49852 48215
rect 35273 47945 35523 47991
rect 35580 47945 35626 47991
rect 35683 47945 35729 47991
rect 35786 47945 35832 47991
rect 35889 47945 35935 47991
rect 35992 47945 36038 47991
rect 36095 47945 36141 47991
rect 36198 47945 36244 47991
rect 36301 47945 36347 47991
rect 36854 47945 36900 47991
rect 36971 47945 37017 47991
rect 37088 47945 37134 47991
rect 37206 47945 37252 47991
rect 37324 47945 37370 47991
rect 37442 47945 37488 47991
rect 39021 47945 39067 47991
rect 39144 47945 39190 47991
rect 39267 47945 39313 47991
rect 44812 48032 44858 48078
rect 44925 48032 44971 48078
rect 45038 48032 45084 48078
rect 45151 48032 45197 48078
rect 45264 48032 45310 48078
rect 51802 48480 53776 48526
rect 51802 48256 53776 48302
rect 48778 47945 48824 47991
rect 48881 47945 48927 47991
rect 48984 47945 49030 47991
rect 49087 47945 49133 47991
rect 49190 47945 49236 47991
rect 49293 47945 49339 47991
rect 49396 47945 49442 47991
rect 49499 47945 49545 47991
rect 49602 47945 49852 47991
rect 51802 48032 53776 48078
rect 29317 47804 29363 47850
rect 29478 47804 29524 47850
rect 29638 47804 29684 47850
rect 29798 47804 29844 47850
rect 29959 47804 30005 47850
rect 30121 47804 30167 47850
rect 30284 47804 30330 47850
rect 54793 47804 54839 47850
rect 54956 47804 55002 47850
rect 55118 47804 55164 47850
rect 55279 47804 55325 47850
rect 55439 47804 55485 47850
rect 55599 47804 55645 47850
rect 55760 47804 55806 47850
rect 31349 47576 33323 47622
rect 35273 47663 35523 47709
rect 35580 47663 35626 47709
rect 35683 47663 35729 47709
rect 35786 47663 35832 47709
rect 35889 47663 35935 47709
rect 35992 47663 36038 47709
rect 36095 47663 36141 47709
rect 36198 47663 36244 47709
rect 36301 47663 36347 47709
rect 36854 47663 36900 47709
rect 36971 47663 37017 47709
rect 37088 47663 37134 47709
rect 37206 47663 37252 47709
rect 37324 47663 37370 47709
rect 37442 47663 37488 47709
rect 39021 47663 39067 47709
rect 39144 47663 39190 47709
rect 39267 47663 39313 47709
rect 31349 47352 33323 47398
rect 31349 47128 33323 47174
rect 29317 46904 29363 46950
rect 29478 46904 29524 46950
rect 29638 46904 29684 46950
rect 29798 46904 29844 46950
rect 29959 46904 30005 46950
rect 30121 46904 30167 46950
rect 30284 46904 30330 46950
rect 35273 47439 35523 47485
rect 35580 47439 35626 47485
rect 35683 47439 35729 47485
rect 35786 47439 35832 47485
rect 35889 47439 35935 47485
rect 35992 47439 36038 47485
rect 36095 47439 36141 47485
rect 36198 47439 36244 47485
rect 36301 47439 36347 47485
rect 36854 47439 36900 47485
rect 36971 47439 37017 47485
rect 37088 47439 37134 47485
rect 37206 47439 37252 47485
rect 37324 47439 37370 47485
rect 37442 47439 37488 47485
rect 48778 47663 48824 47709
rect 48881 47663 48927 47709
rect 48984 47663 49030 47709
rect 49087 47663 49133 47709
rect 49190 47663 49236 47709
rect 49293 47663 49339 47709
rect 49396 47663 49442 47709
rect 49499 47663 49545 47709
rect 49602 47663 49852 47709
rect 44812 47576 44858 47622
rect 44925 47576 44971 47622
rect 45038 47576 45084 47622
rect 45151 47576 45197 47622
rect 45264 47576 45310 47622
rect 39021 47439 39067 47485
rect 39144 47439 39190 47485
rect 39267 47439 39313 47485
rect 44812 47352 44858 47398
rect 44925 47352 44971 47398
rect 45038 47352 45084 47398
rect 45151 47352 45197 47398
rect 45264 47352 45310 47398
rect 48778 47439 48824 47485
rect 48881 47439 48927 47485
rect 48984 47439 49030 47485
rect 49087 47439 49133 47485
rect 49190 47439 49236 47485
rect 49293 47439 49339 47485
rect 49396 47439 49442 47485
rect 49499 47439 49545 47485
rect 49602 47439 49852 47485
rect 51802 47576 53776 47622
rect 35273 47215 35523 47261
rect 35580 47215 35626 47261
rect 35683 47215 35729 47261
rect 35786 47215 35832 47261
rect 35889 47215 35935 47261
rect 35992 47215 36038 47261
rect 36095 47215 36141 47261
rect 36198 47215 36244 47261
rect 36301 47215 36347 47261
rect 36854 47215 36900 47261
rect 36971 47215 37017 47261
rect 37088 47215 37134 47261
rect 37206 47215 37252 47261
rect 37324 47215 37370 47261
rect 37442 47215 37488 47261
rect 48778 47215 48824 47261
rect 48881 47215 48927 47261
rect 48984 47215 49030 47261
rect 49087 47215 49133 47261
rect 49190 47215 49236 47261
rect 49293 47215 49339 47261
rect 49396 47215 49442 47261
rect 49499 47215 49545 47261
rect 49602 47215 49852 47261
rect 44812 47128 44858 47174
rect 44925 47128 44971 47174
rect 45038 47128 45084 47174
rect 45151 47128 45197 47174
rect 45264 47128 45310 47174
rect 31349 46904 33323 46950
rect 31349 46680 33323 46726
rect 31349 46456 33323 46502
rect 51802 47352 53776 47398
rect 51802 47128 53776 47174
rect 44812 46904 44858 46950
rect 44925 46904 44971 46950
rect 45038 46904 45084 46950
rect 45151 46904 45197 46950
rect 45264 46904 45310 46950
rect 51802 46904 53776 46950
rect 35273 46593 35523 46639
rect 35580 46593 35626 46639
rect 35683 46593 35729 46639
rect 35786 46593 35832 46639
rect 35889 46593 35935 46639
rect 35992 46593 36038 46639
rect 36095 46593 36141 46639
rect 36198 46593 36244 46639
rect 36301 46593 36347 46639
rect 36854 46593 36900 46639
rect 36971 46593 37017 46639
rect 37088 46593 37134 46639
rect 37206 46593 37252 46639
rect 37324 46593 37370 46639
rect 37442 46593 37488 46639
rect 44812 46680 44858 46726
rect 44925 46680 44971 46726
rect 45038 46680 45084 46726
rect 45151 46680 45197 46726
rect 45264 46680 45310 46726
rect 54793 46904 54839 46950
rect 54956 46904 55002 46950
rect 55118 46904 55164 46950
rect 55279 46904 55325 46950
rect 55439 46904 55485 46950
rect 55599 46904 55645 46950
rect 55760 46904 55806 46950
rect 31349 46232 33323 46278
rect 35273 46369 35523 46415
rect 35580 46369 35626 46415
rect 35683 46369 35729 46415
rect 35786 46369 35832 46415
rect 35889 46369 35935 46415
rect 35992 46369 36038 46415
rect 36095 46369 36141 46415
rect 36198 46369 36244 46415
rect 36301 46369 36347 46415
rect 48778 46593 48824 46639
rect 48881 46593 48927 46639
rect 48984 46593 49030 46639
rect 49087 46593 49133 46639
rect 49190 46593 49236 46639
rect 49293 46593 49339 46639
rect 49396 46593 49442 46639
rect 49499 46593 49545 46639
rect 49602 46593 49852 46639
rect 36854 46369 36900 46415
rect 36971 46369 37017 46415
rect 37088 46369 37134 46415
rect 37206 46369 37252 46415
rect 37324 46369 37370 46415
rect 37442 46369 37488 46415
rect 39021 46369 39067 46415
rect 39144 46369 39190 46415
rect 39267 46369 39313 46415
rect 44812 46456 44858 46502
rect 44925 46456 44971 46502
rect 45038 46456 45084 46502
rect 45151 46456 45197 46502
rect 45264 46456 45310 46502
rect 48778 46369 48824 46415
rect 48881 46369 48927 46415
rect 48984 46369 49030 46415
rect 49087 46369 49133 46415
rect 49190 46369 49236 46415
rect 49293 46369 49339 46415
rect 49396 46369 49442 46415
rect 49499 46369 49545 46415
rect 49602 46369 49852 46415
rect 35273 46145 35523 46191
rect 35580 46145 35626 46191
rect 35683 46145 35729 46191
rect 35786 46145 35832 46191
rect 35889 46145 35935 46191
rect 35992 46145 36038 46191
rect 36095 46145 36141 46191
rect 36198 46145 36244 46191
rect 36301 46145 36347 46191
rect 36854 46145 36900 46191
rect 36971 46145 37017 46191
rect 37088 46145 37134 46191
rect 37206 46145 37252 46191
rect 37324 46145 37370 46191
rect 37442 46145 37488 46191
rect 39021 46145 39067 46191
rect 39144 46145 39190 46191
rect 39267 46145 39313 46191
rect 44812 46232 44858 46278
rect 44925 46232 44971 46278
rect 45038 46232 45084 46278
rect 45151 46232 45197 46278
rect 45264 46232 45310 46278
rect 51802 46680 53776 46726
rect 51802 46456 53776 46502
rect 48778 46145 48824 46191
rect 48881 46145 48927 46191
rect 48984 46145 49030 46191
rect 49087 46145 49133 46191
rect 49190 46145 49236 46191
rect 49293 46145 49339 46191
rect 49396 46145 49442 46191
rect 49499 46145 49545 46191
rect 49602 46145 49852 46191
rect 51802 46232 53776 46278
rect 29317 46004 29363 46050
rect 29478 46004 29524 46050
rect 29638 46004 29684 46050
rect 29798 46004 29844 46050
rect 29959 46004 30005 46050
rect 30121 46004 30167 46050
rect 30284 46004 30330 46050
rect 54793 46004 54839 46050
rect 54956 46004 55002 46050
rect 55118 46004 55164 46050
rect 55279 46004 55325 46050
rect 55439 46004 55485 46050
rect 55599 46004 55645 46050
rect 55760 46004 55806 46050
rect 31349 45776 33323 45822
rect 35273 45863 35523 45909
rect 35580 45863 35626 45909
rect 35683 45863 35729 45909
rect 35786 45863 35832 45909
rect 35889 45863 35935 45909
rect 35992 45863 36038 45909
rect 36095 45863 36141 45909
rect 36198 45863 36244 45909
rect 36301 45863 36347 45909
rect 36854 45863 36900 45909
rect 36971 45863 37017 45909
rect 37088 45863 37134 45909
rect 37206 45863 37252 45909
rect 37324 45863 37370 45909
rect 37442 45863 37488 45909
rect 39021 45863 39067 45909
rect 39144 45863 39190 45909
rect 39267 45863 39313 45909
rect 31349 45552 33323 45598
rect 31349 45328 33323 45374
rect 29317 45104 29363 45150
rect 29478 45104 29524 45150
rect 29638 45104 29684 45150
rect 29798 45104 29844 45150
rect 29959 45104 30005 45150
rect 30121 45104 30167 45150
rect 30284 45104 30330 45150
rect 35273 45639 35523 45685
rect 35580 45639 35626 45685
rect 35683 45639 35729 45685
rect 35786 45639 35832 45685
rect 35889 45639 35935 45685
rect 35992 45639 36038 45685
rect 36095 45639 36141 45685
rect 36198 45639 36244 45685
rect 36301 45639 36347 45685
rect 36854 45639 36900 45685
rect 36971 45639 37017 45685
rect 37088 45639 37134 45685
rect 37206 45639 37252 45685
rect 37324 45639 37370 45685
rect 37442 45639 37488 45685
rect 48778 45863 48824 45909
rect 48881 45863 48927 45909
rect 48984 45863 49030 45909
rect 49087 45863 49133 45909
rect 49190 45863 49236 45909
rect 49293 45863 49339 45909
rect 49396 45863 49442 45909
rect 49499 45863 49545 45909
rect 49602 45863 49852 45909
rect 44812 45776 44858 45822
rect 44925 45776 44971 45822
rect 45038 45776 45084 45822
rect 45151 45776 45197 45822
rect 45264 45776 45310 45822
rect 39021 45639 39067 45685
rect 39144 45639 39190 45685
rect 39267 45639 39313 45685
rect 44812 45552 44858 45598
rect 44925 45552 44971 45598
rect 45038 45552 45084 45598
rect 45151 45552 45197 45598
rect 45264 45552 45310 45598
rect 48778 45639 48824 45685
rect 48881 45639 48927 45685
rect 48984 45639 49030 45685
rect 49087 45639 49133 45685
rect 49190 45639 49236 45685
rect 49293 45639 49339 45685
rect 49396 45639 49442 45685
rect 49499 45639 49545 45685
rect 49602 45639 49852 45685
rect 51802 45776 53776 45822
rect 35273 45415 35523 45461
rect 35580 45415 35626 45461
rect 35683 45415 35729 45461
rect 35786 45415 35832 45461
rect 35889 45415 35935 45461
rect 35992 45415 36038 45461
rect 36095 45415 36141 45461
rect 36198 45415 36244 45461
rect 36301 45415 36347 45461
rect 36854 45415 36900 45461
rect 36971 45415 37017 45461
rect 37088 45415 37134 45461
rect 37206 45415 37252 45461
rect 37324 45415 37370 45461
rect 37442 45415 37488 45461
rect 48778 45415 48824 45461
rect 48881 45415 48927 45461
rect 48984 45415 49030 45461
rect 49087 45415 49133 45461
rect 49190 45415 49236 45461
rect 49293 45415 49339 45461
rect 49396 45415 49442 45461
rect 49499 45415 49545 45461
rect 49602 45415 49852 45461
rect 44812 45328 44858 45374
rect 44925 45328 44971 45374
rect 45038 45328 45084 45374
rect 45151 45328 45197 45374
rect 45264 45328 45310 45374
rect 31349 45104 33323 45150
rect 31349 44880 33323 44926
rect 31349 44656 33323 44702
rect 51802 45552 53776 45598
rect 51802 45328 53776 45374
rect 44812 45104 44858 45150
rect 44925 45104 44971 45150
rect 45038 45104 45084 45150
rect 45151 45104 45197 45150
rect 45264 45104 45310 45150
rect 51802 45104 53776 45150
rect 35273 44793 35523 44839
rect 35580 44793 35626 44839
rect 35683 44793 35729 44839
rect 35786 44793 35832 44839
rect 35889 44793 35935 44839
rect 35992 44793 36038 44839
rect 36095 44793 36141 44839
rect 36198 44793 36244 44839
rect 36301 44793 36347 44839
rect 36854 44793 36900 44839
rect 36971 44793 37017 44839
rect 37088 44793 37134 44839
rect 37206 44793 37252 44839
rect 37324 44793 37370 44839
rect 37442 44793 37488 44839
rect 44812 44880 44858 44926
rect 44925 44880 44971 44926
rect 45038 44880 45084 44926
rect 45151 44880 45197 44926
rect 45264 44880 45310 44926
rect 54793 45104 54839 45150
rect 54956 45104 55002 45150
rect 55118 45104 55164 45150
rect 55279 45104 55325 45150
rect 55439 45104 55485 45150
rect 55599 45104 55645 45150
rect 55760 45104 55806 45150
rect 31349 44432 33323 44478
rect 35273 44569 35523 44615
rect 35580 44569 35626 44615
rect 35683 44569 35729 44615
rect 35786 44569 35832 44615
rect 35889 44569 35935 44615
rect 35992 44569 36038 44615
rect 36095 44569 36141 44615
rect 36198 44569 36244 44615
rect 36301 44569 36347 44615
rect 48778 44793 48824 44839
rect 48881 44793 48927 44839
rect 48984 44793 49030 44839
rect 49087 44793 49133 44839
rect 49190 44793 49236 44839
rect 49293 44793 49339 44839
rect 49396 44793 49442 44839
rect 49499 44793 49545 44839
rect 49602 44793 49852 44839
rect 36854 44569 36900 44615
rect 36971 44569 37017 44615
rect 37088 44569 37134 44615
rect 37206 44569 37252 44615
rect 37324 44569 37370 44615
rect 37442 44569 37488 44615
rect 39021 44569 39067 44615
rect 39144 44569 39190 44615
rect 39267 44569 39313 44615
rect 44812 44656 44858 44702
rect 44925 44656 44971 44702
rect 45038 44656 45084 44702
rect 45151 44656 45197 44702
rect 45264 44656 45310 44702
rect 48778 44569 48824 44615
rect 48881 44569 48927 44615
rect 48984 44569 49030 44615
rect 49087 44569 49133 44615
rect 49190 44569 49236 44615
rect 49293 44569 49339 44615
rect 49396 44569 49442 44615
rect 49499 44569 49545 44615
rect 49602 44569 49852 44615
rect 35273 44345 35523 44391
rect 35580 44345 35626 44391
rect 35683 44345 35729 44391
rect 35786 44345 35832 44391
rect 35889 44345 35935 44391
rect 35992 44345 36038 44391
rect 36095 44345 36141 44391
rect 36198 44345 36244 44391
rect 36301 44345 36347 44391
rect 36854 44345 36900 44391
rect 36971 44345 37017 44391
rect 37088 44345 37134 44391
rect 37206 44345 37252 44391
rect 37324 44345 37370 44391
rect 37442 44345 37488 44391
rect 39021 44345 39067 44391
rect 39144 44345 39190 44391
rect 39267 44345 39313 44391
rect 44812 44432 44858 44478
rect 44925 44432 44971 44478
rect 45038 44432 45084 44478
rect 45151 44432 45197 44478
rect 45264 44432 45310 44478
rect 51802 44880 53776 44926
rect 51802 44656 53776 44702
rect 48778 44345 48824 44391
rect 48881 44345 48927 44391
rect 48984 44345 49030 44391
rect 49087 44345 49133 44391
rect 49190 44345 49236 44391
rect 49293 44345 49339 44391
rect 49396 44345 49442 44391
rect 49499 44345 49545 44391
rect 49602 44345 49852 44391
rect 51802 44432 53776 44478
rect 29317 44204 29363 44250
rect 29478 44204 29524 44250
rect 29638 44204 29684 44250
rect 29798 44204 29844 44250
rect 29959 44204 30005 44250
rect 30121 44204 30167 44250
rect 30284 44204 30330 44250
rect 54793 44204 54839 44250
rect 54956 44204 55002 44250
rect 55118 44204 55164 44250
rect 55279 44204 55325 44250
rect 55439 44204 55485 44250
rect 55599 44204 55645 44250
rect 55760 44204 55806 44250
rect 31349 43976 33323 44022
rect 35273 44063 35523 44109
rect 35580 44063 35626 44109
rect 35683 44063 35729 44109
rect 35786 44063 35832 44109
rect 35889 44063 35935 44109
rect 35992 44063 36038 44109
rect 36095 44063 36141 44109
rect 36198 44063 36244 44109
rect 36301 44063 36347 44109
rect 36854 44063 36900 44109
rect 36971 44063 37017 44109
rect 37088 44063 37134 44109
rect 37206 44063 37252 44109
rect 37324 44063 37370 44109
rect 37442 44063 37488 44109
rect 39021 44063 39067 44109
rect 39144 44063 39190 44109
rect 39267 44063 39313 44109
rect 31349 43752 33323 43798
rect 31349 43528 33323 43574
rect 29317 43304 29363 43350
rect 29478 43304 29524 43350
rect 29638 43304 29684 43350
rect 29798 43304 29844 43350
rect 29959 43304 30005 43350
rect 30121 43304 30167 43350
rect 30284 43304 30330 43350
rect 35273 43839 35523 43885
rect 35580 43839 35626 43885
rect 35683 43839 35729 43885
rect 35786 43839 35832 43885
rect 35889 43839 35935 43885
rect 35992 43839 36038 43885
rect 36095 43839 36141 43885
rect 36198 43839 36244 43885
rect 36301 43839 36347 43885
rect 36854 43839 36900 43885
rect 36971 43839 37017 43885
rect 37088 43839 37134 43885
rect 37206 43839 37252 43885
rect 37324 43839 37370 43885
rect 37442 43839 37488 43885
rect 48778 44063 48824 44109
rect 48881 44063 48927 44109
rect 48984 44063 49030 44109
rect 49087 44063 49133 44109
rect 49190 44063 49236 44109
rect 49293 44063 49339 44109
rect 49396 44063 49442 44109
rect 49499 44063 49545 44109
rect 49602 44063 49852 44109
rect 44812 43976 44858 44022
rect 44925 43976 44971 44022
rect 45038 43976 45084 44022
rect 45151 43976 45197 44022
rect 45264 43976 45310 44022
rect 39021 43839 39067 43885
rect 39144 43839 39190 43885
rect 39267 43839 39313 43885
rect 44812 43752 44858 43798
rect 44925 43752 44971 43798
rect 45038 43752 45084 43798
rect 45151 43752 45197 43798
rect 45264 43752 45310 43798
rect 48778 43839 48824 43885
rect 48881 43839 48927 43885
rect 48984 43839 49030 43885
rect 49087 43839 49133 43885
rect 49190 43839 49236 43885
rect 49293 43839 49339 43885
rect 49396 43839 49442 43885
rect 49499 43839 49545 43885
rect 49602 43839 49852 43885
rect 51802 43976 53776 44022
rect 35273 43615 35523 43661
rect 35580 43615 35626 43661
rect 35683 43615 35729 43661
rect 35786 43615 35832 43661
rect 35889 43615 35935 43661
rect 35992 43615 36038 43661
rect 36095 43615 36141 43661
rect 36198 43615 36244 43661
rect 36301 43615 36347 43661
rect 36854 43615 36900 43661
rect 36971 43615 37017 43661
rect 37088 43615 37134 43661
rect 37206 43615 37252 43661
rect 37324 43615 37370 43661
rect 37442 43615 37488 43661
rect 48778 43615 48824 43661
rect 48881 43615 48927 43661
rect 48984 43615 49030 43661
rect 49087 43615 49133 43661
rect 49190 43615 49236 43661
rect 49293 43615 49339 43661
rect 49396 43615 49442 43661
rect 49499 43615 49545 43661
rect 49602 43615 49852 43661
rect 44812 43528 44858 43574
rect 44925 43528 44971 43574
rect 45038 43528 45084 43574
rect 45151 43528 45197 43574
rect 45264 43528 45310 43574
rect 31349 43304 33323 43350
rect 31349 43080 33323 43126
rect 31349 42856 33323 42902
rect 51802 43752 53776 43798
rect 51802 43528 53776 43574
rect 44812 43304 44858 43350
rect 44925 43304 44971 43350
rect 45038 43304 45084 43350
rect 45151 43304 45197 43350
rect 45264 43304 45310 43350
rect 51802 43304 53776 43350
rect 35273 42993 35523 43039
rect 35580 42993 35626 43039
rect 35683 42993 35729 43039
rect 35786 42993 35832 43039
rect 35889 42993 35935 43039
rect 35992 42993 36038 43039
rect 36095 42993 36141 43039
rect 36198 42993 36244 43039
rect 36301 42993 36347 43039
rect 36854 42993 36900 43039
rect 36971 42993 37017 43039
rect 37088 42993 37134 43039
rect 37206 42993 37252 43039
rect 37324 42993 37370 43039
rect 37442 42993 37488 43039
rect 44812 43080 44858 43126
rect 44925 43080 44971 43126
rect 45038 43080 45084 43126
rect 45151 43080 45197 43126
rect 45264 43080 45310 43126
rect 54793 43304 54839 43350
rect 54956 43304 55002 43350
rect 55118 43304 55164 43350
rect 55279 43304 55325 43350
rect 55439 43304 55485 43350
rect 55599 43304 55645 43350
rect 55760 43304 55806 43350
rect 31349 42632 33323 42678
rect 35273 42769 35523 42815
rect 35580 42769 35626 42815
rect 35683 42769 35729 42815
rect 35786 42769 35832 42815
rect 35889 42769 35935 42815
rect 35992 42769 36038 42815
rect 36095 42769 36141 42815
rect 36198 42769 36244 42815
rect 36301 42769 36347 42815
rect 48778 42993 48824 43039
rect 48881 42993 48927 43039
rect 48984 42993 49030 43039
rect 49087 42993 49133 43039
rect 49190 42993 49236 43039
rect 49293 42993 49339 43039
rect 49396 42993 49442 43039
rect 49499 42993 49545 43039
rect 49602 42993 49852 43039
rect 36854 42769 36900 42815
rect 36971 42769 37017 42815
rect 37088 42769 37134 42815
rect 37206 42769 37252 42815
rect 37324 42769 37370 42815
rect 37442 42769 37488 42815
rect 39021 42769 39067 42815
rect 39144 42769 39190 42815
rect 39267 42769 39313 42815
rect 44812 42856 44858 42902
rect 44925 42856 44971 42902
rect 45038 42856 45084 42902
rect 45151 42856 45197 42902
rect 45264 42856 45310 42902
rect 48778 42769 48824 42815
rect 48881 42769 48927 42815
rect 48984 42769 49030 42815
rect 49087 42769 49133 42815
rect 49190 42769 49236 42815
rect 49293 42769 49339 42815
rect 49396 42769 49442 42815
rect 49499 42769 49545 42815
rect 49602 42769 49852 42815
rect 35273 42545 35523 42591
rect 35580 42545 35626 42591
rect 35683 42545 35729 42591
rect 35786 42545 35832 42591
rect 35889 42545 35935 42591
rect 35992 42545 36038 42591
rect 36095 42545 36141 42591
rect 36198 42545 36244 42591
rect 36301 42545 36347 42591
rect 36854 42545 36900 42591
rect 36971 42545 37017 42591
rect 37088 42545 37134 42591
rect 37206 42545 37252 42591
rect 37324 42545 37370 42591
rect 37442 42545 37488 42591
rect 39021 42545 39067 42591
rect 39144 42545 39190 42591
rect 39267 42545 39313 42591
rect 44812 42632 44858 42678
rect 44925 42632 44971 42678
rect 45038 42632 45084 42678
rect 45151 42632 45197 42678
rect 45264 42632 45310 42678
rect 51802 43080 53776 43126
rect 51802 42856 53776 42902
rect 48778 42545 48824 42591
rect 48881 42545 48927 42591
rect 48984 42545 49030 42591
rect 49087 42545 49133 42591
rect 49190 42545 49236 42591
rect 49293 42545 49339 42591
rect 49396 42545 49442 42591
rect 49499 42545 49545 42591
rect 49602 42545 49852 42591
rect 51802 42632 53776 42678
rect 29317 42404 29363 42450
rect 29478 42404 29524 42450
rect 29638 42404 29684 42450
rect 29798 42404 29844 42450
rect 29959 42404 30005 42450
rect 30121 42404 30167 42450
rect 30284 42404 30330 42450
rect 54793 42404 54839 42450
rect 54956 42404 55002 42450
rect 55118 42404 55164 42450
rect 55279 42404 55325 42450
rect 55439 42404 55485 42450
rect 55599 42404 55645 42450
rect 55760 42404 55806 42450
rect 31349 42176 33323 42222
rect 35273 42263 35523 42309
rect 35580 42263 35626 42309
rect 35683 42263 35729 42309
rect 35786 42263 35832 42309
rect 35889 42263 35935 42309
rect 35992 42263 36038 42309
rect 36095 42263 36141 42309
rect 36198 42263 36244 42309
rect 36301 42263 36347 42309
rect 36854 42263 36900 42309
rect 36971 42263 37017 42309
rect 37088 42263 37134 42309
rect 37206 42263 37252 42309
rect 37324 42263 37370 42309
rect 37442 42263 37488 42309
rect 39021 42263 39067 42309
rect 39144 42263 39190 42309
rect 39267 42263 39313 42309
rect 31349 41952 33323 41998
rect 31349 41728 33323 41774
rect 29317 41504 29363 41550
rect 29478 41504 29524 41550
rect 29638 41504 29684 41550
rect 29798 41504 29844 41550
rect 29959 41504 30005 41550
rect 30121 41504 30167 41550
rect 30284 41504 30330 41550
rect 35273 42039 35523 42085
rect 35580 42039 35626 42085
rect 35683 42039 35729 42085
rect 35786 42039 35832 42085
rect 35889 42039 35935 42085
rect 35992 42039 36038 42085
rect 36095 42039 36141 42085
rect 36198 42039 36244 42085
rect 36301 42039 36347 42085
rect 36854 42039 36900 42085
rect 36971 42039 37017 42085
rect 37088 42039 37134 42085
rect 37206 42039 37252 42085
rect 37324 42039 37370 42085
rect 37442 42039 37488 42085
rect 48778 42263 48824 42309
rect 48881 42263 48927 42309
rect 48984 42263 49030 42309
rect 49087 42263 49133 42309
rect 49190 42263 49236 42309
rect 49293 42263 49339 42309
rect 49396 42263 49442 42309
rect 49499 42263 49545 42309
rect 49602 42263 49852 42309
rect 44812 42176 44858 42222
rect 44925 42176 44971 42222
rect 45038 42176 45084 42222
rect 45151 42176 45197 42222
rect 45264 42176 45310 42222
rect 39021 42039 39067 42085
rect 39144 42039 39190 42085
rect 39267 42039 39313 42085
rect 44812 41952 44858 41998
rect 44925 41952 44971 41998
rect 45038 41952 45084 41998
rect 45151 41952 45197 41998
rect 45264 41952 45310 41998
rect 48778 42039 48824 42085
rect 48881 42039 48927 42085
rect 48984 42039 49030 42085
rect 49087 42039 49133 42085
rect 49190 42039 49236 42085
rect 49293 42039 49339 42085
rect 49396 42039 49442 42085
rect 49499 42039 49545 42085
rect 49602 42039 49852 42085
rect 51802 42176 53776 42222
rect 35273 41815 35523 41861
rect 35580 41815 35626 41861
rect 35683 41815 35729 41861
rect 35786 41815 35832 41861
rect 35889 41815 35935 41861
rect 35992 41815 36038 41861
rect 36095 41815 36141 41861
rect 36198 41815 36244 41861
rect 36301 41815 36347 41861
rect 36854 41815 36900 41861
rect 36971 41815 37017 41861
rect 37088 41815 37134 41861
rect 37206 41815 37252 41861
rect 37324 41815 37370 41861
rect 37442 41815 37488 41861
rect 48778 41815 48824 41861
rect 48881 41815 48927 41861
rect 48984 41815 49030 41861
rect 49087 41815 49133 41861
rect 49190 41815 49236 41861
rect 49293 41815 49339 41861
rect 49396 41815 49442 41861
rect 49499 41815 49545 41861
rect 49602 41815 49852 41861
rect 44812 41728 44858 41774
rect 44925 41728 44971 41774
rect 45038 41728 45084 41774
rect 45151 41728 45197 41774
rect 45264 41728 45310 41774
rect 31349 41504 33323 41550
rect 31349 41280 33323 41326
rect 31349 41056 33323 41102
rect 51802 41952 53776 41998
rect 51802 41728 53776 41774
rect 44812 41504 44858 41550
rect 44925 41504 44971 41550
rect 45038 41504 45084 41550
rect 45151 41504 45197 41550
rect 45264 41504 45310 41550
rect 51802 41504 53776 41550
rect 35273 41193 35523 41239
rect 35580 41193 35626 41239
rect 35683 41193 35729 41239
rect 35786 41193 35832 41239
rect 35889 41193 35935 41239
rect 35992 41193 36038 41239
rect 36095 41193 36141 41239
rect 36198 41193 36244 41239
rect 36301 41193 36347 41239
rect 36854 41193 36900 41239
rect 36971 41193 37017 41239
rect 37088 41193 37134 41239
rect 37206 41193 37252 41239
rect 37324 41193 37370 41239
rect 37442 41193 37488 41239
rect 44812 41280 44858 41326
rect 44925 41280 44971 41326
rect 45038 41280 45084 41326
rect 45151 41280 45197 41326
rect 45264 41280 45310 41326
rect 54793 41504 54839 41550
rect 54956 41504 55002 41550
rect 55118 41504 55164 41550
rect 55279 41504 55325 41550
rect 55439 41504 55485 41550
rect 55599 41504 55645 41550
rect 55760 41504 55806 41550
rect 31349 40832 33323 40878
rect 35273 40969 35523 41015
rect 35580 40969 35626 41015
rect 35683 40969 35729 41015
rect 35786 40969 35832 41015
rect 35889 40969 35935 41015
rect 35992 40969 36038 41015
rect 36095 40969 36141 41015
rect 36198 40969 36244 41015
rect 36301 40969 36347 41015
rect 48778 41193 48824 41239
rect 48881 41193 48927 41239
rect 48984 41193 49030 41239
rect 49087 41193 49133 41239
rect 49190 41193 49236 41239
rect 49293 41193 49339 41239
rect 49396 41193 49442 41239
rect 49499 41193 49545 41239
rect 49602 41193 49852 41239
rect 36854 40969 36900 41015
rect 36971 40969 37017 41015
rect 37088 40969 37134 41015
rect 37206 40969 37252 41015
rect 37324 40969 37370 41015
rect 37442 40969 37488 41015
rect 39021 40969 39067 41015
rect 39144 40969 39190 41015
rect 39267 40969 39313 41015
rect 44812 41056 44858 41102
rect 44925 41056 44971 41102
rect 45038 41056 45084 41102
rect 45151 41056 45197 41102
rect 45264 41056 45310 41102
rect 48778 40969 48824 41015
rect 48881 40969 48927 41015
rect 48984 40969 49030 41015
rect 49087 40969 49133 41015
rect 49190 40969 49236 41015
rect 49293 40969 49339 41015
rect 49396 40969 49442 41015
rect 49499 40969 49545 41015
rect 49602 40969 49852 41015
rect 35273 40745 35523 40791
rect 35580 40745 35626 40791
rect 35683 40745 35729 40791
rect 35786 40745 35832 40791
rect 35889 40745 35935 40791
rect 35992 40745 36038 40791
rect 36095 40745 36141 40791
rect 36198 40745 36244 40791
rect 36301 40745 36347 40791
rect 36854 40745 36900 40791
rect 36971 40745 37017 40791
rect 37088 40745 37134 40791
rect 37206 40745 37252 40791
rect 37324 40745 37370 40791
rect 37442 40745 37488 40791
rect 39021 40745 39067 40791
rect 39144 40745 39190 40791
rect 39267 40745 39313 40791
rect 44812 40832 44858 40878
rect 44925 40832 44971 40878
rect 45038 40832 45084 40878
rect 45151 40832 45197 40878
rect 45264 40832 45310 40878
rect 51802 41280 53776 41326
rect 51802 41056 53776 41102
rect 48778 40745 48824 40791
rect 48881 40745 48927 40791
rect 48984 40745 49030 40791
rect 49087 40745 49133 40791
rect 49190 40745 49236 40791
rect 49293 40745 49339 40791
rect 49396 40745 49442 40791
rect 49499 40745 49545 40791
rect 49602 40745 49852 40791
rect 51802 40832 53776 40878
rect 29317 40604 29363 40650
rect 29478 40604 29524 40650
rect 29638 40604 29684 40650
rect 29798 40604 29844 40650
rect 29959 40604 30005 40650
rect 30121 40604 30167 40650
rect 30284 40604 30330 40650
rect 54793 40604 54839 40650
rect 54956 40604 55002 40650
rect 55118 40604 55164 40650
rect 55279 40604 55325 40650
rect 55439 40604 55485 40650
rect 55599 40604 55645 40650
rect 55760 40604 55806 40650
rect 31349 40376 33323 40422
rect 35273 40463 35523 40509
rect 35580 40463 35626 40509
rect 35683 40463 35729 40509
rect 35786 40463 35832 40509
rect 35889 40463 35935 40509
rect 35992 40463 36038 40509
rect 36095 40463 36141 40509
rect 36198 40463 36244 40509
rect 36301 40463 36347 40509
rect 36854 40463 36900 40509
rect 36971 40463 37017 40509
rect 37088 40463 37134 40509
rect 37206 40463 37252 40509
rect 37324 40463 37370 40509
rect 37442 40463 37488 40509
rect 39021 40463 39067 40509
rect 39144 40463 39190 40509
rect 39267 40463 39313 40509
rect 31349 40152 33323 40198
rect 31349 39928 33323 39974
rect 29317 39704 29363 39750
rect 29478 39704 29524 39750
rect 29638 39704 29684 39750
rect 29798 39704 29844 39750
rect 29959 39704 30005 39750
rect 30121 39704 30167 39750
rect 30284 39704 30330 39750
rect 35273 40239 35523 40285
rect 35580 40239 35626 40285
rect 35683 40239 35729 40285
rect 35786 40239 35832 40285
rect 35889 40239 35935 40285
rect 35992 40239 36038 40285
rect 36095 40239 36141 40285
rect 36198 40239 36244 40285
rect 36301 40239 36347 40285
rect 36854 40239 36900 40285
rect 36971 40239 37017 40285
rect 37088 40239 37134 40285
rect 37206 40239 37252 40285
rect 37324 40239 37370 40285
rect 37442 40239 37488 40285
rect 48778 40463 48824 40509
rect 48881 40463 48927 40509
rect 48984 40463 49030 40509
rect 49087 40463 49133 40509
rect 49190 40463 49236 40509
rect 49293 40463 49339 40509
rect 49396 40463 49442 40509
rect 49499 40463 49545 40509
rect 49602 40463 49852 40509
rect 44812 40376 44858 40422
rect 44925 40376 44971 40422
rect 45038 40376 45084 40422
rect 45151 40376 45197 40422
rect 45264 40376 45310 40422
rect 39021 40239 39067 40285
rect 39144 40239 39190 40285
rect 39267 40239 39313 40285
rect 44812 40152 44858 40198
rect 44925 40152 44971 40198
rect 45038 40152 45084 40198
rect 45151 40152 45197 40198
rect 45264 40152 45310 40198
rect 48778 40239 48824 40285
rect 48881 40239 48927 40285
rect 48984 40239 49030 40285
rect 49087 40239 49133 40285
rect 49190 40239 49236 40285
rect 49293 40239 49339 40285
rect 49396 40239 49442 40285
rect 49499 40239 49545 40285
rect 49602 40239 49852 40285
rect 51802 40376 53776 40422
rect 35273 40015 35523 40061
rect 35580 40015 35626 40061
rect 35683 40015 35729 40061
rect 35786 40015 35832 40061
rect 35889 40015 35935 40061
rect 35992 40015 36038 40061
rect 36095 40015 36141 40061
rect 36198 40015 36244 40061
rect 36301 40015 36347 40061
rect 36854 40015 36900 40061
rect 36971 40015 37017 40061
rect 37088 40015 37134 40061
rect 37206 40015 37252 40061
rect 37324 40015 37370 40061
rect 37442 40015 37488 40061
rect 48778 40015 48824 40061
rect 48881 40015 48927 40061
rect 48984 40015 49030 40061
rect 49087 40015 49133 40061
rect 49190 40015 49236 40061
rect 49293 40015 49339 40061
rect 49396 40015 49442 40061
rect 49499 40015 49545 40061
rect 49602 40015 49852 40061
rect 44812 39928 44858 39974
rect 44925 39928 44971 39974
rect 45038 39928 45084 39974
rect 45151 39928 45197 39974
rect 45264 39928 45310 39974
rect 31349 39704 33323 39750
rect 31349 39480 33323 39526
rect 31349 39256 33323 39302
rect 51802 40152 53776 40198
rect 51802 39928 53776 39974
rect 44812 39704 44858 39750
rect 44925 39704 44971 39750
rect 45038 39704 45084 39750
rect 45151 39704 45197 39750
rect 45264 39704 45310 39750
rect 51802 39704 53776 39750
rect 35273 39393 35523 39439
rect 35580 39393 35626 39439
rect 35683 39393 35729 39439
rect 35786 39393 35832 39439
rect 35889 39393 35935 39439
rect 35992 39393 36038 39439
rect 36095 39393 36141 39439
rect 36198 39393 36244 39439
rect 36301 39393 36347 39439
rect 36854 39393 36900 39439
rect 36971 39393 37017 39439
rect 37088 39393 37134 39439
rect 37206 39393 37252 39439
rect 37324 39393 37370 39439
rect 37442 39393 37488 39439
rect 44812 39480 44858 39526
rect 44925 39480 44971 39526
rect 45038 39480 45084 39526
rect 45151 39480 45197 39526
rect 45264 39480 45310 39526
rect 54793 39704 54839 39750
rect 54956 39704 55002 39750
rect 55118 39704 55164 39750
rect 55279 39704 55325 39750
rect 55439 39704 55485 39750
rect 55599 39704 55645 39750
rect 55760 39704 55806 39750
rect 31349 39032 33323 39078
rect 35273 39169 35523 39215
rect 35580 39169 35626 39215
rect 35683 39169 35729 39215
rect 35786 39169 35832 39215
rect 35889 39169 35935 39215
rect 35992 39169 36038 39215
rect 36095 39169 36141 39215
rect 36198 39169 36244 39215
rect 36301 39169 36347 39215
rect 48778 39393 48824 39439
rect 48881 39393 48927 39439
rect 48984 39393 49030 39439
rect 49087 39393 49133 39439
rect 49190 39393 49236 39439
rect 49293 39393 49339 39439
rect 49396 39393 49442 39439
rect 49499 39393 49545 39439
rect 49602 39393 49852 39439
rect 36854 39169 36900 39215
rect 36971 39169 37017 39215
rect 37088 39169 37134 39215
rect 37206 39169 37252 39215
rect 37324 39169 37370 39215
rect 37442 39169 37488 39215
rect 39021 39169 39067 39215
rect 39144 39169 39190 39215
rect 39267 39169 39313 39215
rect 44812 39256 44858 39302
rect 44925 39256 44971 39302
rect 45038 39256 45084 39302
rect 45151 39256 45197 39302
rect 45264 39256 45310 39302
rect 48778 39169 48824 39215
rect 48881 39169 48927 39215
rect 48984 39169 49030 39215
rect 49087 39169 49133 39215
rect 49190 39169 49236 39215
rect 49293 39169 49339 39215
rect 49396 39169 49442 39215
rect 49499 39169 49545 39215
rect 49602 39169 49852 39215
rect 35273 38945 35523 38991
rect 35580 38945 35626 38991
rect 35683 38945 35729 38991
rect 35786 38945 35832 38991
rect 35889 38945 35935 38991
rect 35992 38945 36038 38991
rect 36095 38945 36141 38991
rect 36198 38945 36244 38991
rect 36301 38945 36347 38991
rect 36854 38945 36900 38991
rect 36971 38945 37017 38991
rect 37088 38945 37134 38991
rect 37206 38945 37252 38991
rect 37324 38945 37370 38991
rect 37442 38945 37488 38991
rect 39021 38945 39067 38991
rect 39144 38945 39190 38991
rect 39267 38945 39313 38991
rect 44812 39032 44858 39078
rect 44925 39032 44971 39078
rect 45038 39032 45084 39078
rect 45151 39032 45197 39078
rect 45264 39032 45310 39078
rect 51802 39480 53776 39526
rect 51802 39256 53776 39302
rect 48778 38945 48824 38991
rect 48881 38945 48927 38991
rect 48984 38945 49030 38991
rect 49087 38945 49133 38991
rect 49190 38945 49236 38991
rect 49293 38945 49339 38991
rect 49396 38945 49442 38991
rect 49499 38945 49545 38991
rect 49602 38945 49852 38991
rect 51802 39032 53776 39078
rect 29317 38804 29363 38850
rect 29478 38804 29524 38850
rect 29638 38804 29684 38850
rect 29798 38804 29844 38850
rect 29959 38804 30005 38850
rect 30121 38804 30167 38850
rect 30284 38804 30330 38850
rect 54793 38804 54839 38850
rect 54956 38804 55002 38850
rect 55118 38804 55164 38850
rect 55279 38804 55325 38850
rect 55439 38804 55485 38850
rect 55599 38804 55645 38850
rect 55760 38804 55806 38850
rect 31349 38576 33323 38622
rect 35273 38663 35523 38709
rect 35580 38663 35626 38709
rect 35683 38663 35729 38709
rect 35786 38663 35832 38709
rect 35889 38663 35935 38709
rect 35992 38663 36038 38709
rect 36095 38663 36141 38709
rect 36198 38663 36244 38709
rect 36301 38663 36347 38709
rect 36854 38663 36900 38709
rect 36971 38663 37017 38709
rect 37088 38663 37134 38709
rect 37206 38663 37252 38709
rect 37324 38663 37370 38709
rect 37442 38663 37488 38709
rect 39021 38663 39067 38709
rect 39144 38663 39190 38709
rect 39267 38663 39313 38709
rect 31349 38352 33323 38398
rect 31349 38128 33323 38174
rect 29317 37904 29363 37950
rect 29478 37904 29524 37950
rect 29638 37904 29684 37950
rect 29798 37904 29844 37950
rect 29959 37904 30005 37950
rect 30121 37904 30167 37950
rect 30284 37904 30330 37950
rect 35273 38439 35523 38485
rect 35580 38439 35626 38485
rect 35683 38439 35729 38485
rect 35786 38439 35832 38485
rect 35889 38439 35935 38485
rect 35992 38439 36038 38485
rect 36095 38439 36141 38485
rect 36198 38439 36244 38485
rect 36301 38439 36347 38485
rect 36854 38439 36900 38485
rect 36971 38439 37017 38485
rect 37088 38439 37134 38485
rect 37206 38439 37252 38485
rect 37324 38439 37370 38485
rect 37442 38439 37488 38485
rect 48778 38663 48824 38709
rect 48881 38663 48927 38709
rect 48984 38663 49030 38709
rect 49087 38663 49133 38709
rect 49190 38663 49236 38709
rect 49293 38663 49339 38709
rect 49396 38663 49442 38709
rect 49499 38663 49545 38709
rect 49602 38663 49852 38709
rect 44812 38576 44858 38622
rect 44925 38576 44971 38622
rect 45038 38576 45084 38622
rect 45151 38576 45197 38622
rect 45264 38576 45310 38622
rect 39021 38439 39067 38485
rect 39144 38439 39190 38485
rect 39267 38439 39313 38485
rect 44812 38352 44858 38398
rect 44925 38352 44971 38398
rect 45038 38352 45084 38398
rect 45151 38352 45197 38398
rect 45264 38352 45310 38398
rect 48778 38439 48824 38485
rect 48881 38439 48927 38485
rect 48984 38439 49030 38485
rect 49087 38439 49133 38485
rect 49190 38439 49236 38485
rect 49293 38439 49339 38485
rect 49396 38439 49442 38485
rect 49499 38439 49545 38485
rect 49602 38439 49852 38485
rect 51802 38576 53776 38622
rect 35273 38215 35523 38261
rect 35580 38215 35626 38261
rect 35683 38215 35729 38261
rect 35786 38215 35832 38261
rect 35889 38215 35935 38261
rect 35992 38215 36038 38261
rect 36095 38215 36141 38261
rect 36198 38215 36244 38261
rect 36301 38215 36347 38261
rect 36854 38215 36900 38261
rect 36971 38215 37017 38261
rect 37088 38215 37134 38261
rect 37206 38215 37252 38261
rect 37324 38215 37370 38261
rect 37442 38215 37488 38261
rect 48778 38215 48824 38261
rect 48881 38215 48927 38261
rect 48984 38215 49030 38261
rect 49087 38215 49133 38261
rect 49190 38215 49236 38261
rect 49293 38215 49339 38261
rect 49396 38215 49442 38261
rect 49499 38215 49545 38261
rect 49602 38215 49852 38261
rect 44812 38128 44858 38174
rect 44925 38128 44971 38174
rect 45038 38128 45084 38174
rect 45151 38128 45197 38174
rect 45264 38128 45310 38174
rect 31349 37904 33323 37950
rect 31349 37680 33323 37726
rect 31349 37456 33323 37502
rect 51802 38352 53776 38398
rect 51802 38128 53776 38174
rect 44812 37904 44858 37950
rect 44925 37904 44971 37950
rect 45038 37904 45084 37950
rect 45151 37904 45197 37950
rect 45264 37904 45310 37950
rect 51802 37904 53776 37950
rect 35273 37593 35523 37639
rect 35580 37593 35626 37639
rect 35683 37593 35729 37639
rect 35786 37593 35832 37639
rect 35889 37593 35935 37639
rect 35992 37593 36038 37639
rect 36095 37593 36141 37639
rect 36198 37593 36244 37639
rect 36301 37593 36347 37639
rect 36854 37593 36900 37639
rect 36971 37593 37017 37639
rect 37088 37593 37134 37639
rect 37206 37593 37252 37639
rect 37324 37593 37370 37639
rect 37442 37593 37488 37639
rect 44812 37680 44858 37726
rect 44925 37680 44971 37726
rect 45038 37680 45084 37726
rect 45151 37680 45197 37726
rect 45264 37680 45310 37726
rect 54793 37904 54839 37950
rect 54956 37904 55002 37950
rect 55118 37904 55164 37950
rect 55279 37904 55325 37950
rect 55439 37904 55485 37950
rect 55599 37904 55645 37950
rect 55760 37904 55806 37950
rect 31349 37232 33323 37278
rect 35273 37369 35523 37415
rect 35580 37369 35626 37415
rect 35683 37369 35729 37415
rect 35786 37369 35832 37415
rect 35889 37369 35935 37415
rect 35992 37369 36038 37415
rect 36095 37369 36141 37415
rect 36198 37369 36244 37415
rect 36301 37369 36347 37415
rect 48778 37593 48824 37639
rect 48881 37593 48927 37639
rect 48984 37593 49030 37639
rect 49087 37593 49133 37639
rect 49190 37593 49236 37639
rect 49293 37593 49339 37639
rect 49396 37593 49442 37639
rect 49499 37593 49545 37639
rect 49602 37593 49852 37639
rect 36854 37369 36900 37415
rect 36971 37369 37017 37415
rect 37088 37369 37134 37415
rect 37206 37369 37252 37415
rect 37324 37369 37370 37415
rect 37442 37369 37488 37415
rect 39021 37369 39067 37415
rect 39144 37369 39190 37415
rect 39267 37369 39313 37415
rect 44812 37456 44858 37502
rect 44925 37456 44971 37502
rect 45038 37456 45084 37502
rect 45151 37456 45197 37502
rect 45264 37456 45310 37502
rect 48778 37369 48824 37415
rect 48881 37369 48927 37415
rect 48984 37369 49030 37415
rect 49087 37369 49133 37415
rect 49190 37369 49236 37415
rect 49293 37369 49339 37415
rect 49396 37369 49442 37415
rect 49499 37369 49545 37415
rect 49602 37369 49852 37415
rect 35273 37145 35523 37191
rect 35580 37145 35626 37191
rect 35683 37145 35729 37191
rect 35786 37145 35832 37191
rect 35889 37145 35935 37191
rect 35992 37145 36038 37191
rect 36095 37145 36141 37191
rect 36198 37145 36244 37191
rect 36301 37145 36347 37191
rect 36854 37145 36900 37191
rect 36971 37145 37017 37191
rect 37088 37145 37134 37191
rect 37206 37145 37252 37191
rect 37324 37145 37370 37191
rect 37442 37145 37488 37191
rect 39021 37145 39067 37191
rect 39144 37145 39190 37191
rect 39267 37145 39313 37191
rect 44812 37232 44858 37278
rect 44925 37232 44971 37278
rect 45038 37232 45084 37278
rect 45151 37232 45197 37278
rect 45264 37232 45310 37278
rect 51802 37680 53776 37726
rect 51802 37456 53776 37502
rect 48778 37145 48824 37191
rect 48881 37145 48927 37191
rect 48984 37145 49030 37191
rect 49087 37145 49133 37191
rect 49190 37145 49236 37191
rect 49293 37145 49339 37191
rect 49396 37145 49442 37191
rect 49499 37145 49545 37191
rect 49602 37145 49852 37191
rect 51802 37232 53776 37278
rect 29317 37004 29363 37050
rect 29478 37004 29524 37050
rect 29638 37004 29684 37050
rect 29798 37004 29844 37050
rect 29959 37004 30005 37050
rect 30121 37004 30167 37050
rect 30284 37004 30330 37050
rect 54793 37004 54839 37050
rect 54956 37004 55002 37050
rect 55118 37004 55164 37050
rect 55279 37004 55325 37050
rect 55439 37004 55485 37050
rect 55599 37004 55645 37050
rect 55760 37004 55806 37050
rect 31349 36776 33323 36822
rect 35273 36863 35523 36909
rect 35580 36863 35626 36909
rect 35683 36863 35729 36909
rect 35786 36863 35832 36909
rect 35889 36863 35935 36909
rect 35992 36863 36038 36909
rect 36095 36863 36141 36909
rect 36198 36863 36244 36909
rect 36301 36863 36347 36909
rect 36854 36863 36900 36909
rect 36971 36863 37017 36909
rect 37088 36863 37134 36909
rect 37206 36863 37252 36909
rect 37324 36863 37370 36909
rect 37442 36863 37488 36909
rect 39021 36863 39067 36909
rect 39144 36863 39190 36909
rect 39267 36863 39313 36909
rect 31349 36552 33323 36598
rect 31349 36328 33323 36374
rect 29317 36104 29363 36150
rect 29478 36104 29524 36150
rect 29638 36104 29684 36150
rect 29798 36104 29844 36150
rect 29959 36104 30005 36150
rect 30121 36104 30167 36150
rect 30284 36104 30330 36150
rect 35273 36639 35523 36685
rect 35580 36639 35626 36685
rect 35683 36639 35729 36685
rect 35786 36639 35832 36685
rect 35889 36639 35935 36685
rect 35992 36639 36038 36685
rect 36095 36639 36141 36685
rect 36198 36639 36244 36685
rect 36301 36639 36347 36685
rect 36854 36639 36900 36685
rect 36971 36639 37017 36685
rect 37088 36639 37134 36685
rect 37206 36639 37252 36685
rect 37324 36639 37370 36685
rect 37442 36639 37488 36685
rect 48778 36863 48824 36909
rect 48881 36863 48927 36909
rect 48984 36863 49030 36909
rect 49087 36863 49133 36909
rect 49190 36863 49236 36909
rect 49293 36863 49339 36909
rect 49396 36863 49442 36909
rect 49499 36863 49545 36909
rect 49602 36863 49852 36909
rect 44812 36776 44858 36822
rect 44925 36776 44971 36822
rect 45038 36776 45084 36822
rect 45151 36776 45197 36822
rect 45264 36776 45310 36822
rect 39021 36639 39067 36685
rect 39144 36639 39190 36685
rect 39267 36639 39313 36685
rect 44812 36552 44858 36598
rect 44925 36552 44971 36598
rect 45038 36552 45084 36598
rect 45151 36552 45197 36598
rect 45264 36552 45310 36598
rect 48778 36639 48824 36685
rect 48881 36639 48927 36685
rect 48984 36639 49030 36685
rect 49087 36639 49133 36685
rect 49190 36639 49236 36685
rect 49293 36639 49339 36685
rect 49396 36639 49442 36685
rect 49499 36639 49545 36685
rect 49602 36639 49852 36685
rect 51802 36776 53776 36822
rect 35273 36415 35523 36461
rect 35580 36415 35626 36461
rect 35683 36415 35729 36461
rect 35786 36415 35832 36461
rect 35889 36415 35935 36461
rect 35992 36415 36038 36461
rect 36095 36415 36141 36461
rect 36198 36415 36244 36461
rect 36301 36415 36347 36461
rect 36854 36415 36900 36461
rect 36971 36415 37017 36461
rect 37088 36415 37134 36461
rect 37206 36415 37252 36461
rect 37324 36415 37370 36461
rect 37442 36415 37488 36461
rect 48778 36415 48824 36461
rect 48881 36415 48927 36461
rect 48984 36415 49030 36461
rect 49087 36415 49133 36461
rect 49190 36415 49236 36461
rect 49293 36415 49339 36461
rect 49396 36415 49442 36461
rect 49499 36415 49545 36461
rect 49602 36415 49852 36461
rect 44812 36328 44858 36374
rect 44925 36328 44971 36374
rect 45038 36328 45084 36374
rect 45151 36328 45197 36374
rect 45264 36328 45310 36374
rect 31349 36104 33323 36150
rect 51802 36552 53776 36598
rect 51802 36328 53776 36374
rect 44812 36104 44858 36150
rect 44925 36104 44971 36150
rect 45038 36104 45084 36150
rect 45151 36104 45197 36150
rect 45264 36104 45310 36150
rect 51802 36104 53776 36150
rect 54793 36104 54839 36150
rect 54956 36104 55002 36150
rect 55118 36104 55164 36150
rect 55279 36104 55325 36150
rect 55439 36104 55485 36150
rect 55599 36104 55645 36150
rect 55760 36104 55806 36150
<< mvpsubdiff >>
rect 28577 65722 28911 66109
rect 32989 65909 34884 65966
rect 32989 65863 33044 65909
rect 33090 65863 33202 65909
rect 33248 65863 33360 65909
rect 33406 65863 33518 65909
rect 33564 65863 33677 65909
rect 33723 65863 33835 65909
rect 33881 65863 33993 65909
rect 34039 65863 34151 65909
rect 34197 65863 34309 65909
rect 34355 65863 34467 65909
rect 34513 65863 34625 65909
rect 34671 65863 34783 65909
rect 34829 65863 34884 65909
rect 32989 65806 34884 65863
rect 40062 65909 41957 65966
rect 40062 65863 40117 65909
rect 40163 65863 40275 65909
rect 40321 65863 40433 65909
rect 40479 65863 40591 65909
rect 40637 65863 40750 65909
rect 40796 65863 40908 65909
rect 40954 65863 41066 65909
rect 41112 65863 41224 65909
rect 41270 65863 41382 65909
rect 41428 65863 41540 65909
rect 41586 65863 41698 65909
rect 41744 65863 41856 65909
rect 41902 65863 41957 65909
rect 28577 65676 28810 65722
rect 28856 65676 28911 65722
rect 28577 65558 28911 65676
rect 28577 65512 28810 65558
rect 28856 65512 28911 65558
rect 28577 65395 28911 65512
rect 28577 65349 28810 65395
rect 28856 65349 28911 65395
rect 28577 65232 28911 65349
rect 28577 65186 28810 65232
rect 28856 65186 28911 65232
rect 28577 65068 28911 65186
rect 28577 65022 28810 65068
rect 28856 65022 28911 65068
rect 28577 64866 28911 65022
rect 40062 65806 41957 65863
rect 44459 65909 44931 65966
rect 44459 65863 44514 65909
rect 44560 65863 44672 65909
rect 44718 65863 44830 65909
rect 44876 65863 44931 65909
rect 44459 65806 44931 65863
rect 50074 65909 51969 65966
rect 50074 65863 50129 65909
rect 50175 65863 50287 65909
rect 50333 65863 50445 65909
rect 50491 65863 50603 65909
rect 50649 65863 50762 65909
rect 50808 65863 50920 65909
rect 50966 65863 51078 65909
rect 51124 65863 51236 65909
rect 51282 65863 51394 65909
rect 51440 65863 51552 65909
rect 51598 65863 51710 65909
rect 51756 65863 51868 65909
rect 51914 65863 51969 65909
rect 50074 65806 51969 65863
rect 28577 64820 28810 64866
rect 28856 64820 28911 64866
rect 28577 64703 28911 64820
rect 28577 64657 28810 64703
rect 28856 64657 28911 64703
rect 28577 64540 28911 64657
rect 28577 64494 28810 64540
rect 28856 64494 28911 64540
rect 28577 64377 28911 64494
rect 28577 64331 28810 64377
rect 28856 64331 28911 64377
rect 28577 64213 28911 64331
rect 28577 64167 28810 64213
rect 28856 64167 28911 64213
rect 28577 64050 28911 64167
rect 37938 64950 38492 64969
rect 37938 64904 37957 64950
rect 38473 64904 38492 64950
rect 37938 64885 38492 64904
rect 40779 64950 42995 65010
rect 40779 64904 40836 64950
rect 40882 64904 40994 64950
rect 41040 64904 41152 64950
rect 41198 64904 41310 64950
rect 41356 64904 41469 64950
rect 41515 64904 41627 64950
rect 41673 64904 41785 64950
rect 41831 64904 41943 64950
rect 41989 64904 42101 64950
rect 42147 64904 42259 64950
rect 42305 64904 42418 64950
rect 42464 64904 42576 64950
rect 42622 64904 42734 64950
rect 42780 64904 42892 64950
rect 42938 64904 42995 64950
rect 40779 64844 42995 64904
rect 56212 65722 56546 66109
rect 56212 65676 56267 65722
rect 56313 65676 56546 65722
rect 56212 65558 56546 65676
rect 56212 65512 56267 65558
rect 56313 65512 56546 65558
rect 56212 65395 56546 65512
rect 56212 65349 56267 65395
rect 56313 65349 56546 65395
rect 56212 65232 56546 65349
rect 56212 65186 56267 65232
rect 56313 65186 56546 65232
rect 56212 65068 56546 65186
rect 56212 65022 56267 65068
rect 56313 65022 56546 65068
rect 28577 64004 28810 64050
rect 28856 64004 28911 64050
rect 28577 63887 28911 64004
rect 28577 63841 28810 63887
rect 28856 63841 28911 63887
rect 28577 63723 28911 63841
rect 28577 63677 28810 63723
rect 28856 63677 28911 63723
rect 28577 63560 28911 63677
rect 28577 63514 28810 63560
rect 28856 63514 28911 63560
rect 28577 63397 28911 63514
rect 28577 63351 28810 63397
rect 28856 63351 28911 63397
rect 28577 63234 28911 63351
rect 28577 63188 28810 63234
rect 28856 63188 28911 63234
rect 28577 63066 28911 63188
rect 34861 64050 35017 64107
rect 34861 64004 34916 64050
rect 34962 64004 35017 64050
rect 34861 63947 35017 64004
rect 50103 64050 50263 64110
rect 50103 64004 50160 64050
rect 50206 64004 50263 64050
rect 50103 63944 50263 64004
rect 56212 64866 56546 65022
rect 56212 64820 56267 64866
rect 56313 64820 56546 64866
rect 56212 64703 56546 64820
rect 56212 64657 56267 64703
rect 56313 64657 56546 64703
rect 56212 64540 56546 64657
rect 56212 64494 56267 64540
rect 56313 64494 56546 64540
rect 56212 64377 56546 64494
rect 56212 64331 56267 64377
rect 56313 64331 56546 64377
rect 56212 64213 56546 64331
rect 56212 64167 56267 64213
rect 56313 64167 56546 64213
rect 56212 64050 56546 64167
rect 56212 64004 56267 64050
rect 56313 64004 56546 64050
rect 28577 63020 28810 63066
rect 28856 63020 28911 63066
rect 28577 62903 28911 63020
rect 28577 62857 28810 62903
rect 28856 62857 28911 62903
rect 28577 62740 28911 62857
rect 28577 62694 28810 62740
rect 28856 62694 28911 62740
rect 28577 62577 28911 62694
rect 28577 62531 28810 62577
rect 28856 62531 28911 62577
rect 28577 62413 28911 62531
rect 28577 62367 28810 62413
rect 28856 62367 28911 62413
rect 28577 62250 28911 62367
rect 37938 63150 38492 63169
rect 37938 63104 37957 63150
rect 38473 63104 38492 63150
rect 37938 63085 38492 63104
rect 40779 63150 42995 63210
rect 40779 63104 40836 63150
rect 40882 63104 40994 63150
rect 41040 63104 41152 63150
rect 41198 63104 41310 63150
rect 41356 63104 41469 63150
rect 41515 63104 41627 63150
rect 41673 63104 41785 63150
rect 41831 63104 41943 63150
rect 41989 63104 42101 63150
rect 42147 63104 42259 63150
rect 42305 63104 42418 63150
rect 42464 63104 42576 63150
rect 42622 63104 42734 63150
rect 42780 63104 42892 63150
rect 42938 63104 42995 63150
rect 40779 63044 42995 63104
rect 56212 63887 56546 64004
rect 56212 63841 56267 63887
rect 56313 63841 56546 63887
rect 56212 63723 56546 63841
rect 56212 63677 56267 63723
rect 56313 63677 56546 63723
rect 56212 63560 56546 63677
rect 56212 63514 56267 63560
rect 56313 63514 56546 63560
rect 56212 63397 56546 63514
rect 56212 63351 56267 63397
rect 56313 63351 56546 63397
rect 56212 63234 56546 63351
rect 56212 63188 56267 63234
rect 56313 63188 56546 63234
rect 28577 62204 28810 62250
rect 28856 62204 28911 62250
rect 28577 62087 28911 62204
rect 28577 62041 28810 62087
rect 28856 62041 28911 62087
rect 28577 61923 28911 62041
rect 28577 61877 28810 61923
rect 28856 61877 28911 61923
rect 28577 61760 28911 61877
rect 28577 61714 28810 61760
rect 28856 61714 28911 61760
rect 28577 61597 28911 61714
rect 28577 61551 28810 61597
rect 28856 61551 28911 61597
rect 28577 61434 28911 61551
rect 28577 61388 28810 61434
rect 28856 61388 28911 61434
rect 28577 61266 28911 61388
rect 34861 62250 35017 62307
rect 34861 62204 34916 62250
rect 34962 62204 35017 62250
rect 34861 62147 35017 62204
rect 50103 62250 50263 62310
rect 50103 62204 50160 62250
rect 50206 62204 50263 62250
rect 50103 62144 50263 62204
rect 56212 63066 56546 63188
rect 56212 63020 56267 63066
rect 56313 63020 56546 63066
rect 56212 62903 56546 63020
rect 56212 62857 56267 62903
rect 56313 62857 56546 62903
rect 56212 62740 56546 62857
rect 56212 62694 56267 62740
rect 56313 62694 56546 62740
rect 56212 62577 56546 62694
rect 56212 62531 56267 62577
rect 56313 62531 56546 62577
rect 56212 62413 56546 62531
rect 56212 62367 56267 62413
rect 56313 62367 56546 62413
rect 56212 62250 56546 62367
rect 56212 62204 56267 62250
rect 56313 62204 56546 62250
rect 28577 61220 28810 61266
rect 28856 61220 28911 61266
rect 28577 61103 28911 61220
rect 28577 61057 28810 61103
rect 28856 61057 28911 61103
rect 28577 60940 28911 61057
rect 28577 60894 28810 60940
rect 28856 60894 28911 60940
rect 28577 60777 28911 60894
rect 28577 60731 28810 60777
rect 28856 60731 28911 60777
rect 28577 60613 28911 60731
rect 28577 60567 28810 60613
rect 28856 60567 28911 60613
rect 28577 60450 28911 60567
rect 37938 61350 38492 61369
rect 37938 61304 37957 61350
rect 38473 61304 38492 61350
rect 37938 61285 38492 61304
rect 40779 61350 42995 61410
rect 40779 61304 40836 61350
rect 40882 61304 40994 61350
rect 41040 61304 41152 61350
rect 41198 61304 41310 61350
rect 41356 61304 41469 61350
rect 41515 61304 41627 61350
rect 41673 61304 41785 61350
rect 41831 61304 41943 61350
rect 41989 61304 42101 61350
rect 42147 61304 42259 61350
rect 42305 61304 42418 61350
rect 42464 61304 42576 61350
rect 42622 61304 42734 61350
rect 42780 61304 42892 61350
rect 42938 61304 42995 61350
rect 40779 61244 42995 61304
rect 56212 62087 56546 62204
rect 56212 62041 56267 62087
rect 56313 62041 56546 62087
rect 56212 61923 56546 62041
rect 56212 61877 56267 61923
rect 56313 61877 56546 61923
rect 56212 61760 56546 61877
rect 56212 61714 56267 61760
rect 56313 61714 56546 61760
rect 56212 61597 56546 61714
rect 56212 61551 56267 61597
rect 56313 61551 56546 61597
rect 56212 61434 56546 61551
rect 56212 61388 56267 61434
rect 56313 61388 56546 61434
rect 28577 60404 28810 60450
rect 28856 60404 28911 60450
rect 28577 60287 28911 60404
rect 28577 60241 28810 60287
rect 28856 60241 28911 60287
rect 28577 60123 28911 60241
rect 28577 60077 28810 60123
rect 28856 60077 28911 60123
rect 28577 59960 28911 60077
rect 28577 59914 28810 59960
rect 28856 59914 28911 59960
rect 28577 59797 28911 59914
rect 28577 59751 28810 59797
rect 28856 59751 28911 59797
rect 28577 59634 28911 59751
rect 28577 59588 28810 59634
rect 28856 59588 28911 59634
rect 28577 59466 28911 59588
rect 34861 60450 35017 60507
rect 34861 60404 34916 60450
rect 34962 60404 35017 60450
rect 34861 60347 35017 60404
rect 50103 60450 50263 60510
rect 50103 60404 50160 60450
rect 50206 60404 50263 60450
rect 50103 60344 50263 60404
rect 56212 61266 56546 61388
rect 56212 61220 56267 61266
rect 56313 61220 56546 61266
rect 56212 61103 56546 61220
rect 56212 61057 56267 61103
rect 56313 61057 56546 61103
rect 56212 60940 56546 61057
rect 56212 60894 56267 60940
rect 56313 60894 56546 60940
rect 56212 60777 56546 60894
rect 56212 60731 56267 60777
rect 56313 60731 56546 60777
rect 56212 60613 56546 60731
rect 56212 60567 56267 60613
rect 56313 60567 56546 60613
rect 56212 60450 56546 60567
rect 56212 60404 56267 60450
rect 56313 60404 56546 60450
rect 28577 59420 28810 59466
rect 28856 59420 28911 59466
rect 28577 59303 28911 59420
rect 28577 59257 28810 59303
rect 28856 59257 28911 59303
rect 28577 59140 28911 59257
rect 28577 59094 28810 59140
rect 28856 59094 28911 59140
rect 28577 58977 28911 59094
rect 28577 58931 28810 58977
rect 28856 58931 28911 58977
rect 28577 58813 28911 58931
rect 28577 58767 28810 58813
rect 28856 58767 28911 58813
rect 28577 58650 28911 58767
rect 37938 59550 38492 59569
rect 37938 59504 37957 59550
rect 38473 59504 38492 59550
rect 37938 59485 38492 59504
rect 40779 59550 42995 59610
rect 40779 59504 40836 59550
rect 40882 59504 40994 59550
rect 41040 59504 41152 59550
rect 41198 59504 41310 59550
rect 41356 59504 41469 59550
rect 41515 59504 41627 59550
rect 41673 59504 41785 59550
rect 41831 59504 41943 59550
rect 41989 59504 42101 59550
rect 42147 59504 42259 59550
rect 42305 59504 42418 59550
rect 42464 59504 42576 59550
rect 42622 59504 42734 59550
rect 42780 59504 42892 59550
rect 42938 59504 42995 59550
rect 40779 59444 42995 59504
rect 56212 60287 56546 60404
rect 56212 60241 56267 60287
rect 56313 60241 56546 60287
rect 56212 60123 56546 60241
rect 56212 60077 56267 60123
rect 56313 60077 56546 60123
rect 56212 59960 56546 60077
rect 56212 59914 56267 59960
rect 56313 59914 56546 59960
rect 56212 59797 56546 59914
rect 56212 59751 56267 59797
rect 56313 59751 56546 59797
rect 56212 59634 56546 59751
rect 56212 59588 56267 59634
rect 56313 59588 56546 59634
rect 28577 58604 28810 58650
rect 28856 58604 28911 58650
rect 28577 58487 28911 58604
rect 28577 58441 28810 58487
rect 28856 58441 28911 58487
rect 28577 58323 28911 58441
rect 28577 58277 28810 58323
rect 28856 58277 28911 58323
rect 28577 58160 28911 58277
rect 28577 58114 28810 58160
rect 28856 58114 28911 58160
rect 28577 57997 28911 58114
rect 28577 57951 28810 57997
rect 28856 57951 28911 57997
rect 28577 57834 28911 57951
rect 28577 57788 28810 57834
rect 28856 57788 28911 57834
rect 28577 57666 28911 57788
rect 34861 58650 35017 58707
rect 34861 58604 34916 58650
rect 34962 58604 35017 58650
rect 34861 58547 35017 58604
rect 50103 58650 50263 58710
rect 50103 58604 50160 58650
rect 50206 58604 50263 58650
rect 50103 58544 50263 58604
rect 56212 59466 56546 59588
rect 56212 59420 56267 59466
rect 56313 59420 56546 59466
rect 56212 59303 56546 59420
rect 56212 59257 56267 59303
rect 56313 59257 56546 59303
rect 56212 59140 56546 59257
rect 56212 59094 56267 59140
rect 56313 59094 56546 59140
rect 56212 58977 56546 59094
rect 56212 58931 56267 58977
rect 56313 58931 56546 58977
rect 56212 58813 56546 58931
rect 56212 58767 56267 58813
rect 56313 58767 56546 58813
rect 56212 58650 56546 58767
rect 56212 58604 56267 58650
rect 56313 58604 56546 58650
rect 28577 57620 28810 57666
rect 28856 57620 28911 57666
rect 28577 57503 28911 57620
rect 28577 57457 28810 57503
rect 28856 57457 28911 57503
rect 28577 57340 28911 57457
rect 28577 57294 28810 57340
rect 28856 57294 28911 57340
rect 28577 57177 28911 57294
rect 28577 57131 28810 57177
rect 28856 57131 28911 57177
rect 28577 57013 28911 57131
rect 28577 56967 28810 57013
rect 28856 56967 28911 57013
rect 28577 56850 28911 56967
rect 37938 57750 38492 57769
rect 37938 57704 37957 57750
rect 38473 57704 38492 57750
rect 37938 57685 38492 57704
rect 40779 57750 42995 57810
rect 40779 57704 40836 57750
rect 40882 57704 40994 57750
rect 41040 57704 41152 57750
rect 41198 57704 41310 57750
rect 41356 57704 41469 57750
rect 41515 57704 41627 57750
rect 41673 57704 41785 57750
rect 41831 57704 41943 57750
rect 41989 57704 42101 57750
rect 42147 57704 42259 57750
rect 42305 57704 42418 57750
rect 42464 57704 42576 57750
rect 42622 57704 42734 57750
rect 42780 57704 42892 57750
rect 42938 57704 42995 57750
rect 40779 57644 42995 57704
rect 56212 58487 56546 58604
rect 56212 58441 56267 58487
rect 56313 58441 56546 58487
rect 56212 58323 56546 58441
rect 56212 58277 56267 58323
rect 56313 58277 56546 58323
rect 56212 58160 56546 58277
rect 56212 58114 56267 58160
rect 56313 58114 56546 58160
rect 56212 57997 56546 58114
rect 56212 57951 56267 57997
rect 56313 57951 56546 57997
rect 56212 57834 56546 57951
rect 56212 57788 56267 57834
rect 56313 57788 56546 57834
rect 28577 56804 28810 56850
rect 28856 56804 28911 56850
rect 28577 56687 28911 56804
rect 28577 56641 28810 56687
rect 28856 56641 28911 56687
rect 28577 56523 28911 56641
rect 28577 56477 28810 56523
rect 28856 56477 28911 56523
rect 28577 56360 28911 56477
rect 28577 56314 28810 56360
rect 28856 56314 28911 56360
rect 28577 56197 28911 56314
rect 28577 56151 28810 56197
rect 28856 56151 28911 56197
rect 28577 56034 28911 56151
rect 28577 55988 28810 56034
rect 28856 55988 28911 56034
rect 28577 55866 28911 55988
rect 34861 56850 35017 56907
rect 34861 56804 34916 56850
rect 34962 56804 35017 56850
rect 34861 56747 35017 56804
rect 50103 56850 50263 56910
rect 50103 56804 50160 56850
rect 50206 56804 50263 56850
rect 50103 56744 50263 56804
rect 56212 57666 56546 57788
rect 56212 57620 56267 57666
rect 56313 57620 56546 57666
rect 56212 57503 56546 57620
rect 56212 57457 56267 57503
rect 56313 57457 56546 57503
rect 56212 57340 56546 57457
rect 56212 57294 56267 57340
rect 56313 57294 56546 57340
rect 56212 57177 56546 57294
rect 56212 57131 56267 57177
rect 56313 57131 56546 57177
rect 56212 57013 56546 57131
rect 56212 56967 56267 57013
rect 56313 56967 56546 57013
rect 56212 56850 56546 56967
rect 56212 56804 56267 56850
rect 56313 56804 56546 56850
rect 28577 55820 28810 55866
rect 28856 55820 28911 55866
rect 28577 55703 28911 55820
rect 28577 55657 28810 55703
rect 28856 55657 28911 55703
rect 28577 55540 28911 55657
rect 28577 55494 28810 55540
rect 28856 55494 28911 55540
rect 28577 55377 28911 55494
rect 28577 55331 28810 55377
rect 28856 55331 28911 55377
rect 28577 55213 28911 55331
rect 28577 55167 28810 55213
rect 28856 55167 28911 55213
rect 28577 55050 28911 55167
rect 37938 55950 38492 55969
rect 37938 55904 37957 55950
rect 38473 55904 38492 55950
rect 37938 55885 38492 55904
rect 40779 55950 42995 56010
rect 40779 55904 40836 55950
rect 40882 55904 40994 55950
rect 41040 55904 41152 55950
rect 41198 55904 41310 55950
rect 41356 55904 41469 55950
rect 41515 55904 41627 55950
rect 41673 55904 41785 55950
rect 41831 55904 41943 55950
rect 41989 55904 42101 55950
rect 42147 55904 42259 55950
rect 42305 55904 42418 55950
rect 42464 55904 42576 55950
rect 42622 55904 42734 55950
rect 42780 55904 42892 55950
rect 42938 55904 42995 55950
rect 40779 55844 42995 55904
rect 56212 56687 56546 56804
rect 56212 56641 56267 56687
rect 56313 56641 56546 56687
rect 56212 56523 56546 56641
rect 56212 56477 56267 56523
rect 56313 56477 56546 56523
rect 56212 56360 56546 56477
rect 56212 56314 56267 56360
rect 56313 56314 56546 56360
rect 56212 56197 56546 56314
rect 56212 56151 56267 56197
rect 56313 56151 56546 56197
rect 56212 56034 56546 56151
rect 56212 55988 56267 56034
rect 56313 55988 56546 56034
rect 28577 55004 28810 55050
rect 28856 55004 28911 55050
rect 28577 54887 28911 55004
rect 28577 54841 28810 54887
rect 28856 54841 28911 54887
rect 28577 54723 28911 54841
rect 28577 54677 28810 54723
rect 28856 54677 28911 54723
rect 28577 54560 28911 54677
rect 28577 54514 28810 54560
rect 28856 54514 28911 54560
rect 28577 54397 28911 54514
rect 28577 54351 28810 54397
rect 28856 54351 28911 54397
rect 28577 54234 28911 54351
rect 28577 54188 28810 54234
rect 28856 54188 28911 54234
rect 28577 54066 28911 54188
rect 34861 55050 35017 55107
rect 34861 55004 34916 55050
rect 34962 55004 35017 55050
rect 34861 54947 35017 55004
rect 50103 55050 50263 55110
rect 50103 55004 50160 55050
rect 50206 55004 50263 55050
rect 50103 54944 50263 55004
rect 56212 55866 56546 55988
rect 56212 55820 56267 55866
rect 56313 55820 56546 55866
rect 56212 55703 56546 55820
rect 56212 55657 56267 55703
rect 56313 55657 56546 55703
rect 56212 55540 56546 55657
rect 56212 55494 56267 55540
rect 56313 55494 56546 55540
rect 56212 55377 56546 55494
rect 56212 55331 56267 55377
rect 56313 55331 56546 55377
rect 56212 55213 56546 55331
rect 56212 55167 56267 55213
rect 56313 55167 56546 55213
rect 56212 55050 56546 55167
rect 56212 55004 56267 55050
rect 56313 55004 56546 55050
rect 28577 54020 28810 54066
rect 28856 54020 28911 54066
rect 28577 53903 28911 54020
rect 28577 53857 28810 53903
rect 28856 53857 28911 53903
rect 28577 53740 28911 53857
rect 28577 53694 28810 53740
rect 28856 53694 28911 53740
rect 28577 53577 28911 53694
rect 28577 53531 28810 53577
rect 28856 53531 28911 53577
rect 28577 53413 28911 53531
rect 28577 53367 28810 53413
rect 28856 53367 28911 53413
rect 28577 53250 28911 53367
rect 37938 54150 38492 54169
rect 37938 54104 37957 54150
rect 38473 54104 38492 54150
rect 37938 54085 38492 54104
rect 40779 54150 42995 54210
rect 40779 54104 40836 54150
rect 40882 54104 40994 54150
rect 41040 54104 41152 54150
rect 41198 54104 41310 54150
rect 41356 54104 41469 54150
rect 41515 54104 41627 54150
rect 41673 54104 41785 54150
rect 41831 54104 41943 54150
rect 41989 54104 42101 54150
rect 42147 54104 42259 54150
rect 42305 54104 42418 54150
rect 42464 54104 42576 54150
rect 42622 54104 42734 54150
rect 42780 54104 42892 54150
rect 42938 54104 42995 54150
rect 40779 54044 42995 54104
rect 56212 54887 56546 55004
rect 56212 54841 56267 54887
rect 56313 54841 56546 54887
rect 56212 54723 56546 54841
rect 56212 54677 56267 54723
rect 56313 54677 56546 54723
rect 56212 54560 56546 54677
rect 56212 54514 56267 54560
rect 56313 54514 56546 54560
rect 56212 54397 56546 54514
rect 56212 54351 56267 54397
rect 56313 54351 56546 54397
rect 56212 54234 56546 54351
rect 56212 54188 56267 54234
rect 56313 54188 56546 54234
rect 28577 53204 28810 53250
rect 28856 53204 28911 53250
rect 28577 53087 28911 53204
rect 28577 53041 28810 53087
rect 28856 53041 28911 53087
rect 28577 52923 28911 53041
rect 28577 52877 28810 52923
rect 28856 52877 28911 52923
rect 28577 52760 28911 52877
rect 28577 52714 28810 52760
rect 28856 52714 28911 52760
rect 28577 52597 28911 52714
rect 28577 52551 28810 52597
rect 28856 52551 28911 52597
rect 28577 52434 28911 52551
rect 28577 52388 28810 52434
rect 28856 52388 28911 52434
rect 28577 52266 28911 52388
rect 34861 53250 35017 53307
rect 34861 53204 34916 53250
rect 34962 53204 35017 53250
rect 34861 53147 35017 53204
rect 50103 53250 50263 53310
rect 50103 53204 50160 53250
rect 50206 53204 50263 53250
rect 50103 53144 50263 53204
rect 56212 54066 56546 54188
rect 56212 54020 56267 54066
rect 56313 54020 56546 54066
rect 56212 53903 56546 54020
rect 56212 53857 56267 53903
rect 56313 53857 56546 53903
rect 56212 53740 56546 53857
rect 56212 53694 56267 53740
rect 56313 53694 56546 53740
rect 56212 53577 56546 53694
rect 56212 53531 56267 53577
rect 56313 53531 56546 53577
rect 56212 53413 56546 53531
rect 56212 53367 56267 53413
rect 56313 53367 56546 53413
rect 56212 53250 56546 53367
rect 56212 53204 56267 53250
rect 56313 53204 56546 53250
rect 28577 52220 28810 52266
rect 28856 52220 28911 52266
rect 28577 52103 28911 52220
rect 28577 52057 28810 52103
rect 28856 52057 28911 52103
rect 28577 51940 28911 52057
rect 28577 51894 28810 51940
rect 28856 51894 28911 51940
rect 28577 51777 28911 51894
rect 28577 51731 28810 51777
rect 28856 51731 28911 51777
rect 28577 51613 28911 51731
rect 28577 51567 28810 51613
rect 28856 51567 28911 51613
rect 28577 51450 28911 51567
rect 37938 52350 38492 52369
rect 37938 52304 37957 52350
rect 38473 52304 38492 52350
rect 37938 52285 38492 52304
rect 40779 52350 42995 52410
rect 40779 52304 40836 52350
rect 40882 52304 40994 52350
rect 41040 52304 41152 52350
rect 41198 52304 41310 52350
rect 41356 52304 41469 52350
rect 41515 52304 41627 52350
rect 41673 52304 41785 52350
rect 41831 52304 41943 52350
rect 41989 52304 42101 52350
rect 42147 52304 42259 52350
rect 42305 52304 42418 52350
rect 42464 52304 42576 52350
rect 42622 52304 42734 52350
rect 42780 52304 42892 52350
rect 42938 52304 42995 52350
rect 40779 52244 42995 52304
rect 56212 53087 56546 53204
rect 56212 53041 56267 53087
rect 56313 53041 56546 53087
rect 56212 52923 56546 53041
rect 56212 52877 56267 52923
rect 56313 52877 56546 52923
rect 56212 52760 56546 52877
rect 56212 52714 56267 52760
rect 56313 52714 56546 52760
rect 56212 52597 56546 52714
rect 56212 52551 56267 52597
rect 56313 52551 56546 52597
rect 56212 52434 56546 52551
rect 56212 52388 56267 52434
rect 56313 52388 56546 52434
rect 28577 51404 28810 51450
rect 28856 51404 28911 51450
rect 28577 51287 28911 51404
rect 28577 51241 28810 51287
rect 28856 51241 28911 51287
rect 28577 51123 28911 51241
rect 28577 51077 28810 51123
rect 28856 51077 28911 51123
rect 28577 50960 28911 51077
rect 28577 50914 28810 50960
rect 28856 50914 28911 50960
rect 28577 50797 28911 50914
rect 28577 50751 28810 50797
rect 28856 50751 28911 50797
rect 28577 50634 28911 50751
rect 28577 50588 28810 50634
rect 28856 50588 28911 50634
rect 28577 50466 28911 50588
rect 34861 51450 35017 51507
rect 34861 51404 34916 51450
rect 34962 51404 35017 51450
rect 34861 51347 35017 51404
rect 50103 51450 50263 51510
rect 50103 51404 50160 51450
rect 50206 51404 50263 51450
rect 50103 51344 50263 51404
rect 56212 52266 56546 52388
rect 56212 52220 56267 52266
rect 56313 52220 56546 52266
rect 56212 52103 56546 52220
rect 56212 52057 56267 52103
rect 56313 52057 56546 52103
rect 56212 51940 56546 52057
rect 56212 51894 56267 51940
rect 56313 51894 56546 51940
rect 56212 51777 56546 51894
rect 56212 51731 56267 51777
rect 56313 51731 56546 51777
rect 56212 51613 56546 51731
rect 56212 51567 56267 51613
rect 56313 51567 56546 51613
rect 56212 51450 56546 51567
rect 56212 51404 56267 51450
rect 56313 51404 56546 51450
rect 28577 50420 28810 50466
rect 28856 50420 28911 50466
rect 28577 50303 28911 50420
rect 28577 50257 28810 50303
rect 28856 50257 28911 50303
rect 28577 50140 28911 50257
rect 28577 50094 28810 50140
rect 28856 50094 28911 50140
rect 28577 49977 28911 50094
rect 28577 49931 28810 49977
rect 28856 49931 28911 49977
rect 28577 49813 28911 49931
rect 28577 49767 28810 49813
rect 28856 49767 28911 49813
rect 28577 49650 28911 49767
rect 37938 50550 38492 50569
rect 37938 50504 37957 50550
rect 38473 50504 38492 50550
rect 37938 50485 38492 50504
rect 40779 50550 42995 50610
rect 40779 50504 40836 50550
rect 40882 50504 40994 50550
rect 41040 50504 41152 50550
rect 41198 50504 41310 50550
rect 41356 50504 41469 50550
rect 41515 50504 41627 50550
rect 41673 50504 41785 50550
rect 41831 50504 41943 50550
rect 41989 50504 42101 50550
rect 42147 50504 42259 50550
rect 42305 50504 42418 50550
rect 42464 50504 42576 50550
rect 42622 50504 42734 50550
rect 42780 50504 42892 50550
rect 42938 50504 42995 50550
rect 40779 50444 42995 50504
rect 56212 51287 56546 51404
rect 56212 51241 56267 51287
rect 56313 51241 56546 51287
rect 56212 51123 56546 51241
rect 56212 51077 56267 51123
rect 56313 51077 56546 51123
rect 56212 50960 56546 51077
rect 56212 50914 56267 50960
rect 56313 50914 56546 50960
rect 56212 50797 56546 50914
rect 56212 50751 56267 50797
rect 56313 50751 56546 50797
rect 56212 50634 56546 50751
rect 56212 50588 56267 50634
rect 56313 50588 56546 50634
rect 28577 49604 28810 49650
rect 28856 49604 28911 49650
rect 28577 49487 28911 49604
rect 28577 49441 28810 49487
rect 28856 49441 28911 49487
rect 28577 49323 28911 49441
rect 28577 49277 28810 49323
rect 28856 49277 28911 49323
rect 28577 49160 28911 49277
rect 28577 49114 28810 49160
rect 28856 49114 28911 49160
rect 28577 48997 28911 49114
rect 28577 48951 28810 48997
rect 28856 48951 28911 48997
rect 28577 48834 28911 48951
rect 28577 48788 28810 48834
rect 28856 48788 28911 48834
rect 28577 48666 28911 48788
rect 34861 49650 35017 49707
rect 34861 49604 34916 49650
rect 34962 49604 35017 49650
rect 34861 49547 35017 49604
rect 50103 49650 50263 49710
rect 50103 49604 50160 49650
rect 50206 49604 50263 49650
rect 50103 49544 50263 49604
rect 56212 50466 56546 50588
rect 56212 50420 56267 50466
rect 56313 50420 56546 50466
rect 56212 50303 56546 50420
rect 56212 50257 56267 50303
rect 56313 50257 56546 50303
rect 56212 50140 56546 50257
rect 56212 50094 56267 50140
rect 56313 50094 56546 50140
rect 56212 49977 56546 50094
rect 56212 49931 56267 49977
rect 56313 49931 56546 49977
rect 56212 49813 56546 49931
rect 56212 49767 56267 49813
rect 56313 49767 56546 49813
rect 56212 49650 56546 49767
rect 56212 49604 56267 49650
rect 56313 49604 56546 49650
rect 28577 48620 28810 48666
rect 28856 48620 28911 48666
rect 28577 48503 28911 48620
rect 28577 48457 28810 48503
rect 28856 48457 28911 48503
rect 28577 48340 28911 48457
rect 28577 48294 28810 48340
rect 28856 48294 28911 48340
rect 28577 48177 28911 48294
rect 28577 48131 28810 48177
rect 28856 48131 28911 48177
rect 28577 48013 28911 48131
rect 28577 47967 28810 48013
rect 28856 47967 28911 48013
rect 28577 47850 28911 47967
rect 37938 48750 38492 48769
rect 37938 48704 37957 48750
rect 38473 48704 38492 48750
rect 37938 48685 38492 48704
rect 40779 48750 42995 48810
rect 40779 48704 40836 48750
rect 40882 48704 40994 48750
rect 41040 48704 41152 48750
rect 41198 48704 41310 48750
rect 41356 48704 41469 48750
rect 41515 48704 41627 48750
rect 41673 48704 41785 48750
rect 41831 48704 41943 48750
rect 41989 48704 42101 48750
rect 42147 48704 42259 48750
rect 42305 48704 42418 48750
rect 42464 48704 42576 48750
rect 42622 48704 42734 48750
rect 42780 48704 42892 48750
rect 42938 48704 42995 48750
rect 40779 48644 42995 48704
rect 56212 49487 56546 49604
rect 56212 49441 56267 49487
rect 56313 49441 56546 49487
rect 56212 49323 56546 49441
rect 56212 49277 56267 49323
rect 56313 49277 56546 49323
rect 56212 49160 56546 49277
rect 56212 49114 56267 49160
rect 56313 49114 56546 49160
rect 56212 48997 56546 49114
rect 56212 48951 56267 48997
rect 56313 48951 56546 48997
rect 56212 48834 56546 48951
rect 56212 48788 56267 48834
rect 56313 48788 56546 48834
rect 28577 47804 28810 47850
rect 28856 47804 28911 47850
rect 28577 47687 28911 47804
rect 28577 47641 28810 47687
rect 28856 47641 28911 47687
rect 28577 47523 28911 47641
rect 28577 47477 28810 47523
rect 28856 47477 28911 47523
rect 28577 47360 28911 47477
rect 28577 47314 28810 47360
rect 28856 47314 28911 47360
rect 28577 47197 28911 47314
rect 28577 47151 28810 47197
rect 28856 47151 28911 47197
rect 28577 47034 28911 47151
rect 28577 46988 28810 47034
rect 28856 46988 28911 47034
rect 28577 46866 28911 46988
rect 34861 47850 35017 47907
rect 34861 47804 34916 47850
rect 34962 47804 35017 47850
rect 34861 47747 35017 47804
rect 50103 47850 50263 47910
rect 50103 47804 50160 47850
rect 50206 47804 50263 47850
rect 50103 47744 50263 47804
rect 56212 48666 56546 48788
rect 56212 48620 56267 48666
rect 56313 48620 56546 48666
rect 56212 48503 56546 48620
rect 56212 48457 56267 48503
rect 56313 48457 56546 48503
rect 56212 48340 56546 48457
rect 56212 48294 56267 48340
rect 56313 48294 56546 48340
rect 56212 48177 56546 48294
rect 56212 48131 56267 48177
rect 56313 48131 56546 48177
rect 56212 48013 56546 48131
rect 56212 47967 56267 48013
rect 56313 47967 56546 48013
rect 56212 47850 56546 47967
rect 56212 47804 56267 47850
rect 56313 47804 56546 47850
rect 28577 46820 28810 46866
rect 28856 46820 28911 46866
rect 28577 46703 28911 46820
rect 28577 46657 28810 46703
rect 28856 46657 28911 46703
rect 28577 46540 28911 46657
rect 28577 46494 28810 46540
rect 28856 46494 28911 46540
rect 28577 46377 28911 46494
rect 28577 46331 28810 46377
rect 28856 46331 28911 46377
rect 28577 46213 28911 46331
rect 28577 46167 28810 46213
rect 28856 46167 28911 46213
rect 28577 46050 28911 46167
rect 37938 46950 38492 46969
rect 37938 46904 37957 46950
rect 38473 46904 38492 46950
rect 37938 46885 38492 46904
rect 40779 46950 42995 47010
rect 40779 46904 40836 46950
rect 40882 46904 40994 46950
rect 41040 46904 41152 46950
rect 41198 46904 41310 46950
rect 41356 46904 41469 46950
rect 41515 46904 41627 46950
rect 41673 46904 41785 46950
rect 41831 46904 41943 46950
rect 41989 46904 42101 46950
rect 42147 46904 42259 46950
rect 42305 46904 42418 46950
rect 42464 46904 42576 46950
rect 42622 46904 42734 46950
rect 42780 46904 42892 46950
rect 42938 46904 42995 46950
rect 40779 46844 42995 46904
rect 56212 47687 56546 47804
rect 56212 47641 56267 47687
rect 56313 47641 56546 47687
rect 56212 47523 56546 47641
rect 56212 47477 56267 47523
rect 56313 47477 56546 47523
rect 56212 47360 56546 47477
rect 56212 47314 56267 47360
rect 56313 47314 56546 47360
rect 56212 47197 56546 47314
rect 56212 47151 56267 47197
rect 56313 47151 56546 47197
rect 56212 47034 56546 47151
rect 56212 46988 56267 47034
rect 56313 46988 56546 47034
rect 28577 46004 28810 46050
rect 28856 46004 28911 46050
rect 28577 45887 28911 46004
rect 28577 45841 28810 45887
rect 28856 45841 28911 45887
rect 28577 45723 28911 45841
rect 28577 45677 28810 45723
rect 28856 45677 28911 45723
rect 28577 45560 28911 45677
rect 28577 45514 28810 45560
rect 28856 45514 28911 45560
rect 28577 45397 28911 45514
rect 28577 45351 28810 45397
rect 28856 45351 28911 45397
rect 28577 45234 28911 45351
rect 28577 45188 28810 45234
rect 28856 45188 28911 45234
rect 28577 45066 28911 45188
rect 34861 46050 35017 46107
rect 34861 46004 34916 46050
rect 34962 46004 35017 46050
rect 34861 45947 35017 46004
rect 50103 46050 50263 46110
rect 50103 46004 50160 46050
rect 50206 46004 50263 46050
rect 50103 45944 50263 46004
rect 56212 46866 56546 46988
rect 56212 46820 56267 46866
rect 56313 46820 56546 46866
rect 56212 46703 56546 46820
rect 56212 46657 56267 46703
rect 56313 46657 56546 46703
rect 56212 46540 56546 46657
rect 56212 46494 56267 46540
rect 56313 46494 56546 46540
rect 56212 46377 56546 46494
rect 56212 46331 56267 46377
rect 56313 46331 56546 46377
rect 56212 46213 56546 46331
rect 56212 46167 56267 46213
rect 56313 46167 56546 46213
rect 56212 46050 56546 46167
rect 56212 46004 56267 46050
rect 56313 46004 56546 46050
rect 28577 45020 28810 45066
rect 28856 45020 28911 45066
rect 28577 44903 28911 45020
rect 28577 44857 28810 44903
rect 28856 44857 28911 44903
rect 28577 44740 28911 44857
rect 28577 44694 28810 44740
rect 28856 44694 28911 44740
rect 28577 44577 28911 44694
rect 28577 44531 28810 44577
rect 28856 44531 28911 44577
rect 28577 44413 28911 44531
rect 28577 44367 28810 44413
rect 28856 44367 28911 44413
rect 28577 44250 28911 44367
rect 37938 45150 38492 45169
rect 37938 45104 37957 45150
rect 38473 45104 38492 45150
rect 37938 45085 38492 45104
rect 40779 45150 42995 45210
rect 40779 45104 40836 45150
rect 40882 45104 40994 45150
rect 41040 45104 41152 45150
rect 41198 45104 41310 45150
rect 41356 45104 41469 45150
rect 41515 45104 41627 45150
rect 41673 45104 41785 45150
rect 41831 45104 41943 45150
rect 41989 45104 42101 45150
rect 42147 45104 42259 45150
rect 42305 45104 42418 45150
rect 42464 45104 42576 45150
rect 42622 45104 42734 45150
rect 42780 45104 42892 45150
rect 42938 45104 42995 45150
rect 40779 45044 42995 45104
rect 56212 45887 56546 46004
rect 56212 45841 56267 45887
rect 56313 45841 56546 45887
rect 56212 45723 56546 45841
rect 56212 45677 56267 45723
rect 56313 45677 56546 45723
rect 56212 45560 56546 45677
rect 56212 45514 56267 45560
rect 56313 45514 56546 45560
rect 56212 45397 56546 45514
rect 56212 45351 56267 45397
rect 56313 45351 56546 45397
rect 56212 45234 56546 45351
rect 56212 45188 56267 45234
rect 56313 45188 56546 45234
rect 28577 44204 28810 44250
rect 28856 44204 28911 44250
rect 28577 44087 28911 44204
rect 28577 44041 28810 44087
rect 28856 44041 28911 44087
rect 28577 43923 28911 44041
rect 28577 43877 28810 43923
rect 28856 43877 28911 43923
rect 28577 43760 28911 43877
rect 28577 43714 28810 43760
rect 28856 43714 28911 43760
rect 28577 43597 28911 43714
rect 28577 43551 28810 43597
rect 28856 43551 28911 43597
rect 28577 43434 28911 43551
rect 28577 43388 28810 43434
rect 28856 43388 28911 43434
rect 28577 43266 28911 43388
rect 34861 44250 35017 44307
rect 34861 44204 34916 44250
rect 34962 44204 35017 44250
rect 34861 44147 35017 44204
rect 50103 44250 50263 44310
rect 50103 44204 50160 44250
rect 50206 44204 50263 44250
rect 50103 44144 50263 44204
rect 56212 45066 56546 45188
rect 56212 45020 56267 45066
rect 56313 45020 56546 45066
rect 56212 44903 56546 45020
rect 56212 44857 56267 44903
rect 56313 44857 56546 44903
rect 56212 44740 56546 44857
rect 56212 44694 56267 44740
rect 56313 44694 56546 44740
rect 56212 44577 56546 44694
rect 56212 44531 56267 44577
rect 56313 44531 56546 44577
rect 56212 44413 56546 44531
rect 56212 44367 56267 44413
rect 56313 44367 56546 44413
rect 56212 44250 56546 44367
rect 56212 44204 56267 44250
rect 56313 44204 56546 44250
rect 28577 43220 28810 43266
rect 28856 43220 28911 43266
rect 28577 43103 28911 43220
rect 28577 43057 28810 43103
rect 28856 43057 28911 43103
rect 28577 42940 28911 43057
rect 28577 42894 28810 42940
rect 28856 42894 28911 42940
rect 28577 42777 28911 42894
rect 28577 42731 28810 42777
rect 28856 42731 28911 42777
rect 28577 42613 28911 42731
rect 28577 42567 28810 42613
rect 28856 42567 28911 42613
rect 28577 42450 28911 42567
rect 37938 43350 38492 43369
rect 37938 43304 37957 43350
rect 38473 43304 38492 43350
rect 37938 43285 38492 43304
rect 40779 43350 42995 43410
rect 40779 43304 40836 43350
rect 40882 43304 40994 43350
rect 41040 43304 41152 43350
rect 41198 43304 41310 43350
rect 41356 43304 41469 43350
rect 41515 43304 41627 43350
rect 41673 43304 41785 43350
rect 41831 43304 41943 43350
rect 41989 43304 42101 43350
rect 42147 43304 42259 43350
rect 42305 43304 42418 43350
rect 42464 43304 42576 43350
rect 42622 43304 42734 43350
rect 42780 43304 42892 43350
rect 42938 43304 42995 43350
rect 40779 43244 42995 43304
rect 56212 44087 56546 44204
rect 56212 44041 56267 44087
rect 56313 44041 56546 44087
rect 56212 43923 56546 44041
rect 56212 43877 56267 43923
rect 56313 43877 56546 43923
rect 56212 43760 56546 43877
rect 56212 43714 56267 43760
rect 56313 43714 56546 43760
rect 56212 43597 56546 43714
rect 56212 43551 56267 43597
rect 56313 43551 56546 43597
rect 56212 43434 56546 43551
rect 56212 43388 56267 43434
rect 56313 43388 56546 43434
rect 28577 42404 28810 42450
rect 28856 42404 28911 42450
rect 28577 42287 28911 42404
rect 28577 42241 28810 42287
rect 28856 42241 28911 42287
rect 28577 42123 28911 42241
rect 28577 42077 28810 42123
rect 28856 42077 28911 42123
rect 28577 41960 28911 42077
rect 28577 41914 28810 41960
rect 28856 41914 28911 41960
rect 28577 41797 28911 41914
rect 28577 41751 28810 41797
rect 28856 41751 28911 41797
rect 28577 41634 28911 41751
rect 28577 41588 28810 41634
rect 28856 41588 28911 41634
rect 28577 41466 28911 41588
rect 34861 42450 35017 42507
rect 34861 42404 34916 42450
rect 34962 42404 35017 42450
rect 34861 42347 35017 42404
rect 50103 42450 50263 42510
rect 50103 42404 50160 42450
rect 50206 42404 50263 42450
rect 50103 42344 50263 42404
rect 56212 43266 56546 43388
rect 56212 43220 56267 43266
rect 56313 43220 56546 43266
rect 56212 43103 56546 43220
rect 56212 43057 56267 43103
rect 56313 43057 56546 43103
rect 56212 42940 56546 43057
rect 56212 42894 56267 42940
rect 56313 42894 56546 42940
rect 56212 42777 56546 42894
rect 56212 42731 56267 42777
rect 56313 42731 56546 42777
rect 56212 42613 56546 42731
rect 56212 42567 56267 42613
rect 56313 42567 56546 42613
rect 56212 42450 56546 42567
rect 56212 42404 56267 42450
rect 56313 42404 56546 42450
rect 28577 41420 28810 41466
rect 28856 41420 28911 41466
rect 28577 41303 28911 41420
rect 28577 41257 28810 41303
rect 28856 41257 28911 41303
rect 28577 41140 28911 41257
rect 28577 41094 28810 41140
rect 28856 41094 28911 41140
rect 28577 40977 28911 41094
rect 28577 40931 28810 40977
rect 28856 40931 28911 40977
rect 28577 40813 28911 40931
rect 28577 40767 28810 40813
rect 28856 40767 28911 40813
rect 28577 40650 28911 40767
rect 37938 41550 38492 41569
rect 37938 41504 37957 41550
rect 38473 41504 38492 41550
rect 37938 41485 38492 41504
rect 40779 41550 42995 41610
rect 40779 41504 40836 41550
rect 40882 41504 40994 41550
rect 41040 41504 41152 41550
rect 41198 41504 41310 41550
rect 41356 41504 41469 41550
rect 41515 41504 41627 41550
rect 41673 41504 41785 41550
rect 41831 41504 41943 41550
rect 41989 41504 42101 41550
rect 42147 41504 42259 41550
rect 42305 41504 42418 41550
rect 42464 41504 42576 41550
rect 42622 41504 42734 41550
rect 42780 41504 42892 41550
rect 42938 41504 42995 41550
rect 40779 41444 42995 41504
rect 56212 42287 56546 42404
rect 56212 42241 56267 42287
rect 56313 42241 56546 42287
rect 56212 42123 56546 42241
rect 56212 42077 56267 42123
rect 56313 42077 56546 42123
rect 56212 41960 56546 42077
rect 56212 41914 56267 41960
rect 56313 41914 56546 41960
rect 56212 41797 56546 41914
rect 56212 41751 56267 41797
rect 56313 41751 56546 41797
rect 56212 41634 56546 41751
rect 56212 41588 56267 41634
rect 56313 41588 56546 41634
rect 28577 40604 28810 40650
rect 28856 40604 28911 40650
rect 28577 40487 28911 40604
rect 28577 40441 28810 40487
rect 28856 40441 28911 40487
rect 28577 40323 28911 40441
rect 28577 40277 28810 40323
rect 28856 40277 28911 40323
rect 28577 40160 28911 40277
rect 28577 40114 28810 40160
rect 28856 40114 28911 40160
rect 28577 39997 28911 40114
rect 28577 39951 28810 39997
rect 28856 39951 28911 39997
rect 28577 39834 28911 39951
rect 28577 39788 28810 39834
rect 28856 39788 28911 39834
rect 28577 39666 28911 39788
rect 34861 40650 35017 40707
rect 34861 40604 34916 40650
rect 34962 40604 35017 40650
rect 34861 40547 35017 40604
rect 50103 40650 50263 40710
rect 50103 40604 50160 40650
rect 50206 40604 50263 40650
rect 50103 40544 50263 40604
rect 56212 41466 56546 41588
rect 56212 41420 56267 41466
rect 56313 41420 56546 41466
rect 56212 41303 56546 41420
rect 56212 41257 56267 41303
rect 56313 41257 56546 41303
rect 56212 41140 56546 41257
rect 56212 41094 56267 41140
rect 56313 41094 56546 41140
rect 56212 40977 56546 41094
rect 56212 40931 56267 40977
rect 56313 40931 56546 40977
rect 56212 40813 56546 40931
rect 56212 40767 56267 40813
rect 56313 40767 56546 40813
rect 56212 40650 56546 40767
rect 56212 40604 56267 40650
rect 56313 40604 56546 40650
rect 28577 39620 28810 39666
rect 28856 39620 28911 39666
rect 28577 39503 28911 39620
rect 28577 39457 28810 39503
rect 28856 39457 28911 39503
rect 28577 39340 28911 39457
rect 28577 39294 28810 39340
rect 28856 39294 28911 39340
rect 28577 39177 28911 39294
rect 28577 39131 28810 39177
rect 28856 39131 28911 39177
rect 28577 39013 28911 39131
rect 28577 38967 28810 39013
rect 28856 38967 28911 39013
rect 28577 38850 28911 38967
rect 37938 39750 38492 39769
rect 37938 39704 37957 39750
rect 38473 39704 38492 39750
rect 37938 39685 38492 39704
rect 40779 39750 42995 39810
rect 40779 39704 40836 39750
rect 40882 39704 40994 39750
rect 41040 39704 41152 39750
rect 41198 39704 41310 39750
rect 41356 39704 41469 39750
rect 41515 39704 41627 39750
rect 41673 39704 41785 39750
rect 41831 39704 41943 39750
rect 41989 39704 42101 39750
rect 42147 39704 42259 39750
rect 42305 39704 42418 39750
rect 42464 39704 42576 39750
rect 42622 39704 42734 39750
rect 42780 39704 42892 39750
rect 42938 39704 42995 39750
rect 40779 39644 42995 39704
rect 56212 40487 56546 40604
rect 56212 40441 56267 40487
rect 56313 40441 56546 40487
rect 56212 40323 56546 40441
rect 56212 40277 56267 40323
rect 56313 40277 56546 40323
rect 56212 40160 56546 40277
rect 56212 40114 56267 40160
rect 56313 40114 56546 40160
rect 56212 39997 56546 40114
rect 56212 39951 56267 39997
rect 56313 39951 56546 39997
rect 56212 39834 56546 39951
rect 56212 39788 56267 39834
rect 56313 39788 56546 39834
rect 28577 38804 28810 38850
rect 28856 38804 28911 38850
rect 28577 38687 28911 38804
rect 28577 38641 28810 38687
rect 28856 38641 28911 38687
rect 28577 38523 28911 38641
rect 28577 38477 28810 38523
rect 28856 38477 28911 38523
rect 28577 38360 28911 38477
rect 28577 38314 28810 38360
rect 28856 38314 28911 38360
rect 28577 38197 28911 38314
rect 28577 38151 28810 38197
rect 28856 38151 28911 38197
rect 28577 38034 28911 38151
rect 28577 37988 28810 38034
rect 28856 37988 28911 38034
rect 28577 37866 28911 37988
rect 34861 38850 35017 38907
rect 34861 38804 34916 38850
rect 34962 38804 35017 38850
rect 34861 38747 35017 38804
rect 50103 38850 50263 38910
rect 50103 38804 50160 38850
rect 50206 38804 50263 38850
rect 50103 38744 50263 38804
rect 56212 39666 56546 39788
rect 56212 39620 56267 39666
rect 56313 39620 56546 39666
rect 56212 39503 56546 39620
rect 56212 39457 56267 39503
rect 56313 39457 56546 39503
rect 56212 39340 56546 39457
rect 56212 39294 56267 39340
rect 56313 39294 56546 39340
rect 56212 39177 56546 39294
rect 56212 39131 56267 39177
rect 56313 39131 56546 39177
rect 56212 39013 56546 39131
rect 56212 38967 56267 39013
rect 56313 38967 56546 39013
rect 56212 38850 56546 38967
rect 56212 38804 56267 38850
rect 56313 38804 56546 38850
rect 28577 37820 28810 37866
rect 28856 37820 28911 37866
rect 28577 37703 28911 37820
rect 28577 37657 28810 37703
rect 28856 37657 28911 37703
rect 28577 37540 28911 37657
rect 28577 37494 28810 37540
rect 28856 37494 28911 37540
rect 28577 37377 28911 37494
rect 28577 37331 28810 37377
rect 28856 37331 28911 37377
rect 28577 37213 28911 37331
rect 28577 37167 28810 37213
rect 28856 37167 28911 37213
rect 28577 37050 28911 37167
rect 37938 37950 38492 37969
rect 37938 37904 37957 37950
rect 38473 37904 38492 37950
rect 37938 37885 38492 37904
rect 40779 37950 42995 38010
rect 40779 37904 40836 37950
rect 40882 37904 40994 37950
rect 41040 37904 41152 37950
rect 41198 37904 41310 37950
rect 41356 37904 41469 37950
rect 41515 37904 41627 37950
rect 41673 37904 41785 37950
rect 41831 37904 41943 37950
rect 41989 37904 42101 37950
rect 42147 37904 42259 37950
rect 42305 37904 42418 37950
rect 42464 37904 42576 37950
rect 42622 37904 42734 37950
rect 42780 37904 42892 37950
rect 42938 37904 42995 37950
rect 40779 37844 42995 37904
rect 56212 38687 56546 38804
rect 56212 38641 56267 38687
rect 56313 38641 56546 38687
rect 56212 38523 56546 38641
rect 56212 38477 56267 38523
rect 56313 38477 56546 38523
rect 56212 38360 56546 38477
rect 56212 38314 56267 38360
rect 56313 38314 56546 38360
rect 56212 38197 56546 38314
rect 56212 38151 56267 38197
rect 56313 38151 56546 38197
rect 56212 38034 56546 38151
rect 56212 37988 56267 38034
rect 56313 37988 56546 38034
rect 28577 37004 28810 37050
rect 28856 37004 28911 37050
rect 28577 36887 28911 37004
rect 28577 36841 28810 36887
rect 28856 36841 28911 36887
rect 28577 36723 28911 36841
rect 28577 36677 28810 36723
rect 28856 36677 28911 36723
rect 28577 36560 28911 36677
rect 28577 36514 28810 36560
rect 28856 36514 28911 36560
rect 28577 36397 28911 36514
rect 28577 36351 28810 36397
rect 28856 36351 28911 36397
rect 28577 36234 28911 36351
rect 28577 36188 28810 36234
rect 28856 36188 28911 36234
rect 28577 35977 28911 36188
rect 34861 37050 35017 37107
rect 34861 37004 34916 37050
rect 34962 37004 35017 37050
rect 34861 36947 35017 37004
rect 50103 37050 50263 37110
rect 50103 37004 50160 37050
rect 50206 37004 50263 37050
rect 50103 36944 50263 37004
rect 56212 37866 56546 37988
rect 56212 37820 56267 37866
rect 56313 37820 56546 37866
rect 56212 37703 56546 37820
rect 56212 37657 56267 37703
rect 56313 37657 56546 37703
rect 56212 37540 56546 37657
rect 56212 37494 56267 37540
rect 56313 37494 56546 37540
rect 56212 37377 56546 37494
rect 56212 37331 56267 37377
rect 56313 37331 56546 37377
rect 56212 37213 56546 37331
rect 56212 37167 56267 37213
rect 56313 37167 56546 37213
rect 56212 37050 56546 37167
rect 56212 37004 56267 37050
rect 56313 37004 56546 37050
rect 37938 36150 38492 36169
rect 37938 36104 37957 36150
rect 38473 36104 38492 36150
rect 37938 36085 38492 36104
rect 40779 36150 42995 36210
rect 40779 36104 40836 36150
rect 40882 36104 40994 36150
rect 41040 36104 41152 36150
rect 41198 36104 41310 36150
rect 41356 36104 41469 36150
rect 41515 36104 41627 36150
rect 41673 36104 41785 36150
rect 41831 36104 41943 36150
rect 41989 36104 42101 36150
rect 42147 36104 42259 36150
rect 42305 36104 42418 36150
rect 42464 36104 42576 36150
rect 42622 36104 42734 36150
rect 42780 36104 42892 36150
rect 42938 36104 42995 36150
rect 40779 36044 42995 36104
rect 56212 36887 56546 37004
rect 56212 36841 56267 36887
rect 56313 36841 56546 36887
rect 56212 36723 56546 36841
rect 56212 36677 56267 36723
rect 56313 36677 56546 36723
rect 56212 36560 56546 36677
rect 56212 36514 56267 36560
rect 56313 36514 56546 36560
rect 56212 36397 56546 36514
rect 56212 36351 56267 36397
rect 56313 36351 56546 36397
rect 56212 36234 56546 36351
rect 56212 36188 56267 36234
rect 56313 36188 56546 36234
rect 56212 35977 56546 36188
rect 27751 34223 57297 34607
rect 28620 3906 40188 3925
rect 28620 3860 28639 3906
rect 28685 3860 28755 3906
rect 28801 3860 28871 3906
rect 28917 3860 28987 3906
rect 29033 3860 29103 3906
rect 29149 3860 29219 3906
rect 29265 3860 29335 3906
rect 29381 3860 29451 3906
rect 29497 3860 29567 3906
rect 29613 3860 29683 3906
rect 29729 3860 29799 3906
rect 29845 3860 29915 3906
rect 29961 3860 30031 3906
rect 30077 3860 30147 3906
rect 30193 3860 30263 3906
rect 30309 3860 30379 3906
rect 30425 3860 30495 3906
rect 30541 3860 30611 3906
rect 30657 3860 30727 3906
rect 30773 3860 30843 3906
rect 30889 3860 30959 3906
rect 31005 3860 31075 3906
rect 31121 3860 31191 3906
rect 31237 3860 31307 3906
rect 31353 3860 31423 3906
rect 31469 3860 31539 3906
rect 31585 3860 31655 3906
rect 31701 3860 31771 3906
rect 31817 3860 31887 3906
rect 31933 3860 32003 3906
rect 32049 3860 32119 3906
rect 32165 3860 32235 3906
rect 32281 3860 32351 3906
rect 32397 3860 32467 3906
rect 32513 3860 32583 3906
rect 32629 3860 32699 3906
rect 32745 3860 32815 3906
rect 32861 3860 32931 3906
rect 32977 3860 33047 3906
rect 33093 3860 33163 3906
rect 33209 3860 33279 3906
rect 33325 3860 33395 3906
rect 33441 3860 33511 3906
rect 33557 3860 33627 3906
rect 33673 3860 33743 3906
rect 33789 3860 33859 3906
rect 33905 3860 33975 3906
rect 34021 3860 34091 3906
rect 34137 3860 34207 3906
rect 34253 3860 34323 3906
rect 34369 3860 34439 3906
rect 34485 3860 34555 3906
rect 34601 3860 34671 3906
rect 34717 3860 34787 3906
rect 34833 3860 34903 3906
rect 34949 3860 35019 3906
rect 35065 3860 35135 3906
rect 35181 3860 35251 3906
rect 35297 3860 35367 3906
rect 35413 3860 35483 3906
rect 35529 3860 35599 3906
rect 35645 3860 35715 3906
rect 35761 3860 35831 3906
rect 35877 3860 35947 3906
rect 35993 3860 36063 3906
rect 36109 3860 36179 3906
rect 36225 3860 36295 3906
rect 36341 3860 36411 3906
rect 36457 3860 36527 3906
rect 36573 3860 36643 3906
rect 36689 3860 36759 3906
rect 36805 3860 36875 3906
rect 36921 3860 36991 3906
rect 37037 3860 37107 3906
rect 37153 3860 37223 3906
rect 37269 3860 37339 3906
rect 37385 3860 37455 3906
rect 37501 3860 37571 3906
rect 37617 3860 37687 3906
rect 37733 3860 37803 3906
rect 37849 3860 37919 3906
rect 37965 3860 38035 3906
rect 38081 3860 38151 3906
rect 38197 3860 38267 3906
rect 38313 3860 38383 3906
rect 38429 3860 38499 3906
rect 38545 3860 38615 3906
rect 38661 3860 38731 3906
rect 38777 3860 38847 3906
rect 38893 3860 38963 3906
rect 39009 3860 39079 3906
rect 39125 3860 39195 3906
rect 39241 3860 39311 3906
rect 39357 3860 39427 3906
rect 39473 3860 39543 3906
rect 39589 3860 39659 3906
rect 39705 3860 39775 3906
rect 39821 3860 39891 3906
rect 39937 3860 40007 3906
rect 40053 3860 40123 3906
rect 40169 3860 40188 3906
rect 28620 3790 40188 3860
rect 28620 3744 28639 3790
rect 28685 3744 28755 3790
rect 28801 3744 28871 3790
rect 28917 3744 28987 3790
rect 29033 3744 29103 3790
rect 29149 3744 29219 3790
rect 29265 3744 29335 3790
rect 29381 3744 29451 3790
rect 29497 3744 29567 3790
rect 29613 3744 29683 3790
rect 29729 3744 29799 3790
rect 29845 3744 29915 3790
rect 29961 3744 30031 3790
rect 30077 3744 30147 3790
rect 30193 3744 30263 3790
rect 30309 3744 30379 3790
rect 30425 3744 30495 3790
rect 30541 3744 30611 3790
rect 30657 3744 30727 3790
rect 30773 3744 30843 3790
rect 30889 3744 30959 3790
rect 31005 3744 31075 3790
rect 31121 3744 31191 3790
rect 31237 3744 31307 3790
rect 31353 3744 31423 3790
rect 31469 3744 31539 3790
rect 31585 3744 31655 3790
rect 31701 3744 31771 3790
rect 31817 3744 31887 3790
rect 31933 3744 32003 3790
rect 32049 3744 32119 3790
rect 32165 3744 32235 3790
rect 32281 3744 32351 3790
rect 32397 3744 32467 3790
rect 32513 3744 32583 3790
rect 32629 3744 32699 3790
rect 32745 3744 32815 3790
rect 32861 3744 32931 3790
rect 32977 3744 33047 3790
rect 33093 3744 33163 3790
rect 33209 3744 33279 3790
rect 33325 3744 33395 3790
rect 33441 3744 33511 3790
rect 33557 3744 33627 3790
rect 33673 3744 33743 3790
rect 33789 3744 33859 3790
rect 33905 3744 33975 3790
rect 34021 3744 34091 3790
rect 34137 3744 34207 3790
rect 34253 3744 34323 3790
rect 34369 3744 34439 3790
rect 34485 3744 34555 3790
rect 34601 3744 34671 3790
rect 34717 3744 34787 3790
rect 34833 3744 34903 3790
rect 34949 3744 35019 3790
rect 35065 3744 35135 3790
rect 35181 3744 35251 3790
rect 35297 3744 35367 3790
rect 35413 3744 35483 3790
rect 35529 3744 35599 3790
rect 35645 3744 35715 3790
rect 35761 3744 35831 3790
rect 35877 3744 35947 3790
rect 35993 3744 36063 3790
rect 36109 3744 36179 3790
rect 36225 3744 36295 3790
rect 36341 3744 36411 3790
rect 36457 3744 36527 3790
rect 36573 3744 36643 3790
rect 36689 3744 36759 3790
rect 36805 3744 36875 3790
rect 36921 3744 36991 3790
rect 37037 3744 37107 3790
rect 37153 3744 37223 3790
rect 37269 3744 37339 3790
rect 37385 3744 37455 3790
rect 37501 3744 37571 3790
rect 37617 3744 37687 3790
rect 37733 3744 37803 3790
rect 37849 3744 37919 3790
rect 37965 3744 38035 3790
rect 38081 3744 38151 3790
rect 38197 3744 38267 3790
rect 38313 3744 38383 3790
rect 38429 3744 38499 3790
rect 38545 3744 38615 3790
rect 38661 3744 38731 3790
rect 38777 3744 38847 3790
rect 38893 3744 38963 3790
rect 39009 3744 39079 3790
rect 39125 3744 39195 3790
rect 39241 3744 39311 3790
rect 39357 3744 39427 3790
rect 39473 3744 39543 3790
rect 39589 3744 39659 3790
rect 39705 3744 39775 3790
rect 39821 3744 39891 3790
rect 39937 3744 40007 3790
rect 40053 3744 40123 3790
rect 40169 3744 40188 3790
rect 28620 3674 40188 3744
rect 28620 3628 28639 3674
rect 28685 3628 28755 3674
rect 28801 3628 28871 3674
rect 28917 3628 28987 3674
rect 29033 3628 29103 3674
rect 29149 3628 29219 3674
rect 29265 3628 29335 3674
rect 29381 3628 29451 3674
rect 29497 3628 29567 3674
rect 29613 3628 29683 3674
rect 29729 3628 29799 3674
rect 29845 3628 29915 3674
rect 29961 3628 30031 3674
rect 30077 3628 30147 3674
rect 30193 3628 30263 3674
rect 30309 3628 30379 3674
rect 30425 3628 30495 3674
rect 30541 3628 30611 3674
rect 30657 3628 30727 3674
rect 30773 3628 30843 3674
rect 30889 3628 30959 3674
rect 31005 3628 31075 3674
rect 31121 3628 31191 3674
rect 31237 3628 31307 3674
rect 31353 3628 31423 3674
rect 31469 3628 31539 3674
rect 31585 3628 31655 3674
rect 31701 3628 31771 3674
rect 31817 3628 31887 3674
rect 31933 3628 32003 3674
rect 32049 3628 32119 3674
rect 32165 3628 32235 3674
rect 32281 3628 32351 3674
rect 32397 3628 32467 3674
rect 32513 3628 32583 3674
rect 32629 3628 32699 3674
rect 32745 3628 32815 3674
rect 32861 3628 32931 3674
rect 32977 3628 33047 3674
rect 33093 3628 33163 3674
rect 33209 3628 33279 3674
rect 33325 3628 33395 3674
rect 33441 3628 33511 3674
rect 33557 3628 33627 3674
rect 33673 3628 33743 3674
rect 33789 3628 33859 3674
rect 33905 3628 33975 3674
rect 34021 3628 34091 3674
rect 34137 3628 34207 3674
rect 34253 3628 34323 3674
rect 34369 3628 34439 3674
rect 34485 3628 34555 3674
rect 34601 3628 34671 3674
rect 34717 3628 34787 3674
rect 34833 3628 34903 3674
rect 34949 3628 35019 3674
rect 35065 3628 35135 3674
rect 35181 3628 35251 3674
rect 35297 3628 35367 3674
rect 35413 3628 35483 3674
rect 35529 3628 35599 3674
rect 35645 3628 35715 3674
rect 35761 3628 35831 3674
rect 35877 3628 35947 3674
rect 35993 3628 36063 3674
rect 36109 3628 36179 3674
rect 36225 3628 36295 3674
rect 36341 3628 36411 3674
rect 36457 3628 36527 3674
rect 36573 3628 36643 3674
rect 36689 3628 36759 3674
rect 36805 3628 36875 3674
rect 36921 3628 36991 3674
rect 37037 3628 37107 3674
rect 37153 3628 37223 3674
rect 37269 3628 37339 3674
rect 37385 3628 37455 3674
rect 37501 3628 37571 3674
rect 37617 3628 37687 3674
rect 37733 3628 37803 3674
rect 37849 3628 37919 3674
rect 37965 3628 38035 3674
rect 38081 3628 38151 3674
rect 38197 3628 38267 3674
rect 38313 3628 38383 3674
rect 38429 3628 38499 3674
rect 38545 3628 38615 3674
rect 38661 3628 38731 3674
rect 38777 3628 38847 3674
rect 38893 3628 38963 3674
rect 39009 3628 39079 3674
rect 39125 3628 39195 3674
rect 39241 3628 39311 3674
rect 39357 3628 39427 3674
rect 39473 3628 39543 3674
rect 39589 3628 39659 3674
rect 39705 3628 39775 3674
rect 39821 3628 39891 3674
rect 39937 3628 40007 3674
rect 40053 3628 40123 3674
rect 40169 3628 40188 3674
rect 28620 3558 40188 3628
rect 28620 3512 28639 3558
rect 28685 3512 28755 3558
rect 28801 3512 28871 3558
rect 28917 3512 28987 3558
rect 29033 3512 29103 3558
rect 29149 3512 29219 3558
rect 29265 3512 29335 3558
rect 29381 3512 29451 3558
rect 29497 3512 29567 3558
rect 29613 3512 29683 3558
rect 29729 3512 29799 3558
rect 29845 3512 29915 3558
rect 29961 3512 30031 3558
rect 30077 3512 30147 3558
rect 30193 3512 30263 3558
rect 30309 3512 30379 3558
rect 30425 3512 30495 3558
rect 30541 3512 30611 3558
rect 30657 3512 30727 3558
rect 30773 3512 30843 3558
rect 30889 3512 30959 3558
rect 31005 3512 31075 3558
rect 31121 3512 31191 3558
rect 31237 3512 31307 3558
rect 31353 3512 31423 3558
rect 31469 3512 31539 3558
rect 31585 3512 31655 3558
rect 31701 3512 31771 3558
rect 31817 3512 31887 3558
rect 31933 3512 32003 3558
rect 32049 3512 32119 3558
rect 32165 3512 32235 3558
rect 32281 3512 32351 3558
rect 32397 3512 32467 3558
rect 32513 3512 32583 3558
rect 32629 3512 32699 3558
rect 32745 3512 32815 3558
rect 32861 3512 32931 3558
rect 32977 3512 33047 3558
rect 33093 3512 33163 3558
rect 33209 3512 33279 3558
rect 33325 3512 33395 3558
rect 33441 3512 33511 3558
rect 33557 3512 33627 3558
rect 33673 3512 33743 3558
rect 33789 3512 33859 3558
rect 33905 3512 33975 3558
rect 34021 3512 34091 3558
rect 34137 3512 34207 3558
rect 34253 3512 34323 3558
rect 34369 3512 34439 3558
rect 34485 3512 34555 3558
rect 34601 3512 34671 3558
rect 34717 3512 34787 3558
rect 34833 3512 34903 3558
rect 34949 3512 35019 3558
rect 35065 3512 35135 3558
rect 35181 3512 35251 3558
rect 35297 3512 35367 3558
rect 35413 3512 35483 3558
rect 35529 3512 35599 3558
rect 35645 3512 35715 3558
rect 35761 3512 35831 3558
rect 35877 3512 35947 3558
rect 35993 3512 36063 3558
rect 36109 3512 36179 3558
rect 36225 3512 36295 3558
rect 36341 3512 36411 3558
rect 36457 3512 36527 3558
rect 36573 3512 36643 3558
rect 36689 3512 36759 3558
rect 36805 3512 36875 3558
rect 36921 3512 36991 3558
rect 37037 3512 37107 3558
rect 37153 3512 37223 3558
rect 37269 3512 37339 3558
rect 37385 3512 37455 3558
rect 37501 3512 37571 3558
rect 37617 3512 37687 3558
rect 37733 3512 37803 3558
rect 37849 3512 37919 3558
rect 37965 3512 38035 3558
rect 38081 3512 38151 3558
rect 38197 3512 38267 3558
rect 38313 3512 38383 3558
rect 38429 3512 38499 3558
rect 38545 3512 38615 3558
rect 38661 3512 38731 3558
rect 38777 3512 38847 3558
rect 38893 3512 38963 3558
rect 39009 3512 39079 3558
rect 39125 3512 39195 3558
rect 39241 3512 39311 3558
rect 39357 3512 39427 3558
rect 39473 3512 39543 3558
rect 39589 3512 39659 3558
rect 39705 3512 39775 3558
rect 39821 3512 39891 3558
rect 39937 3512 40007 3558
rect 40053 3512 40123 3558
rect 40169 3512 40188 3558
rect 28620 3442 40188 3512
rect 28620 3396 28639 3442
rect 28685 3396 28755 3442
rect 28801 3396 28871 3442
rect 28917 3396 28987 3442
rect 29033 3396 29103 3442
rect 29149 3396 29219 3442
rect 29265 3396 29335 3442
rect 29381 3396 29451 3442
rect 29497 3396 29567 3442
rect 29613 3396 29683 3442
rect 29729 3396 29799 3442
rect 29845 3396 29915 3442
rect 29961 3396 30031 3442
rect 30077 3396 30147 3442
rect 30193 3396 30263 3442
rect 30309 3396 30379 3442
rect 30425 3396 30495 3442
rect 30541 3396 30611 3442
rect 30657 3396 30727 3442
rect 30773 3396 30843 3442
rect 30889 3396 30959 3442
rect 31005 3396 31075 3442
rect 31121 3396 31191 3442
rect 31237 3396 31307 3442
rect 31353 3396 31423 3442
rect 31469 3396 31539 3442
rect 31585 3396 31655 3442
rect 31701 3396 31771 3442
rect 31817 3396 31887 3442
rect 31933 3396 32003 3442
rect 32049 3396 32119 3442
rect 32165 3396 32235 3442
rect 32281 3396 32351 3442
rect 32397 3396 32467 3442
rect 32513 3396 32583 3442
rect 32629 3396 32699 3442
rect 32745 3396 32815 3442
rect 32861 3396 32931 3442
rect 32977 3396 33047 3442
rect 33093 3396 33163 3442
rect 33209 3396 33279 3442
rect 33325 3396 33395 3442
rect 33441 3396 33511 3442
rect 33557 3396 33627 3442
rect 33673 3396 33743 3442
rect 33789 3396 33859 3442
rect 33905 3396 33975 3442
rect 34021 3396 34091 3442
rect 34137 3396 34207 3442
rect 34253 3396 34323 3442
rect 34369 3396 34439 3442
rect 34485 3396 34555 3442
rect 34601 3396 34671 3442
rect 34717 3396 34787 3442
rect 34833 3396 34903 3442
rect 34949 3396 35019 3442
rect 35065 3396 35135 3442
rect 35181 3396 35251 3442
rect 35297 3396 35367 3442
rect 35413 3396 35483 3442
rect 35529 3396 35599 3442
rect 35645 3396 35715 3442
rect 35761 3396 35831 3442
rect 35877 3396 35947 3442
rect 35993 3396 36063 3442
rect 36109 3396 36179 3442
rect 36225 3396 36295 3442
rect 36341 3396 36411 3442
rect 36457 3396 36527 3442
rect 36573 3396 36643 3442
rect 36689 3396 36759 3442
rect 36805 3396 36875 3442
rect 36921 3396 36991 3442
rect 37037 3396 37107 3442
rect 37153 3396 37223 3442
rect 37269 3396 37339 3442
rect 37385 3396 37455 3442
rect 37501 3396 37571 3442
rect 37617 3396 37687 3442
rect 37733 3396 37803 3442
rect 37849 3396 37919 3442
rect 37965 3396 38035 3442
rect 38081 3396 38151 3442
rect 38197 3396 38267 3442
rect 38313 3396 38383 3442
rect 38429 3396 38499 3442
rect 38545 3396 38615 3442
rect 38661 3396 38731 3442
rect 38777 3396 38847 3442
rect 38893 3396 38963 3442
rect 39009 3396 39079 3442
rect 39125 3396 39195 3442
rect 39241 3396 39311 3442
rect 39357 3396 39427 3442
rect 39473 3396 39543 3442
rect 39589 3396 39659 3442
rect 39705 3396 39775 3442
rect 39821 3396 39891 3442
rect 39937 3396 40007 3442
rect 40053 3396 40123 3442
rect 40169 3396 40188 3442
rect 28620 3326 40188 3396
rect 28620 3280 28639 3326
rect 28685 3280 28755 3326
rect 28801 3280 28871 3326
rect 28917 3280 28987 3326
rect 29033 3280 29103 3326
rect 29149 3280 29219 3326
rect 29265 3280 29335 3326
rect 29381 3280 29451 3326
rect 29497 3280 29567 3326
rect 29613 3280 29683 3326
rect 29729 3280 29799 3326
rect 29845 3280 29915 3326
rect 29961 3280 30031 3326
rect 30077 3280 30147 3326
rect 30193 3280 30263 3326
rect 30309 3280 30379 3326
rect 30425 3280 30495 3326
rect 30541 3280 30611 3326
rect 30657 3280 30727 3326
rect 30773 3280 30843 3326
rect 30889 3280 30959 3326
rect 31005 3280 31075 3326
rect 31121 3280 31191 3326
rect 31237 3280 31307 3326
rect 31353 3280 31423 3326
rect 31469 3280 31539 3326
rect 31585 3280 31655 3326
rect 31701 3280 31771 3326
rect 31817 3280 31887 3326
rect 31933 3280 32003 3326
rect 32049 3280 32119 3326
rect 32165 3280 32235 3326
rect 32281 3280 32351 3326
rect 32397 3280 32467 3326
rect 32513 3280 32583 3326
rect 32629 3280 32699 3326
rect 32745 3280 32815 3326
rect 32861 3280 32931 3326
rect 32977 3280 33047 3326
rect 33093 3280 33163 3326
rect 33209 3280 33279 3326
rect 33325 3280 33395 3326
rect 33441 3280 33511 3326
rect 33557 3280 33627 3326
rect 33673 3280 33743 3326
rect 33789 3280 33859 3326
rect 33905 3280 33975 3326
rect 34021 3280 34091 3326
rect 34137 3280 34207 3326
rect 34253 3280 34323 3326
rect 34369 3280 34439 3326
rect 34485 3280 34555 3326
rect 34601 3280 34671 3326
rect 34717 3280 34787 3326
rect 34833 3280 34903 3326
rect 34949 3280 35019 3326
rect 35065 3280 35135 3326
rect 35181 3280 35251 3326
rect 35297 3280 35367 3326
rect 35413 3280 35483 3326
rect 35529 3280 35599 3326
rect 35645 3280 35715 3326
rect 35761 3280 35831 3326
rect 35877 3280 35947 3326
rect 35993 3280 36063 3326
rect 36109 3280 36179 3326
rect 36225 3280 36295 3326
rect 36341 3280 36411 3326
rect 36457 3280 36527 3326
rect 36573 3280 36643 3326
rect 36689 3280 36759 3326
rect 36805 3280 36875 3326
rect 36921 3280 36991 3326
rect 37037 3280 37107 3326
rect 37153 3280 37223 3326
rect 37269 3280 37339 3326
rect 37385 3280 37455 3326
rect 37501 3280 37571 3326
rect 37617 3280 37687 3326
rect 37733 3280 37803 3326
rect 37849 3280 37919 3326
rect 37965 3280 38035 3326
rect 38081 3280 38151 3326
rect 38197 3280 38267 3326
rect 38313 3280 38383 3326
rect 38429 3280 38499 3326
rect 38545 3280 38615 3326
rect 38661 3280 38731 3326
rect 38777 3280 38847 3326
rect 38893 3280 38963 3326
rect 39009 3280 39079 3326
rect 39125 3280 39195 3326
rect 39241 3280 39311 3326
rect 39357 3280 39427 3326
rect 39473 3280 39543 3326
rect 39589 3280 39659 3326
rect 39705 3280 39775 3326
rect 39821 3280 39891 3326
rect 39937 3280 40007 3326
rect 40053 3280 40123 3326
rect 40169 3280 40188 3326
rect 28620 3210 40188 3280
rect 28620 3164 28639 3210
rect 28685 3164 28755 3210
rect 28801 3164 28871 3210
rect 28917 3164 28987 3210
rect 29033 3164 29103 3210
rect 29149 3164 29219 3210
rect 29265 3164 29335 3210
rect 29381 3164 29451 3210
rect 29497 3164 29567 3210
rect 29613 3164 29683 3210
rect 29729 3164 29799 3210
rect 29845 3164 29915 3210
rect 29961 3164 30031 3210
rect 30077 3164 30147 3210
rect 30193 3164 30263 3210
rect 30309 3164 30379 3210
rect 30425 3164 30495 3210
rect 30541 3164 30611 3210
rect 30657 3164 30727 3210
rect 30773 3164 30843 3210
rect 30889 3164 30959 3210
rect 31005 3164 31075 3210
rect 31121 3164 31191 3210
rect 31237 3164 31307 3210
rect 31353 3164 31423 3210
rect 31469 3164 31539 3210
rect 31585 3164 31655 3210
rect 31701 3164 31771 3210
rect 31817 3164 31887 3210
rect 31933 3164 32003 3210
rect 32049 3164 32119 3210
rect 32165 3164 32235 3210
rect 32281 3164 32351 3210
rect 32397 3164 32467 3210
rect 32513 3164 32583 3210
rect 32629 3164 32699 3210
rect 32745 3164 32815 3210
rect 32861 3164 32931 3210
rect 32977 3164 33047 3210
rect 33093 3164 33163 3210
rect 33209 3164 33279 3210
rect 33325 3164 33395 3210
rect 33441 3164 33511 3210
rect 33557 3164 33627 3210
rect 33673 3164 33743 3210
rect 33789 3164 33859 3210
rect 33905 3164 33975 3210
rect 34021 3164 34091 3210
rect 34137 3164 34207 3210
rect 34253 3164 34323 3210
rect 34369 3164 34439 3210
rect 34485 3164 34555 3210
rect 34601 3164 34671 3210
rect 34717 3164 34787 3210
rect 34833 3164 34903 3210
rect 34949 3164 35019 3210
rect 35065 3164 35135 3210
rect 35181 3164 35251 3210
rect 35297 3164 35367 3210
rect 35413 3164 35483 3210
rect 35529 3164 35599 3210
rect 35645 3164 35715 3210
rect 35761 3164 35831 3210
rect 35877 3164 35947 3210
rect 35993 3164 36063 3210
rect 36109 3164 36179 3210
rect 36225 3164 36295 3210
rect 36341 3164 36411 3210
rect 36457 3164 36527 3210
rect 36573 3164 36643 3210
rect 36689 3164 36759 3210
rect 36805 3164 36875 3210
rect 36921 3164 36991 3210
rect 37037 3164 37107 3210
rect 37153 3164 37223 3210
rect 37269 3164 37339 3210
rect 37385 3164 37455 3210
rect 37501 3164 37571 3210
rect 37617 3164 37687 3210
rect 37733 3164 37803 3210
rect 37849 3164 37919 3210
rect 37965 3164 38035 3210
rect 38081 3164 38151 3210
rect 38197 3164 38267 3210
rect 38313 3164 38383 3210
rect 38429 3164 38499 3210
rect 38545 3164 38615 3210
rect 38661 3164 38731 3210
rect 38777 3164 38847 3210
rect 38893 3164 38963 3210
rect 39009 3164 39079 3210
rect 39125 3164 39195 3210
rect 39241 3164 39311 3210
rect 39357 3164 39427 3210
rect 39473 3164 39543 3210
rect 39589 3164 39659 3210
rect 39705 3164 39775 3210
rect 39821 3164 39891 3210
rect 39937 3164 40007 3210
rect 40053 3164 40123 3210
rect 40169 3164 40188 3210
rect 28620 3094 40188 3164
rect 28620 3048 28639 3094
rect 28685 3048 28755 3094
rect 28801 3048 28871 3094
rect 28917 3048 28987 3094
rect 29033 3048 29103 3094
rect 29149 3048 29219 3094
rect 29265 3048 29335 3094
rect 29381 3048 29451 3094
rect 29497 3048 29567 3094
rect 29613 3048 29683 3094
rect 29729 3048 29799 3094
rect 29845 3048 29915 3094
rect 29961 3048 30031 3094
rect 30077 3048 30147 3094
rect 30193 3048 30263 3094
rect 30309 3048 30379 3094
rect 30425 3048 30495 3094
rect 30541 3048 30611 3094
rect 30657 3048 30727 3094
rect 30773 3048 30843 3094
rect 30889 3048 30959 3094
rect 31005 3048 31075 3094
rect 31121 3048 31191 3094
rect 31237 3048 31307 3094
rect 31353 3048 31423 3094
rect 31469 3048 31539 3094
rect 31585 3048 31655 3094
rect 31701 3048 31771 3094
rect 31817 3048 31887 3094
rect 31933 3048 32003 3094
rect 32049 3048 32119 3094
rect 32165 3048 32235 3094
rect 32281 3048 32351 3094
rect 32397 3048 32467 3094
rect 32513 3048 32583 3094
rect 32629 3048 32699 3094
rect 32745 3048 32815 3094
rect 32861 3048 32931 3094
rect 32977 3048 33047 3094
rect 33093 3048 33163 3094
rect 33209 3048 33279 3094
rect 33325 3048 33395 3094
rect 33441 3048 33511 3094
rect 33557 3048 33627 3094
rect 33673 3048 33743 3094
rect 33789 3048 33859 3094
rect 33905 3048 33975 3094
rect 34021 3048 34091 3094
rect 34137 3048 34207 3094
rect 34253 3048 34323 3094
rect 34369 3048 34439 3094
rect 34485 3048 34555 3094
rect 34601 3048 34671 3094
rect 34717 3048 34787 3094
rect 34833 3048 34903 3094
rect 34949 3048 35019 3094
rect 35065 3048 35135 3094
rect 35181 3048 35251 3094
rect 35297 3048 35367 3094
rect 35413 3048 35483 3094
rect 35529 3048 35599 3094
rect 35645 3048 35715 3094
rect 35761 3048 35831 3094
rect 35877 3048 35947 3094
rect 35993 3048 36063 3094
rect 36109 3048 36179 3094
rect 36225 3048 36295 3094
rect 36341 3048 36411 3094
rect 36457 3048 36527 3094
rect 36573 3048 36643 3094
rect 36689 3048 36759 3094
rect 36805 3048 36875 3094
rect 36921 3048 36991 3094
rect 37037 3048 37107 3094
rect 37153 3048 37223 3094
rect 37269 3048 37339 3094
rect 37385 3048 37455 3094
rect 37501 3048 37571 3094
rect 37617 3048 37687 3094
rect 37733 3048 37803 3094
rect 37849 3048 37919 3094
rect 37965 3048 38035 3094
rect 38081 3048 38151 3094
rect 38197 3048 38267 3094
rect 38313 3048 38383 3094
rect 38429 3048 38499 3094
rect 38545 3048 38615 3094
rect 38661 3048 38731 3094
rect 38777 3048 38847 3094
rect 38893 3048 38963 3094
rect 39009 3048 39079 3094
rect 39125 3048 39195 3094
rect 39241 3048 39311 3094
rect 39357 3048 39427 3094
rect 39473 3048 39543 3094
rect 39589 3048 39659 3094
rect 39705 3048 39775 3094
rect 39821 3048 39891 3094
rect 39937 3048 40007 3094
rect 40053 3048 40123 3094
rect 40169 3048 40188 3094
rect 28620 2978 40188 3048
rect 28620 2932 28639 2978
rect 28685 2932 28755 2978
rect 28801 2932 28871 2978
rect 28917 2932 28987 2978
rect 29033 2932 29103 2978
rect 29149 2932 29219 2978
rect 29265 2932 29335 2978
rect 29381 2932 29451 2978
rect 29497 2932 29567 2978
rect 29613 2932 29683 2978
rect 29729 2932 29799 2978
rect 29845 2932 29915 2978
rect 29961 2932 30031 2978
rect 30077 2932 30147 2978
rect 30193 2932 30263 2978
rect 30309 2932 30379 2978
rect 30425 2932 30495 2978
rect 30541 2932 30611 2978
rect 30657 2932 30727 2978
rect 30773 2932 30843 2978
rect 30889 2932 30959 2978
rect 31005 2932 31075 2978
rect 31121 2932 31191 2978
rect 31237 2932 31307 2978
rect 31353 2932 31423 2978
rect 31469 2932 31539 2978
rect 31585 2932 31655 2978
rect 31701 2932 31771 2978
rect 31817 2932 31887 2978
rect 31933 2932 32003 2978
rect 32049 2932 32119 2978
rect 32165 2932 32235 2978
rect 32281 2932 32351 2978
rect 32397 2932 32467 2978
rect 32513 2932 32583 2978
rect 32629 2932 32699 2978
rect 32745 2932 32815 2978
rect 32861 2932 32931 2978
rect 32977 2932 33047 2978
rect 33093 2932 33163 2978
rect 33209 2932 33279 2978
rect 33325 2932 33395 2978
rect 33441 2932 33511 2978
rect 33557 2932 33627 2978
rect 33673 2932 33743 2978
rect 33789 2932 33859 2978
rect 33905 2932 33975 2978
rect 34021 2932 34091 2978
rect 34137 2932 34207 2978
rect 34253 2932 34323 2978
rect 34369 2932 34439 2978
rect 34485 2932 34555 2978
rect 34601 2932 34671 2978
rect 34717 2932 34787 2978
rect 34833 2932 34903 2978
rect 34949 2932 35019 2978
rect 35065 2932 35135 2978
rect 35181 2932 35251 2978
rect 35297 2932 35367 2978
rect 35413 2932 35483 2978
rect 35529 2932 35599 2978
rect 35645 2932 35715 2978
rect 35761 2932 35831 2978
rect 35877 2932 35947 2978
rect 35993 2932 36063 2978
rect 36109 2932 36179 2978
rect 36225 2932 36295 2978
rect 36341 2932 36411 2978
rect 36457 2932 36527 2978
rect 36573 2932 36643 2978
rect 36689 2932 36759 2978
rect 36805 2932 36875 2978
rect 36921 2932 36991 2978
rect 37037 2932 37107 2978
rect 37153 2932 37223 2978
rect 37269 2932 37339 2978
rect 37385 2932 37455 2978
rect 37501 2932 37571 2978
rect 37617 2932 37687 2978
rect 37733 2932 37803 2978
rect 37849 2932 37919 2978
rect 37965 2932 38035 2978
rect 38081 2932 38151 2978
rect 38197 2932 38267 2978
rect 38313 2932 38383 2978
rect 38429 2932 38499 2978
rect 38545 2932 38615 2978
rect 38661 2932 38731 2978
rect 38777 2932 38847 2978
rect 38893 2932 38963 2978
rect 39009 2932 39079 2978
rect 39125 2932 39195 2978
rect 39241 2932 39311 2978
rect 39357 2932 39427 2978
rect 39473 2932 39543 2978
rect 39589 2932 39659 2978
rect 39705 2932 39775 2978
rect 39821 2932 39891 2978
rect 39937 2932 40007 2978
rect 40053 2932 40123 2978
rect 40169 2932 40188 2978
rect 28620 2862 40188 2932
rect 28620 2816 28639 2862
rect 28685 2816 28755 2862
rect 28801 2816 28871 2862
rect 28917 2816 28987 2862
rect 29033 2816 29103 2862
rect 29149 2816 29219 2862
rect 29265 2816 29335 2862
rect 29381 2816 29451 2862
rect 29497 2816 29567 2862
rect 29613 2816 29683 2862
rect 29729 2816 29799 2862
rect 29845 2816 29915 2862
rect 29961 2816 30031 2862
rect 30077 2816 30147 2862
rect 30193 2816 30263 2862
rect 30309 2816 30379 2862
rect 30425 2816 30495 2862
rect 30541 2816 30611 2862
rect 30657 2816 30727 2862
rect 30773 2816 30843 2862
rect 30889 2816 30959 2862
rect 31005 2816 31075 2862
rect 31121 2816 31191 2862
rect 31237 2816 31307 2862
rect 31353 2816 31423 2862
rect 31469 2816 31539 2862
rect 31585 2816 31655 2862
rect 31701 2816 31771 2862
rect 31817 2816 31887 2862
rect 31933 2816 32003 2862
rect 32049 2816 32119 2862
rect 32165 2816 32235 2862
rect 32281 2816 32351 2862
rect 32397 2816 32467 2862
rect 32513 2816 32583 2862
rect 32629 2816 32699 2862
rect 32745 2816 32815 2862
rect 32861 2816 32931 2862
rect 32977 2816 33047 2862
rect 33093 2816 33163 2862
rect 33209 2816 33279 2862
rect 33325 2816 33395 2862
rect 33441 2816 33511 2862
rect 33557 2816 33627 2862
rect 33673 2816 33743 2862
rect 33789 2816 33859 2862
rect 33905 2816 33975 2862
rect 34021 2816 34091 2862
rect 34137 2816 34207 2862
rect 34253 2816 34323 2862
rect 34369 2816 34439 2862
rect 34485 2816 34555 2862
rect 34601 2816 34671 2862
rect 34717 2816 34787 2862
rect 34833 2816 34903 2862
rect 34949 2816 35019 2862
rect 35065 2816 35135 2862
rect 35181 2816 35251 2862
rect 35297 2816 35367 2862
rect 35413 2816 35483 2862
rect 35529 2816 35599 2862
rect 35645 2816 35715 2862
rect 35761 2816 35831 2862
rect 35877 2816 35947 2862
rect 35993 2816 36063 2862
rect 36109 2816 36179 2862
rect 36225 2816 36295 2862
rect 36341 2816 36411 2862
rect 36457 2816 36527 2862
rect 36573 2816 36643 2862
rect 36689 2816 36759 2862
rect 36805 2816 36875 2862
rect 36921 2816 36991 2862
rect 37037 2816 37107 2862
rect 37153 2816 37223 2862
rect 37269 2816 37339 2862
rect 37385 2816 37455 2862
rect 37501 2816 37571 2862
rect 37617 2816 37687 2862
rect 37733 2816 37803 2862
rect 37849 2816 37919 2862
rect 37965 2816 38035 2862
rect 38081 2816 38151 2862
rect 38197 2816 38267 2862
rect 38313 2816 38383 2862
rect 38429 2816 38499 2862
rect 38545 2816 38615 2862
rect 38661 2816 38731 2862
rect 38777 2816 38847 2862
rect 38893 2816 38963 2862
rect 39009 2816 39079 2862
rect 39125 2816 39195 2862
rect 39241 2816 39311 2862
rect 39357 2816 39427 2862
rect 39473 2816 39543 2862
rect 39589 2816 39659 2862
rect 39705 2816 39775 2862
rect 39821 2816 39891 2862
rect 39937 2816 40007 2862
rect 40053 2816 40123 2862
rect 40169 2816 40188 2862
rect 28620 2746 40188 2816
rect 28620 2700 28639 2746
rect 28685 2700 28755 2746
rect 28801 2700 28871 2746
rect 28917 2700 28987 2746
rect 29033 2700 29103 2746
rect 29149 2700 29219 2746
rect 29265 2700 29335 2746
rect 29381 2700 29451 2746
rect 29497 2700 29567 2746
rect 29613 2700 29683 2746
rect 29729 2700 29799 2746
rect 29845 2700 29915 2746
rect 29961 2700 30031 2746
rect 30077 2700 30147 2746
rect 30193 2700 30263 2746
rect 30309 2700 30379 2746
rect 30425 2700 30495 2746
rect 30541 2700 30611 2746
rect 30657 2700 30727 2746
rect 30773 2700 30843 2746
rect 30889 2700 30959 2746
rect 31005 2700 31075 2746
rect 31121 2700 31191 2746
rect 31237 2700 31307 2746
rect 31353 2700 31423 2746
rect 31469 2700 31539 2746
rect 31585 2700 31655 2746
rect 31701 2700 31771 2746
rect 31817 2700 31887 2746
rect 31933 2700 32003 2746
rect 32049 2700 32119 2746
rect 32165 2700 32235 2746
rect 32281 2700 32351 2746
rect 32397 2700 32467 2746
rect 32513 2700 32583 2746
rect 32629 2700 32699 2746
rect 32745 2700 32815 2746
rect 32861 2700 32931 2746
rect 32977 2700 33047 2746
rect 33093 2700 33163 2746
rect 33209 2700 33279 2746
rect 33325 2700 33395 2746
rect 33441 2700 33511 2746
rect 33557 2700 33627 2746
rect 33673 2700 33743 2746
rect 33789 2700 33859 2746
rect 33905 2700 33975 2746
rect 34021 2700 34091 2746
rect 34137 2700 34207 2746
rect 34253 2700 34323 2746
rect 34369 2700 34439 2746
rect 34485 2700 34555 2746
rect 34601 2700 34671 2746
rect 34717 2700 34787 2746
rect 34833 2700 34903 2746
rect 34949 2700 35019 2746
rect 35065 2700 35135 2746
rect 35181 2700 35251 2746
rect 35297 2700 35367 2746
rect 35413 2700 35483 2746
rect 35529 2700 35599 2746
rect 35645 2700 35715 2746
rect 35761 2700 35831 2746
rect 35877 2700 35947 2746
rect 35993 2700 36063 2746
rect 36109 2700 36179 2746
rect 36225 2700 36295 2746
rect 36341 2700 36411 2746
rect 36457 2700 36527 2746
rect 36573 2700 36643 2746
rect 36689 2700 36759 2746
rect 36805 2700 36875 2746
rect 36921 2700 36991 2746
rect 37037 2700 37107 2746
rect 37153 2700 37223 2746
rect 37269 2700 37339 2746
rect 37385 2700 37455 2746
rect 37501 2700 37571 2746
rect 37617 2700 37687 2746
rect 37733 2700 37803 2746
rect 37849 2700 37919 2746
rect 37965 2700 38035 2746
rect 38081 2700 38151 2746
rect 38197 2700 38267 2746
rect 38313 2700 38383 2746
rect 38429 2700 38499 2746
rect 38545 2700 38615 2746
rect 38661 2700 38731 2746
rect 38777 2700 38847 2746
rect 38893 2700 38963 2746
rect 39009 2700 39079 2746
rect 39125 2700 39195 2746
rect 39241 2700 39311 2746
rect 39357 2700 39427 2746
rect 39473 2700 39543 2746
rect 39589 2700 39659 2746
rect 39705 2700 39775 2746
rect 39821 2700 39891 2746
rect 39937 2700 40007 2746
rect 40053 2700 40123 2746
rect 40169 2700 40188 2746
rect 28620 2630 40188 2700
rect 28620 2584 28639 2630
rect 28685 2584 28755 2630
rect 28801 2584 28871 2630
rect 28917 2584 28987 2630
rect 29033 2584 29103 2630
rect 29149 2584 29219 2630
rect 29265 2584 29335 2630
rect 29381 2584 29451 2630
rect 29497 2584 29567 2630
rect 29613 2584 29683 2630
rect 29729 2584 29799 2630
rect 29845 2584 29915 2630
rect 29961 2584 30031 2630
rect 30077 2584 30147 2630
rect 30193 2584 30263 2630
rect 30309 2584 30379 2630
rect 30425 2584 30495 2630
rect 30541 2584 30611 2630
rect 30657 2584 30727 2630
rect 30773 2584 30843 2630
rect 30889 2584 30959 2630
rect 31005 2584 31075 2630
rect 31121 2584 31191 2630
rect 31237 2584 31307 2630
rect 31353 2584 31423 2630
rect 31469 2584 31539 2630
rect 31585 2584 31655 2630
rect 31701 2584 31771 2630
rect 31817 2584 31887 2630
rect 31933 2584 32003 2630
rect 32049 2584 32119 2630
rect 32165 2584 32235 2630
rect 32281 2584 32351 2630
rect 32397 2584 32467 2630
rect 32513 2584 32583 2630
rect 32629 2584 32699 2630
rect 32745 2584 32815 2630
rect 32861 2584 32931 2630
rect 32977 2584 33047 2630
rect 33093 2584 33163 2630
rect 33209 2584 33279 2630
rect 33325 2584 33395 2630
rect 33441 2584 33511 2630
rect 33557 2584 33627 2630
rect 33673 2584 33743 2630
rect 33789 2584 33859 2630
rect 33905 2584 33975 2630
rect 34021 2584 34091 2630
rect 34137 2584 34207 2630
rect 34253 2584 34323 2630
rect 34369 2584 34439 2630
rect 34485 2584 34555 2630
rect 34601 2584 34671 2630
rect 34717 2584 34787 2630
rect 34833 2584 34903 2630
rect 34949 2584 35019 2630
rect 35065 2584 35135 2630
rect 35181 2584 35251 2630
rect 35297 2584 35367 2630
rect 35413 2584 35483 2630
rect 35529 2584 35599 2630
rect 35645 2584 35715 2630
rect 35761 2584 35831 2630
rect 35877 2584 35947 2630
rect 35993 2584 36063 2630
rect 36109 2584 36179 2630
rect 36225 2584 36295 2630
rect 36341 2584 36411 2630
rect 36457 2584 36527 2630
rect 36573 2584 36643 2630
rect 36689 2584 36759 2630
rect 36805 2584 36875 2630
rect 36921 2584 36991 2630
rect 37037 2584 37107 2630
rect 37153 2584 37223 2630
rect 37269 2584 37339 2630
rect 37385 2584 37455 2630
rect 37501 2584 37571 2630
rect 37617 2584 37687 2630
rect 37733 2584 37803 2630
rect 37849 2584 37919 2630
rect 37965 2584 38035 2630
rect 38081 2584 38151 2630
rect 38197 2584 38267 2630
rect 38313 2584 38383 2630
rect 38429 2584 38499 2630
rect 38545 2584 38615 2630
rect 38661 2584 38731 2630
rect 38777 2584 38847 2630
rect 38893 2584 38963 2630
rect 39009 2584 39079 2630
rect 39125 2584 39195 2630
rect 39241 2584 39311 2630
rect 39357 2584 39427 2630
rect 39473 2584 39543 2630
rect 39589 2584 39659 2630
rect 39705 2584 39775 2630
rect 39821 2584 39891 2630
rect 39937 2584 40007 2630
rect 40053 2584 40123 2630
rect 40169 2584 40188 2630
rect 28620 2514 40188 2584
rect 28620 2468 28639 2514
rect 28685 2468 28755 2514
rect 28801 2468 28871 2514
rect 28917 2468 28987 2514
rect 29033 2468 29103 2514
rect 29149 2468 29219 2514
rect 29265 2468 29335 2514
rect 29381 2468 29451 2514
rect 29497 2468 29567 2514
rect 29613 2468 29683 2514
rect 29729 2468 29799 2514
rect 29845 2468 29915 2514
rect 29961 2468 30031 2514
rect 30077 2468 30147 2514
rect 30193 2468 30263 2514
rect 30309 2468 30379 2514
rect 30425 2468 30495 2514
rect 30541 2468 30611 2514
rect 30657 2468 30727 2514
rect 30773 2468 30843 2514
rect 30889 2468 30959 2514
rect 31005 2468 31075 2514
rect 31121 2468 31191 2514
rect 31237 2468 31307 2514
rect 31353 2468 31423 2514
rect 31469 2468 31539 2514
rect 31585 2468 31655 2514
rect 31701 2468 31771 2514
rect 31817 2468 31887 2514
rect 31933 2468 32003 2514
rect 32049 2468 32119 2514
rect 32165 2468 32235 2514
rect 32281 2468 32351 2514
rect 32397 2468 32467 2514
rect 32513 2468 32583 2514
rect 32629 2468 32699 2514
rect 32745 2468 32815 2514
rect 32861 2468 32931 2514
rect 32977 2468 33047 2514
rect 33093 2468 33163 2514
rect 33209 2468 33279 2514
rect 33325 2468 33395 2514
rect 33441 2468 33511 2514
rect 33557 2468 33627 2514
rect 33673 2468 33743 2514
rect 33789 2468 33859 2514
rect 33905 2468 33975 2514
rect 34021 2468 34091 2514
rect 34137 2468 34207 2514
rect 34253 2468 34323 2514
rect 34369 2468 34439 2514
rect 34485 2468 34555 2514
rect 34601 2468 34671 2514
rect 34717 2468 34787 2514
rect 34833 2468 34903 2514
rect 34949 2468 35019 2514
rect 35065 2468 35135 2514
rect 35181 2468 35251 2514
rect 35297 2468 35367 2514
rect 35413 2468 35483 2514
rect 35529 2468 35599 2514
rect 35645 2468 35715 2514
rect 35761 2468 35831 2514
rect 35877 2468 35947 2514
rect 35993 2468 36063 2514
rect 36109 2468 36179 2514
rect 36225 2468 36295 2514
rect 36341 2468 36411 2514
rect 36457 2468 36527 2514
rect 36573 2468 36643 2514
rect 36689 2468 36759 2514
rect 36805 2468 36875 2514
rect 36921 2468 36991 2514
rect 37037 2468 37107 2514
rect 37153 2468 37223 2514
rect 37269 2468 37339 2514
rect 37385 2468 37455 2514
rect 37501 2468 37571 2514
rect 37617 2468 37687 2514
rect 37733 2468 37803 2514
rect 37849 2468 37919 2514
rect 37965 2468 38035 2514
rect 38081 2468 38151 2514
rect 38197 2468 38267 2514
rect 38313 2468 38383 2514
rect 38429 2468 38499 2514
rect 38545 2468 38615 2514
rect 38661 2468 38731 2514
rect 38777 2468 38847 2514
rect 38893 2468 38963 2514
rect 39009 2468 39079 2514
rect 39125 2468 39195 2514
rect 39241 2468 39311 2514
rect 39357 2468 39427 2514
rect 39473 2468 39543 2514
rect 39589 2468 39659 2514
rect 39705 2468 39775 2514
rect 39821 2468 39891 2514
rect 39937 2468 40007 2514
rect 40053 2468 40123 2514
rect 40169 2468 40188 2514
rect 28620 2398 40188 2468
rect 28620 2352 28639 2398
rect 28685 2352 28755 2398
rect 28801 2352 28871 2398
rect 28917 2352 28987 2398
rect 29033 2352 29103 2398
rect 29149 2352 29219 2398
rect 29265 2352 29335 2398
rect 29381 2352 29451 2398
rect 29497 2352 29567 2398
rect 29613 2352 29683 2398
rect 29729 2352 29799 2398
rect 29845 2352 29915 2398
rect 29961 2352 30031 2398
rect 30077 2352 30147 2398
rect 30193 2352 30263 2398
rect 30309 2352 30379 2398
rect 30425 2352 30495 2398
rect 30541 2352 30611 2398
rect 30657 2352 30727 2398
rect 30773 2352 30843 2398
rect 30889 2352 30959 2398
rect 31005 2352 31075 2398
rect 31121 2352 31191 2398
rect 31237 2352 31307 2398
rect 31353 2352 31423 2398
rect 31469 2352 31539 2398
rect 31585 2352 31655 2398
rect 31701 2352 31771 2398
rect 31817 2352 31887 2398
rect 31933 2352 32003 2398
rect 32049 2352 32119 2398
rect 32165 2352 32235 2398
rect 32281 2352 32351 2398
rect 32397 2352 32467 2398
rect 32513 2352 32583 2398
rect 32629 2352 32699 2398
rect 32745 2352 32815 2398
rect 32861 2352 32931 2398
rect 32977 2352 33047 2398
rect 33093 2352 33163 2398
rect 33209 2352 33279 2398
rect 33325 2352 33395 2398
rect 33441 2352 33511 2398
rect 33557 2352 33627 2398
rect 33673 2352 33743 2398
rect 33789 2352 33859 2398
rect 33905 2352 33975 2398
rect 34021 2352 34091 2398
rect 34137 2352 34207 2398
rect 34253 2352 34323 2398
rect 34369 2352 34439 2398
rect 34485 2352 34555 2398
rect 34601 2352 34671 2398
rect 34717 2352 34787 2398
rect 34833 2352 34903 2398
rect 34949 2352 35019 2398
rect 35065 2352 35135 2398
rect 35181 2352 35251 2398
rect 35297 2352 35367 2398
rect 35413 2352 35483 2398
rect 35529 2352 35599 2398
rect 35645 2352 35715 2398
rect 35761 2352 35831 2398
rect 35877 2352 35947 2398
rect 35993 2352 36063 2398
rect 36109 2352 36179 2398
rect 36225 2352 36295 2398
rect 36341 2352 36411 2398
rect 36457 2352 36527 2398
rect 36573 2352 36643 2398
rect 36689 2352 36759 2398
rect 36805 2352 36875 2398
rect 36921 2352 36991 2398
rect 37037 2352 37107 2398
rect 37153 2352 37223 2398
rect 37269 2352 37339 2398
rect 37385 2352 37455 2398
rect 37501 2352 37571 2398
rect 37617 2352 37687 2398
rect 37733 2352 37803 2398
rect 37849 2352 37919 2398
rect 37965 2352 38035 2398
rect 38081 2352 38151 2398
rect 38197 2352 38267 2398
rect 38313 2352 38383 2398
rect 38429 2352 38499 2398
rect 38545 2352 38615 2398
rect 38661 2352 38731 2398
rect 38777 2352 38847 2398
rect 38893 2352 38963 2398
rect 39009 2352 39079 2398
rect 39125 2352 39195 2398
rect 39241 2352 39311 2398
rect 39357 2352 39427 2398
rect 39473 2352 39543 2398
rect 39589 2352 39659 2398
rect 39705 2352 39775 2398
rect 39821 2352 39891 2398
rect 39937 2352 40007 2398
rect 40053 2352 40123 2398
rect 40169 2352 40188 2398
rect 28620 2282 40188 2352
rect 28620 2236 28639 2282
rect 28685 2236 28755 2282
rect 28801 2236 28871 2282
rect 28917 2236 28987 2282
rect 29033 2236 29103 2282
rect 29149 2236 29219 2282
rect 29265 2236 29335 2282
rect 29381 2236 29451 2282
rect 29497 2236 29567 2282
rect 29613 2236 29683 2282
rect 29729 2236 29799 2282
rect 29845 2236 29915 2282
rect 29961 2236 30031 2282
rect 30077 2236 30147 2282
rect 30193 2236 30263 2282
rect 30309 2236 30379 2282
rect 30425 2236 30495 2282
rect 30541 2236 30611 2282
rect 30657 2236 30727 2282
rect 30773 2236 30843 2282
rect 30889 2236 30959 2282
rect 31005 2236 31075 2282
rect 31121 2236 31191 2282
rect 31237 2236 31307 2282
rect 31353 2236 31423 2282
rect 31469 2236 31539 2282
rect 31585 2236 31655 2282
rect 31701 2236 31771 2282
rect 31817 2236 31887 2282
rect 31933 2236 32003 2282
rect 32049 2236 32119 2282
rect 32165 2236 32235 2282
rect 32281 2236 32351 2282
rect 32397 2236 32467 2282
rect 32513 2236 32583 2282
rect 32629 2236 32699 2282
rect 32745 2236 32815 2282
rect 32861 2236 32931 2282
rect 32977 2236 33047 2282
rect 33093 2236 33163 2282
rect 33209 2236 33279 2282
rect 33325 2236 33395 2282
rect 33441 2236 33511 2282
rect 33557 2236 33627 2282
rect 33673 2236 33743 2282
rect 33789 2236 33859 2282
rect 33905 2236 33975 2282
rect 34021 2236 34091 2282
rect 34137 2236 34207 2282
rect 34253 2236 34323 2282
rect 34369 2236 34439 2282
rect 34485 2236 34555 2282
rect 34601 2236 34671 2282
rect 34717 2236 34787 2282
rect 34833 2236 34903 2282
rect 34949 2236 35019 2282
rect 35065 2236 35135 2282
rect 35181 2236 35251 2282
rect 35297 2236 35367 2282
rect 35413 2236 35483 2282
rect 35529 2236 35599 2282
rect 35645 2236 35715 2282
rect 35761 2236 35831 2282
rect 35877 2236 35947 2282
rect 35993 2236 36063 2282
rect 36109 2236 36179 2282
rect 36225 2236 36295 2282
rect 36341 2236 36411 2282
rect 36457 2236 36527 2282
rect 36573 2236 36643 2282
rect 36689 2236 36759 2282
rect 36805 2236 36875 2282
rect 36921 2236 36991 2282
rect 37037 2236 37107 2282
rect 37153 2236 37223 2282
rect 37269 2236 37339 2282
rect 37385 2236 37455 2282
rect 37501 2236 37571 2282
rect 37617 2236 37687 2282
rect 37733 2236 37803 2282
rect 37849 2236 37919 2282
rect 37965 2236 38035 2282
rect 38081 2236 38151 2282
rect 38197 2236 38267 2282
rect 38313 2236 38383 2282
rect 38429 2236 38499 2282
rect 38545 2236 38615 2282
rect 38661 2236 38731 2282
rect 38777 2236 38847 2282
rect 38893 2236 38963 2282
rect 39009 2236 39079 2282
rect 39125 2236 39195 2282
rect 39241 2236 39311 2282
rect 39357 2236 39427 2282
rect 39473 2236 39543 2282
rect 39589 2236 39659 2282
rect 39705 2236 39775 2282
rect 39821 2236 39891 2282
rect 39937 2236 40007 2282
rect 40053 2236 40123 2282
rect 40169 2236 40188 2282
rect 28620 2166 40188 2236
rect 28620 2120 28639 2166
rect 28685 2120 28755 2166
rect 28801 2120 28871 2166
rect 28917 2120 28987 2166
rect 29033 2120 29103 2166
rect 29149 2120 29219 2166
rect 29265 2120 29335 2166
rect 29381 2120 29451 2166
rect 29497 2120 29567 2166
rect 29613 2120 29683 2166
rect 29729 2120 29799 2166
rect 29845 2120 29915 2166
rect 29961 2120 30031 2166
rect 30077 2120 30147 2166
rect 30193 2120 30263 2166
rect 30309 2120 30379 2166
rect 30425 2120 30495 2166
rect 30541 2120 30611 2166
rect 30657 2120 30727 2166
rect 30773 2120 30843 2166
rect 30889 2120 30959 2166
rect 31005 2120 31075 2166
rect 31121 2120 31191 2166
rect 31237 2120 31307 2166
rect 31353 2120 31423 2166
rect 31469 2120 31539 2166
rect 31585 2120 31655 2166
rect 31701 2120 31771 2166
rect 31817 2120 31887 2166
rect 31933 2120 32003 2166
rect 32049 2120 32119 2166
rect 32165 2120 32235 2166
rect 32281 2120 32351 2166
rect 32397 2120 32467 2166
rect 32513 2120 32583 2166
rect 32629 2120 32699 2166
rect 32745 2120 32815 2166
rect 32861 2120 32931 2166
rect 32977 2120 33047 2166
rect 33093 2120 33163 2166
rect 33209 2120 33279 2166
rect 33325 2120 33395 2166
rect 33441 2120 33511 2166
rect 33557 2120 33627 2166
rect 33673 2120 33743 2166
rect 33789 2120 33859 2166
rect 33905 2120 33975 2166
rect 34021 2120 34091 2166
rect 34137 2120 34207 2166
rect 34253 2120 34323 2166
rect 34369 2120 34439 2166
rect 34485 2120 34555 2166
rect 34601 2120 34671 2166
rect 34717 2120 34787 2166
rect 34833 2120 34903 2166
rect 34949 2120 35019 2166
rect 35065 2120 35135 2166
rect 35181 2120 35251 2166
rect 35297 2120 35367 2166
rect 35413 2120 35483 2166
rect 35529 2120 35599 2166
rect 35645 2120 35715 2166
rect 35761 2120 35831 2166
rect 35877 2120 35947 2166
rect 35993 2120 36063 2166
rect 36109 2120 36179 2166
rect 36225 2120 36295 2166
rect 36341 2120 36411 2166
rect 36457 2120 36527 2166
rect 36573 2120 36643 2166
rect 36689 2120 36759 2166
rect 36805 2120 36875 2166
rect 36921 2120 36991 2166
rect 37037 2120 37107 2166
rect 37153 2120 37223 2166
rect 37269 2120 37339 2166
rect 37385 2120 37455 2166
rect 37501 2120 37571 2166
rect 37617 2120 37687 2166
rect 37733 2120 37803 2166
rect 37849 2120 37919 2166
rect 37965 2120 38035 2166
rect 38081 2120 38151 2166
rect 38197 2120 38267 2166
rect 38313 2120 38383 2166
rect 38429 2120 38499 2166
rect 38545 2120 38615 2166
rect 38661 2120 38731 2166
rect 38777 2120 38847 2166
rect 38893 2120 38963 2166
rect 39009 2120 39079 2166
rect 39125 2120 39195 2166
rect 39241 2120 39311 2166
rect 39357 2120 39427 2166
rect 39473 2120 39543 2166
rect 39589 2120 39659 2166
rect 39705 2120 39775 2166
rect 39821 2120 39891 2166
rect 39937 2120 40007 2166
rect 40053 2120 40123 2166
rect 40169 2120 40188 2166
rect 28620 2050 40188 2120
rect 28620 2004 28639 2050
rect 28685 2004 28755 2050
rect 28801 2004 28871 2050
rect 28917 2004 28987 2050
rect 29033 2004 29103 2050
rect 29149 2004 29219 2050
rect 29265 2004 29335 2050
rect 29381 2004 29451 2050
rect 29497 2004 29567 2050
rect 29613 2004 29683 2050
rect 29729 2004 29799 2050
rect 29845 2004 29915 2050
rect 29961 2004 30031 2050
rect 30077 2004 30147 2050
rect 30193 2004 30263 2050
rect 30309 2004 30379 2050
rect 30425 2004 30495 2050
rect 30541 2004 30611 2050
rect 30657 2004 30727 2050
rect 30773 2004 30843 2050
rect 30889 2004 30959 2050
rect 31005 2004 31075 2050
rect 31121 2004 31191 2050
rect 31237 2004 31307 2050
rect 31353 2004 31423 2050
rect 31469 2004 31539 2050
rect 31585 2004 31655 2050
rect 31701 2004 31771 2050
rect 31817 2004 31887 2050
rect 31933 2004 32003 2050
rect 32049 2004 32119 2050
rect 32165 2004 32235 2050
rect 32281 2004 32351 2050
rect 32397 2004 32467 2050
rect 32513 2004 32583 2050
rect 32629 2004 32699 2050
rect 32745 2004 32815 2050
rect 32861 2004 32931 2050
rect 32977 2004 33047 2050
rect 33093 2004 33163 2050
rect 33209 2004 33279 2050
rect 33325 2004 33395 2050
rect 33441 2004 33511 2050
rect 33557 2004 33627 2050
rect 33673 2004 33743 2050
rect 33789 2004 33859 2050
rect 33905 2004 33975 2050
rect 34021 2004 34091 2050
rect 34137 2004 34207 2050
rect 34253 2004 34323 2050
rect 34369 2004 34439 2050
rect 34485 2004 34555 2050
rect 34601 2004 34671 2050
rect 34717 2004 34787 2050
rect 34833 2004 34903 2050
rect 34949 2004 35019 2050
rect 35065 2004 35135 2050
rect 35181 2004 35251 2050
rect 35297 2004 35367 2050
rect 35413 2004 35483 2050
rect 35529 2004 35599 2050
rect 35645 2004 35715 2050
rect 35761 2004 35831 2050
rect 35877 2004 35947 2050
rect 35993 2004 36063 2050
rect 36109 2004 36179 2050
rect 36225 2004 36295 2050
rect 36341 2004 36411 2050
rect 36457 2004 36527 2050
rect 36573 2004 36643 2050
rect 36689 2004 36759 2050
rect 36805 2004 36875 2050
rect 36921 2004 36991 2050
rect 37037 2004 37107 2050
rect 37153 2004 37223 2050
rect 37269 2004 37339 2050
rect 37385 2004 37455 2050
rect 37501 2004 37571 2050
rect 37617 2004 37687 2050
rect 37733 2004 37803 2050
rect 37849 2004 37919 2050
rect 37965 2004 38035 2050
rect 38081 2004 38151 2050
rect 38197 2004 38267 2050
rect 38313 2004 38383 2050
rect 38429 2004 38499 2050
rect 38545 2004 38615 2050
rect 38661 2004 38731 2050
rect 38777 2004 38847 2050
rect 38893 2004 38963 2050
rect 39009 2004 39079 2050
rect 39125 2004 39195 2050
rect 39241 2004 39311 2050
rect 39357 2004 39427 2050
rect 39473 2004 39543 2050
rect 39589 2004 39659 2050
rect 39705 2004 39775 2050
rect 39821 2004 39891 2050
rect 39937 2004 40007 2050
rect 40053 2004 40123 2050
rect 40169 2004 40188 2050
rect 28620 1934 40188 2004
rect 28620 1888 28639 1934
rect 28685 1888 28755 1934
rect 28801 1888 28871 1934
rect 28917 1888 28987 1934
rect 29033 1888 29103 1934
rect 29149 1888 29219 1934
rect 29265 1888 29335 1934
rect 29381 1888 29451 1934
rect 29497 1888 29567 1934
rect 29613 1888 29683 1934
rect 29729 1888 29799 1934
rect 29845 1888 29915 1934
rect 29961 1888 30031 1934
rect 30077 1888 30147 1934
rect 30193 1888 30263 1934
rect 30309 1888 30379 1934
rect 30425 1888 30495 1934
rect 30541 1888 30611 1934
rect 30657 1888 30727 1934
rect 30773 1888 30843 1934
rect 30889 1888 30959 1934
rect 31005 1888 31075 1934
rect 31121 1888 31191 1934
rect 31237 1888 31307 1934
rect 31353 1888 31423 1934
rect 31469 1888 31539 1934
rect 31585 1888 31655 1934
rect 31701 1888 31771 1934
rect 31817 1888 31887 1934
rect 31933 1888 32003 1934
rect 32049 1888 32119 1934
rect 32165 1888 32235 1934
rect 32281 1888 32351 1934
rect 32397 1888 32467 1934
rect 32513 1888 32583 1934
rect 32629 1888 32699 1934
rect 32745 1888 32815 1934
rect 32861 1888 32931 1934
rect 32977 1888 33047 1934
rect 33093 1888 33163 1934
rect 33209 1888 33279 1934
rect 33325 1888 33395 1934
rect 33441 1888 33511 1934
rect 33557 1888 33627 1934
rect 33673 1888 33743 1934
rect 33789 1888 33859 1934
rect 33905 1888 33975 1934
rect 34021 1888 34091 1934
rect 34137 1888 34207 1934
rect 34253 1888 34323 1934
rect 34369 1888 34439 1934
rect 34485 1888 34555 1934
rect 34601 1888 34671 1934
rect 34717 1888 34787 1934
rect 34833 1888 34903 1934
rect 34949 1888 35019 1934
rect 35065 1888 35135 1934
rect 35181 1888 35251 1934
rect 35297 1888 35367 1934
rect 35413 1888 35483 1934
rect 35529 1888 35599 1934
rect 35645 1888 35715 1934
rect 35761 1888 35831 1934
rect 35877 1888 35947 1934
rect 35993 1888 36063 1934
rect 36109 1888 36179 1934
rect 36225 1888 36295 1934
rect 36341 1888 36411 1934
rect 36457 1888 36527 1934
rect 36573 1888 36643 1934
rect 36689 1888 36759 1934
rect 36805 1888 36875 1934
rect 36921 1888 36991 1934
rect 37037 1888 37107 1934
rect 37153 1888 37223 1934
rect 37269 1888 37339 1934
rect 37385 1888 37455 1934
rect 37501 1888 37571 1934
rect 37617 1888 37687 1934
rect 37733 1888 37803 1934
rect 37849 1888 37919 1934
rect 37965 1888 38035 1934
rect 38081 1888 38151 1934
rect 38197 1888 38267 1934
rect 38313 1888 38383 1934
rect 38429 1888 38499 1934
rect 38545 1888 38615 1934
rect 38661 1888 38731 1934
rect 38777 1888 38847 1934
rect 38893 1888 38963 1934
rect 39009 1888 39079 1934
rect 39125 1888 39195 1934
rect 39241 1888 39311 1934
rect 39357 1888 39427 1934
rect 39473 1888 39543 1934
rect 39589 1888 39659 1934
rect 39705 1888 39775 1934
rect 39821 1888 39891 1934
rect 39937 1888 40007 1934
rect 40053 1888 40123 1934
rect 40169 1888 40188 1934
rect 28620 1818 40188 1888
rect 28620 1772 28639 1818
rect 28685 1772 28755 1818
rect 28801 1772 28871 1818
rect 28917 1772 28987 1818
rect 29033 1772 29103 1818
rect 29149 1772 29219 1818
rect 29265 1772 29335 1818
rect 29381 1772 29451 1818
rect 29497 1772 29567 1818
rect 29613 1772 29683 1818
rect 29729 1772 29799 1818
rect 29845 1772 29915 1818
rect 29961 1772 30031 1818
rect 30077 1772 30147 1818
rect 30193 1772 30263 1818
rect 30309 1772 30379 1818
rect 30425 1772 30495 1818
rect 30541 1772 30611 1818
rect 30657 1772 30727 1818
rect 30773 1772 30843 1818
rect 30889 1772 30959 1818
rect 31005 1772 31075 1818
rect 31121 1772 31191 1818
rect 31237 1772 31307 1818
rect 31353 1772 31423 1818
rect 31469 1772 31539 1818
rect 31585 1772 31655 1818
rect 31701 1772 31771 1818
rect 31817 1772 31887 1818
rect 31933 1772 32003 1818
rect 32049 1772 32119 1818
rect 32165 1772 32235 1818
rect 32281 1772 32351 1818
rect 32397 1772 32467 1818
rect 32513 1772 32583 1818
rect 32629 1772 32699 1818
rect 32745 1772 32815 1818
rect 32861 1772 32931 1818
rect 32977 1772 33047 1818
rect 33093 1772 33163 1818
rect 33209 1772 33279 1818
rect 33325 1772 33395 1818
rect 33441 1772 33511 1818
rect 33557 1772 33627 1818
rect 33673 1772 33743 1818
rect 33789 1772 33859 1818
rect 33905 1772 33975 1818
rect 34021 1772 34091 1818
rect 34137 1772 34207 1818
rect 34253 1772 34323 1818
rect 34369 1772 34439 1818
rect 34485 1772 34555 1818
rect 34601 1772 34671 1818
rect 34717 1772 34787 1818
rect 34833 1772 34903 1818
rect 34949 1772 35019 1818
rect 35065 1772 35135 1818
rect 35181 1772 35251 1818
rect 35297 1772 35367 1818
rect 35413 1772 35483 1818
rect 35529 1772 35599 1818
rect 35645 1772 35715 1818
rect 35761 1772 35831 1818
rect 35877 1772 35947 1818
rect 35993 1772 36063 1818
rect 36109 1772 36179 1818
rect 36225 1772 36295 1818
rect 36341 1772 36411 1818
rect 36457 1772 36527 1818
rect 36573 1772 36643 1818
rect 36689 1772 36759 1818
rect 36805 1772 36875 1818
rect 36921 1772 36991 1818
rect 37037 1772 37107 1818
rect 37153 1772 37223 1818
rect 37269 1772 37339 1818
rect 37385 1772 37455 1818
rect 37501 1772 37571 1818
rect 37617 1772 37687 1818
rect 37733 1772 37803 1818
rect 37849 1772 37919 1818
rect 37965 1772 38035 1818
rect 38081 1772 38151 1818
rect 38197 1772 38267 1818
rect 38313 1772 38383 1818
rect 38429 1772 38499 1818
rect 38545 1772 38615 1818
rect 38661 1772 38731 1818
rect 38777 1772 38847 1818
rect 38893 1772 38963 1818
rect 39009 1772 39079 1818
rect 39125 1772 39195 1818
rect 39241 1772 39311 1818
rect 39357 1772 39427 1818
rect 39473 1772 39543 1818
rect 39589 1772 39659 1818
rect 39705 1772 39775 1818
rect 39821 1772 39891 1818
rect 39937 1772 40007 1818
rect 40053 1772 40123 1818
rect 40169 1772 40188 1818
rect 28620 1702 40188 1772
rect 28620 1656 28639 1702
rect 28685 1656 28755 1702
rect 28801 1656 28871 1702
rect 28917 1656 28987 1702
rect 29033 1656 29103 1702
rect 29149 1656 29219 1702
rect 29265 1656 29335 1702
rect 29381 1656 29451 1702
rect 29497 1656 29567 1702
rect 29613 1656 29683 1702
rect 29729 1656 29799 1702
rect 29845 1656 29915 1702
rect 29961 1656 30031 1702
rect 30077 1656 30147 1702
rect 30193 1656 30263 1702
rect 30309 1656 30379 1702
rect 30425 1656 30495 1702
rect 30541 1656 30611 1702
rect 30657 1656 30727 1702
rect 30773 1656 30843 1702
rect 30889 1656 30959 1702
rect 31005 1656 31075 1702
rect 31121 1656 31191 1702
rect 31237 1656 31307 1702
rect 31353 1656 31423 1702
rect 31469 1656 31539 1702
rect 31585 1656 31655 1702
rect 31701 1656 31771 1702
rect 31817 1656 31887 1702
rect 31933 1656 32003 1702
rect 32049 1656 32119 1702
rect 32165 1656 32235 1702
rect 32281 1656 32351 1702
rect 32397 1656 32467 1702
rect 32513 1656 32583 1702
rect 32629 1656 32699 1702
rect 32745 1656 32815 1702
rect 32861 1656 32931 1702
rect 32977 1656 33047 1702
rect 33093 1656 33163 1702
rect 33209 1656 33279 1702
rect 33325 1656 33395 1702
rect 33441 1656 33511 1702
rect 33557 1656 33627 1702
rect 33673 1656 33743 1702
rect 33789 1656 33859 1702
rect 33905 1656 33975 1702
rect 34021 1656 34091 1702
rect 34137 1656 34207 1702
rect 34253 1656 34323 1702
rect 34369 1656 34439 1702
rect 34485 1656 34555 1702
rect 34601 1656 34671 1702
rect 34717 1656 34787 1702
rect 34833 1656 34903 1702
rect 34949 1656 35019 1702
rect 35065 1656 35135 1702
rect 35181 1656 35251 1702
rect 35297 1656 35367 1702
rect 35413 1656 35483 1702
rect 35529 1656 35599 1702
rect 35645 1656 35715 1702
rect 35761 1656 35831 1702
rect 35877 1656 35947 1702
rect 35993 1656 36063 1702
rect 36109 1656 36179 1702
rect 36225 1656 36295 1702
rect 36341 1656 36411 1702
rect 36457 1656 36527 1702
rect 36573 1656 36643 1702
rect 36689 1656 36759 1702
rect 36805 1656 36875 1702
rect 36921 1656 36991 1702
rect 37037 1656 37107 1702
rect 37153 1656 37223 1702
rect 37269 1656 37339 1702
rect 37385 1656 37455 1702
rect 37501 1656 37571 1702
rect 37617 1656 37687 1702
rect 37733 1656 37803 1702
rect 37849 1656 37919 1702
rect 37965 1656 38035 1702
rect 38081 1656 38151 1702
rect 38197 1656 38267 1702
rect 38313 1656 38383 1702
rect 38429 1656 38499 1702
rect 38545 1656 38615 1702
rect 38661 1656 38731 1702
rect 38777 1656 38847 1702
rect 38893 1656 38963 1702
rect 39009 1656 39079 1702
rect 39125 1656 39195 1702
rect 39241 1656 39311 1702
rect 39357 1656 39427 1702
rect 39473 1656 39543 1702
rect 39589 1656 39659 1702
rect 39705 1656 39775 1702
rect 39821 1656 39891 1702
rect 39937 1656 40007 1702
rect 40053 1656 40123 1702
rect 40169 1656 40188 1702
rect 28620 1637 40188 1656
rect 50826 3906 56594 3925
rect 50826 3860 50845 3906
rect 50891 3860 50961 3906
rect 51007 3860 51077 3906
rect 51123 3860 51193 3906
rect 51239 3860 51309 3906
rect 51355 3860 51425 3906
rect 51471 3860 51541 3906
rect 51587 3860 51657 3906
rect 51703 3860 51773 3906
rect 51819 3860 51889 3906
rect 51935 3860 52005 3906
rect 52051 3860 52121 3906
rect 52167 3860 52237 3906
rect 52283 3860 52353 3906
rect 52399 3860 52469 3906
rect 52515 3860 52585 3906
rect 52631 3860 52701 3906
rect 52747 3860 52817 3906
rect 52863 3860 52933 3906
rect 52979 3860 53049 3906
rect 53095 3860 53165 3906
rect 53211 3860 53281 3906
rect 53327 3860 53397 3906
rect 53443 3860 53513 3906
rect 53559 3860 53629 3906
rect 53675 3860 53745 3906
rect 53791 3860 53861 3906
rect 53907 3860 53977 3906
rect 54023 3860 54093 3906
rect 54139 3860 54209 3906
rect 54255 3860 54325 3906
rect 54371 3860 54441 3906
rect 54487 3860 54557 3906
rect 54603 3860 54673 3906
rect 54719 3860 54789 3906
rect 54835 3860 54905 3906
rect 54951 3860 55021 3906
rect 55067 3860 55137 3906
rect 55183 3860 55253 3906
rect 55299 3860 55369 3906
rect 55415 3860 55485 3906
rect 55531 3860 55601 3906
rect 55647 3860 55717 3906
rect 55763 3860 55833 3906
rect 55879 3860 55949 3906
rect 55995 3860 56065 3906
rect 56111 3860 56181 3906
rect 56227 3860 56297 3906
rect 56343 3860 56413 3906
rect 56459 3860 56529 3906
rect 56575 3860 56594 3906
rect 50826 3790 56594 3860
rect 50826 3744 50845 3790
rect 50891 3744 50961 3790
rect 51007 3744 51077 3790
rect 51123 3744 51193 3790
rect 51239 3744 51309 3790
rect 51355 3744 51425 3790
rect 51471 3744 51541 3790
rect 51587 3744 51657 3790
rect 51703 3744 51773 3790
rect 51819 3744 51889 3790
rect 51935 3744 52005 3790
rect 52051 3744 52121 3790
rect 52167 3744 52237 3790
rect 52283 3744 52353 3790
rect 52399 3744 52469 3790
rect 52515 3744 52585 3790
rect 52631 3744 52701 3790
rect 52747 3744 52817 3790
rect 52863 3744 52933 3790
rect 52979 3744 53049 3790
rect 53095 3744 53165 3790
rect 53211 3744 53281 3790
rect 53327 3744 53397 3790
rect 53443 3744 53513 3790
rect 53559 3744 53629 3790
rect 53675 3744 53745 3790
rect 53791 3744 53861 3790
rect 53907 3744 53977 3790
rect 54023 3744 54093 3790
rect 54139 3744 54209 3790
rect 54255 3744 54325 3790
rect 54371 3744 54441 3790
rect 54487 3744 54557 3790
rect 54603 3744 54673 3790
rect 54719 3744 54789 3790
rect 54835 3744 54905 3790
rect 54951 3744 55021 3790
rect 55067 3744 55137 3790
rect 55183 3744 55253 3790
rect 55299 3744 55369 3790
rect 55415 3744 55485 3790
rect 55531 3744 55601 3790
rect 55647 3744 55717 3790
rect 55763 3744 55833 3790
rect 55879 3744 55949 3790
rect 55995 3744 56065 3790
rect 56111 3744 56181 3790
rect 56227 3744 56297 3790
rect 56343 3744 56413 3790
rect 56459 3744 56529 3790
rect 56575 3744 56594 3790
rect 50826 3674 56594 3744
rect 50826 3628 50845 3674
rect 50891 3628 50961 3674
rect 51007 3628 51077 3674
rect 51123 3628 51193 3674
rect 51239 3628 51309 3674
rect 51355 3628 51425 3674
rect 51471 3628 51541 3674
rect 51587 3628 51657 3674
rect 51703 3628 51773 3674
rect 51819 3628 51889 3674
rect 51935 3628 52005 3674
rect 52051 3628 52121 3674
rect 52167 3628 52237 3674
rect 52283 3628 52353 3674
rect 52399 3628 52469 3674
rect 52515 3628 52585 3674
rect 52631 3628 52701 3674
rect 52747 3628 52817 3674
rect 52863 3628 52933 3674
rect 52979 3628 53049 3674
rect 53095 3628 53165 3674
rect 53211 3628 53281 3674
rect 53327 3628 53397 3674
rect 53443 3628 53513 3674
rect 53559 3628 53629 3674
rect 53675 3628 53745 3674
rect 53791 3628 53861 3674
rect 53907 3628 53977 3674
rect 54023 3628 54093 3674
rect 54139 3628 54209 3674
rect 54255 3628 54325 3674
rect 54371 3628 54441 3674
rect 54487 3628 54557 3674
rect 54603 3628 54673 3674
rect 54719 3628 54789 3674
rect 54835 3628 54905 3674
rect 54951 3628 55021 3674
rect 55067 3628 55137 3674
rect 55183 3628 55253 3674
rect 55299 3628 55369 3674
rect 55415 3628 55485 3674
rect 55531 3628 55601 3674
rect 55647 3628 55717 3674
rect 55763 3628 55833 3674
rect 55879 3628 55949 3674
rect 55995 3628 56065 3674
rect 56111 3628 56181 3674
rect 56227 3628 56297 3674
rect 56343 3628 56413 3674
rect 56459 3628 56529 3674
rect 56575 3628 56594 3674
rect 50826 3558 56594 3628
rect 50826 3512 50845 3558
rect 50891 3512 50961 3558
rect 51007 3512 51077 3558
rect 51123 3512 51193 3558
rect 51239 3512 51309 3558
rect 51355 3512 51425 3558
rect 51471 3512 51541 3558
rect 51587 3512 51657 3558
rect 51703 3512 51773 3558
rect 51819 3512 51889 3558
rect 51935 3512 52005 3558
rect 52051 3512 52121 3558
rect 52167 3512 52237 3558
rect 52283 3512 52353 3558
rect 52399 3512 52469 3558
rect 52515 3512 52585 3558
rect 52631 3512 52701 3558
rect 52747 3512 52817 3558
rect 52863 3512 52933 3558
rect 52979 3512 53049 3558
rect 53095 3512 53165 3558
rect 53211 3512 53281 3558
rect 53327 3512 53397 3558
rect 53443 3512 53513 3558
rect 53559 3512 53629 3558
rect 53675 3512 53745 3558
rect 53791 3512 53861 3558
rect 53907 3512 53977 3558
rect 54023 3512 54093 3558
rect 54139 3512 54209 3558
rect 54255 3512 54325 3558
rect 54371 3512 54441 3558
rect 54487 3512 54557 3558
rect 54603 3512 54673 3558
rect 54719 3512 54789 3558
rect 54835 3512 54905 3558
rect 54951 3512 55021 3558
rect 55067 3512 55137 3558
rect 55183 3512 55253 3558
rect 55299 3512 55369 3558
rect 55415 3512 55485 3558
rect 55531 3512 55601 3558
rect 55647 3512 55717 3558
rect 55763 3512 55833 3558
rect 55879 3512 55949 3558
rect 55995 3512 56065 3558
rect 56111 3512 56181 3558
rect 56227 3512 56297 3558
rect 56343 3512 56413 3558
rect 56459 3512 56529 3558
rect 56575 3512 56594 3558
rect 50826 3442 56594 3512
rect 50826 3396 50845 3442
rect 50891 3396 50961 3442
rect 51007 3396 51077 3442
rect 51123 3396 51193 3442
rect 51239 3396 51309 3442
rect 51355 3396 51425 3442
rect 51471 3396 51541 3442
rect 51587 3396 51657 3442
rect 51703 3396 51773 3442
rect 51819 3396 51889 3442
rect 51935 3396 52005 3442
rect 52051 3396 52121 3442
rect 52167 3396 52237 3442
rect 52283 3396 52353 3442
rect 52399 3396 52469 3442
rect 52515 3396 52585 3442
rect 52631 3396 52701 3442
rect 52747 3396 52817 3442
rect 52863 3396 52933 3442
rect 52979 3396 53049 3442
rect 53095 3396 53165 3442
rect 53211 3396 53281 3442
rect 53327 3396 53397 3442
rect 53443 3396 53513 3442
rect 53559 3396 53629 3442
rect 53675 3396 53745 3442
rect 53791 3396 53861 3442
rect 53907 3396 53977 3442
rect 54023 3396 54093 3442
rect 54139 3396 54209 3442
rect 54255 3396 54325 3442
rect 54371 3396 54441 3442
rect 54487 3396 54557 3442
rect 54603 3396 54673 3442
rect 54719 3396 54789 3442
rect 54835 3396 54905 3442
rect 54951 3396 55021 3442
rect 55067 3396 55137 3442
rect 55183 3396 55253 3442
rect 55299 3396 55369 3442
rect 55415 3396 55485 3442
rect 55531 3396 55601 3442
rect 55647 3396 55717 3442
rect 55763 3396 55833 3442
rect 55879 3396 55949 3442
rect 55995 3396 56065 3442
rect 56111 3396 56181 3442
rect 56227 3396 56297 3442
rect 56343 3396 56413 3442
rect 56459 3396 56529 3442
rect 56575 3396 56594 3442
rect 50826 3326 56594 3396
rect 50826 3280 50845 3326
rect 50891 3280 50961 3326
rect 51007 3280 51077 3326
rect 51123 3280 51193 3326
rect 51239 3280 51309 3326
rect 51355 3280 51425 3326
rect 51471 3280 51541 3326
rect 51587 3280 51657 3326
rect 51703 3280 51773 3326
rect 51819 3280 51889 3326
rect 51935 3280 52005 3326
rect 52051 3280 52121 3326
rect 52167 3280 52237 3326
rect 52283 3280 52353 3326
rect 52399 3280 52469 3326
rect 52515 3280 52585 3326
rect 52631 3280 52701 3326
rect 52747 3280 52817 3326
rect 52863 3280 52933 3326
rect 52979 3280 53049 3326
rect 53095 3280 53165 3326
rect 53211 3280 53281 3326
rect 53327 3280 53397 3326
rect 53443 3280 53513 3326
rect 53559 3280 53629 3326
rect 53675 3280 53745 3326
rect 53791 3280 53861 3326
rect 53907 3280 53977 3326
rect 54023 3280 54093 3326
rect 54139 3280 54209 3326
rect 54255 3280 54325 3326
rect 54371 3280 54441 3326
rect 54487 3280 54557 3326
rect 54603 3280 54673 3326
rect 54719 3280 54789 3326
rect 54835 3280 54905 3326
rect 54951 3280 55021 3326
rect 55067 3280 55137 3326
rect 55183 3280 55253 3326
rect 55299 3280 55369 3326
rect 55415 3280 55485 3326
rect 55531 3280 55601 3326
rect 55647 3280 55717 3326
rect 55763 3280 55833 3326
rect 55879 3280 55949 3326
rect 55995 3280 56065 3326
rect 56111 3280 56181 3326
rect 56227 3280 56297 3326
rect 56343 3280 56413 3326
rect 56459 3280 56529 3326
rect 56575 3280 56594 3326
rect 50826 3210 56594 3280
rect 50826 3164 50845 3210
rect 50891 3164 50961 3210
rect 51007 3164 51077 3210
rect 51123 3164 51193 3210
rect 51239 3164 51309 3210
rect 51355 3164 51425 3210
rect 51471 3164 51541 3210
rect 51587 3164 51657 3210
rect 51703 3164 51773 3210
rect 51819 3164 51889 3210
rect 51935 3164 52005 3210
rect 52051 3164 52121 3210
rect 52167 3164 52237 3210
rect 52283 3164 52353 3210
rect 52399 3164 52469 3210
rect 52515 3164 52585 3210
rect 52631 3164 52701 3210
rect 52747 3164 52817 3210
rect 52863 3164 52933 3210
rect 52979 3164 53049 3210
rect 53095 3164 53165 3210
rect 53211 3164 53281 3210
rect 53327 3164 53397 3210
rect 53443 3164 53513 3210
rect 53559 3164 53629 3210
rect 53675 3164 53745 3210
rect 53791 3164 53861 3210
rect 53907 3164 53977 3210
rect 54023 3164 54093 3210
rect 54139 3164 54209 3210
rect 54255 3164 54325 3210
rect 54371 3164 54441 3210
rect 54487 3164 54557 3210
rect 54603 3164 54673 3210
rect 54719 3164 54789 3210
rect 54835 3164 54905 3210
rect 54951 3164 55021 3210
rect 55067 3164 55137 3210
rect 55183 3164 55253 3210
rect 55299 3164 55369 3210
rect 55415 3164 55485 3210
rect 55531 3164 55601 3210
rect 55647 3164 55717 3210
rect 55763 3164 55833 3210
rect 55879 3164 55949 3210
rect 55995 3164 56065 3210
rect 56111 3164 56181 3210
rect 56227 3164 56297 3210
rect 56343 3164 56413 3210
rect 56459 3164 56529 3210
rect 56575 3164 56594 3210
rect 50826 3094 56594 3164
rect 50826 3048 50845 3094
rect 50891 3048 50961 3094
rect 51007 3048 51077 3094
rect 51123 3048 51193 3094
rect 51239 3048 51309 3094
rect 51355 3048 51425 3094
rect 51471 3048 51541 3094
rect 51587 3048 51657 3094
rect 51703 3048 51773 3094
rect 51819 3048 51889 3094
rect 51935 3048 52005 3094
rect 52051 3048 52121 3094
rect 52167 3048 52237 3094
rect 52283 3048 52353 3094
rect 52399 3048 52469 3094
rect 52515 3048 52585 3094
rect 52631 3048 52701 3094
rect 52747 3048 52817 3094
rect 52863 3048 52933 3094
rect 52979 3048 53049 3094
rect 53095 3048 53165 3094
rect 53211 3048 53281 3094
rect 53327 3048 53397 3094
rect 53443 3048 53513 3094
rect 53559 3048 53629 3094
rect 53675 3048 53745 3094
rect 53791 3048 53861 3094
rect 53907 3048 53977 3094
rect 54023 3048 54093 3094
rect 54139 3048 54209 3094
rect 54255 3048 54325 3094
rect 54371 3048 54441 3094
rect 54487 3048 54557 3094
rect 54603 3048 54673 3094
rect 54719 3048 54789 3094
rect 54835 3048 54905 3094
rect 54951 3048 55021 3094
rect 55067 3048 55137 3094
rect 55183 3048 55253 3094
rect 55299 3048 55369 3094
rect 55415 3048 55485 3094
rect 55531 3048 55601 3094
rect 55647 3048 55717 3094
rect 55763 3048 55833 3094
rect 55879 3048 55949 3094
rect 55995 3048 56065 3094
rect 56111 3048 56181 3094
rect 56227 3048 56297 3094
rect 56343 3048 56413 3094
rect 56459 3048 56529 3094
rect 56575 3048 56594 3094
rect 50826 2978 56594 3048
rect 50826 2932 50845 2978
rect 50891 2932 50961 2978
rect 51007 2932 51077 2978
rect 51123 2932 51193 2978
rect 51239 2932 51309 2978
rect 51355 2932 51425 2978
rect 51471 2932 51541 2978
rect 51587 2932 51657 2978
rect 51703 2932 51773 2978
rect 51819 2932 51889 2978
rect 51935 2932 52005 2978
rect 52051 2932 52121 2978
rect 52167 2932 52237 2978
rect 52283 2932 52353 2978
rect 52399 2932 52469 2978
rect 52515 2932 52585 2978
rect 52631 2932 52701 2978
rect 52747 2932 52817 2978
rect 52863 2932 52933 2978
rect 52979 2932 53049 2978
rect 53095 2932 53165 2978
rect 53211 2932 53281 2978
rect 53327 2932 53397 2978
rect 53443 2932 53513 2978
rect 53559 2932 53629 2978
rect 53675 2932 53745 2978
rect 53791 2932 53861 2978
rect 53907 2932 53977 2978
rect 54023 2932 54093 2978
rect 54139 2932 54209 2978
rect 54255 2932 54325 2978
rect 54371 2932 54441 2978
rect 54487 2932 54557 2978
rect 54603 2932 54673 2978
rect 54719 2932 54789 2978
rect 54835 2932 54905 2978
rect 54951 2932 55021 2978
rect 55067 2932 55137 2978
rect 55183 2932 55253 2978
rect 55299 2932 55369 2978
rect 55415 2932 55485 2978
rect 55531 2932 55601 2978
rect 55647 2932 55717 2978
rect 55763 2932 55833 2978
rect 55879 2932 55949 2978
rect 55995 2932 56065 2978
rect 56111 2932 56181 2978
rect 56227 2932 56297 2978
rect 56343 2932 56413 2978
rect 56459 2932 56529 2978
rect 56575 2932 56594 2978
rect 50826 2862 56594 2932
rect 50826 2816 50845 2862
rect 50891 2816 50961 2862
rect 51007 2816 51077 2862
rect 51123 2816 51193 2862
rect 51239 2816 51309 2862
rect 51355 2816 51425 2862
rect 51471 2816 51541 2862
rect 51587 2816 51657 2862
rect 51703 2816 51773 2862
rect 51819 2816 51889 2862
rect 51935 2816 52005 2862
rect 52051 2816 52121 2862
rect 52167 2816 52237 2862
rect 52283 2816 52353 2862
rect 52399 2816 52469 2862
rect 52515 2816 52585 2862
rect 52631 2816 52701 2862
rect 52747 2816 52817 2862
rect 52863 2816 52933 2862
rect 52979 2816 53049 2862
rect 53095 2816 53165 2862
rect 53211 2816 53281 2862
rect 53327 2816 53397 2862
rect 53443 2816 53513 2862
rect 53559 2816 53629 2862
rect 53675 2816 53745 2862
rect 53791 2816 53861 2862
rect 53907 2816 53977 2862
rect 54023 2816 54093 2862
rect 54139 2816 54209 2862
rect 54255 2816 54325 2862
rect 54371 2816 54441 2862
rect 54487 2816 54557 2862
rect 54603 2816 54673 2862
rect 54719 2816 54789 2862
rect 54835 2816 54905 2862
rect 54951 2816 55021 2862
rect 55067 2816 55137 2862
rect 55183 2816 55253 2862
rect 55299 2816 55369 2862
rect 55415 2816 55485 2862
rect 55531 2816 55601 2862
rect 55647 2816 55717 2862
rect 55763 2816 55833 2862
rect 55879 2816 55949 2862
rect 55995 2816 56065 2862
rect 56111 2816 56181 2862
rect 56227 2816 56297 2862
rect 56343 2816 56413 2862
rect 56459 2816 56529 2862
rect 56575 2816 56594 2862
rect 50826 2746 56594 2816
rect 50826 2700 50845 2746
rect 50891 2700 50961 2746
rect 51007 2700 51077 2746
rect 51123 2700 51193 2746
rect 51239 2700 51309 2746
rect 51355 2700 51425 2746
rect 51471 2700 51541 2746
rect 51587 2700 51657 2746
rect 51703 2700 51773 2746
rect 51819 2700 51889 2746
rect 51935 2700 52005 2746
rect 52051 2700 52121 2746
rect 52167 2700 52237 2746
rect 52283 2700 52353 2746
rect 52399 2700 52469 2746
rect 52515 2700 52585 2746
rect 52631 2700 52701 2746
rect 52747 2700 52817 2746
rect 52863 2700 52933 2746
rect 52979 2700 53049 2746
rect 53095 2700 53165 2746
rect 53211 2700 53281 2746
rect 53327 2700 53397 2746
rect 53443 2700 53513 2746
rect 53559 2700 53629 2746
rect 53675 2700 53745 2746
rect 53791 2700 53861 2746
rect 53907 2700 53977 2746
rect 54023 2700 54093 2746
rect 54139 2700 54209 2746
rect 54255 2700 54325 2746
rect 54371 2700 54441 2746
rect 54487 2700 54557 2746
rect 54603 2700 54673 2746
rect 54719 2700 54789 2746
rect 54835 2700 54905 2746
rect 54951 2700 55021 2746
rect 55067 2700 55137 2746
rect 55183 2700 55253 2746
rect 55299 2700 55369 2746
rect 55415 2700 55485 2746
rect 55531 2700 55601 2746
rect 55647 2700 55717 2746
rect 55763 2700 55833 2746
rect 55879 2700 55949 2746
rect 55995 2700 56065 2746
rect 56111 2700 56181 2746
rect 56227 2700 56297 2746
rect 56343 2700 56413 2746
rect 56459 2700 56529 2746
rect 56575 2700 56594 2746
rect 50826 2630 56594 2700
rect 50826 2584 50845 2630
rect 50891 2584 50961 2630
rect 51007 2584 51077 2630
rect 51123 2584 51193 2630
rect 51239 2584 51309 2630
rect 51355 2584 51425 2630
rect 51471 2584 51541 2630
rect 51587 2584 51657 2630
rect 51703 2584 51773 2630
rect 51819 2584 51889 2630
rect 51935 2584 52005 2630
rect 52051 2584 52121 2630
rect 52167 2584 52237 2630
rect 52283 2584 52353 2630
rect 52399 2584 52469 2630
rect 52515 2584 52585 2630
rect 52631 2584 52701 2630
rect 52747 2584 52817 2630
rect 52863 2584 52933 2630
rect 52979 2584 53049 2630
rect 53095 2584 53165 2630
rect 53211 2584 53281 2630
rect 53327 2584 53397 2630
rect 53443 2584 53513 2630
rect 53559 2584 53629 2630
rect 53675 2584 53745 2630
rect 53791 2584 53861 2630
rect 53907 2584 53977 2630
rect 54023 2584 54093 2630
rect 54139 2584 54209 2630
rect 54255 2584 54325 2630
rect 54371 2584 54441 2630
rect 54487 2584 54557 2630
rect 54603 2584 54673 2630
rect 54719 2584 54789 2630
rect 54835 2584 54905 2630
rect 54951 2584 55021 2630
rect 55067 2584 55137 2630
rect 55183 2584 55253 2630
rect 55299 2584 55369 2630
rect 55415 2584 55485 2630
rect 55531 2584 55601 2630
rect 55647 2584 55717 2630
rect 55763 2584 55833 2630
rect 55879 2584 55949 2630
rect 55995 2584 56065 2630
rect 56111 2584 56181 2630
rect 56227 2584 56297 2630
rect 56343 2584 56413 2630
rect 56459 2584 56529 2630
rect 56575 2584 56594 2630
rect 50826 2514 56594 2584
rect 50826 2468 50845 2514
rect 50891 2468 50961 2514
rect 51007 2468 51077 2514
rect 51123 2468 51193 2514
rect 51239 2468 51309 2514
rect 51355 2468 51425 2514
rect 51471 2468 51541 2514
rect 51587 2468 51657 2514
rect 51703 2468 51773 2514
rect 51819 2468 51889 2514
rect 51935 2468 52005 2514
rect 52051 2468 52121 2514
rect 52167 2468 52237 2514
rect 52283 2468 52353 2514
rect 52399 2468 52469 2514
rect 52515 2468 52585 2514
rect 52631 2468 52701 2514
rect 52747 2468 52817 2514
rect 52863 2468 52933 2514
rect 52979 2468 53049 2514
rect 53095 2468 53165 2514
rect 53211 2468 53281 2514
rect 53327 2468 53397 2514
rect 53443 2468 53513 2514
rect 53559 2468 53629 2514
rect 53675 2468 53745 2514
rect 53791 2468 53861 2514
rect 53907 2468 53977 2514
rect 54023 2468 54093 2514
rect 54139 2468 54209 2514
rect 54255 2468 54325 2514
rect 54371 2468 54441 2514
rect 54487 2468 54557 2514
rect 54603 2468 54673 2514
rect 54719 2468 54789 2514
rect 54835 2468 54905 2514
rect 54951 2468 55021 2514
rect 55067 2468 55137 2514
rect 55183 2468 55253 2514
rect 55299 2468 55369 2514
rect 55415 2468 55485 2514
rect 55531 2468 55601 2514
rect 55647 2468 55717 2514
rect 55763 2468 55833 2514
rect 55879 2468 55949 2514
rect 55995 2468 56065 2514
rect 56111 2468 56181 2514
rect 56227 2468 56297 2514
rect 56343 2468 56413 2514
rect 56459 2468 56529 2514
rect 56575 2468 56594 2514
rect 50826 2398 56594 2468
rect 50826 2352 50845 2398
rect 50891 2352 50961 2398
rect 51007 2352 51077 2398
rect 51123 2352 51193 2398
rect 51239 2352 51309 2398
rect 51355 2352 51425 2398
rect 51471 2352 51541 2398
rect 51587 2352 51657 2398
rect 51703 2352 51773 2398
rect 51819 2352 51889 2398
rect 51935 2352 52005 2398
rect 52051 2352 52121 2398
rect 52167 2352 52237 2398
rect 52283 2352 52353 2398
rect 52399 2352 52469 2398
rect 52515 2352 52585 2398
rect 52631 2352 52701 2398
rect 52747 2352 52817 2398
rect 52863 2352 52933 2398
rect 52979 2352 53049 2398
rect 53095 2352 53165 2398
rect 53211 2352 53281 2398
rect 53327 2352 53397 2398
rect 53443 2352 53513 2398
rect 53559 2352 53629 2398
rect 53675 2352 53745 2398
rect 53791 2352 53861 2398
rect 53907 2352 53977 2398
rect 54023 2352 54093 2398
rect 54139 2352 54209 2398
rect 54255 2352 54325 2398
rect 54371 2352 54441 2398
rect 54487 2352 54557 2398
rect 54603 2352 54673 2398
rect 54719 2352 54789 2398
rect 54835 2352 54905 2398
rect 54951 2352 55021 2398
rect 55067 2352 55137 2398
rect 55183 2352 55253 2398
rect 55299 2352 55369 2398
rect 55415 2352 55485 2398
rect 55531 2352 55601 2398
rect 55647 2352 55717 2398
rect 55763 2352 55833 2398
rect 55879 2352 55949 2398
rect 55995 2352 56065 2398
rect 56111 2352 56181 2398
rect 56227 2352 56297 2398
rect 56343 2352 56413 2398
rect 56459 2352 56529 2398
rect 56575 2352 56594 2398
rect 50826 2282 56594 2352
rect 50826 2236 50845 2282
rect 50891 2236 50961 2282
rect 51007 2236 51077 2282
rect 51123 2236 51193 2282
rect 51239 2236 51309 2282
rect 51355 2236 51425 2282
rect 51471 2236 51541 2282
rect 51587 2236 51657 2282
rect 51703 2236 51773 2282
rect 51819 2236 51889 2282
rect 51935 2236 52005 2282
rect 52051 2236 52121 2282
rect 52167 2236 52237 2282
rect 52283 2236 52353 2282
rect 52399 2236 52469 2282
rect 52515 2236 52585 2282
rect 52631 2236 52701 2282
rect 52747 2236 52817 2282
rect 52863 2236 52933 2282
rect 52979 2236 53049 2282
rect 53095 2236 53165 2282
rect 53211 2236 53281 2282
rect 53327 2236 53397 2282
rect 53443 2236 53513 2282
rect 53559 2236 53629 2282
rect 53675 2236 53745 2282
rect 53791 2236 53861 2282
rect 53907 2236 53977 2282
rect 54023 2236 54093 2282
rect 54139 2236 54209 2282
rect 54255 2236 54325 2282
rect 54371 2236 54441 2282
rect 54487 2236 54557 2282
rect 54603 2236 54673 2282
rect 54719 2236 54789 2282
rect 54835 2236 54905 2282
rect 54951 2236 55021 2282
rect 55067 2236 55137 2282
rect 55183 2236 55253 2282
rect 55299 2236 55369 2282
rect 55415 2236 55485 2282
rect 55531 2236 55601 2282
rect 55647 2236 55717 2282
rect 55763 2236 55833 2282
rect 55879 2236 55949 2282
rect 55995 2236 56065 2282
rect 56111 2236 56181 2282
rect 56227 2236 56297 2282
rect 56343 2236 56413 2282
rect 56459 2236 56529 2282
rect 56575 2236 56594 2282
rect 50826 2166 56594 2236
rect 50826 2120 50845 2166
rect 50891 2120 50961 2166
rect 51007 2120 51077 2166
rect 51123 2120 51193 2166
rect 51239 2120 51309 2166
rect 51355 2120 51425 2166
rect 51471 2120 51541 2166
rect 51587 2120 51657 2166
rect 51703 2120 51773 2166
rect 51819 2120 51889 2166
rect 51935 2120 52005 2166
rect 52051 2120 52121 2166
rect 52167 2120 52237 2166
rect 52283 2120 52353 2166
rect 52399 2120 52469 2166
rect 52515 2120 52585 2166
rect 52631 2120 52701 2166
rect 52747 2120 52817 2166
rect 52863 2120 52933 2166
rect 52979 2120 53049 2166
rect 53095 2120 53165 2166
rect 53211 2120 53281 2166
rect 53327 2120 53397 2166
rect 53443 2120 53513 2166
rect 53559 2120 53629 2166
rect 53675 2120 53745 2166
rect 53791 2120 53861 2166
rect 53907 2120 53977 2166
rect 54023 2120 54093 2166
rect 54139 2120 54209 2166
rect 54255 2120 54325 2166
rect 54371 2120 54441 2166
rect 54487 2120 54557 2166
rect 54603 2120 54673 2166
rect 54719 2120 54789 2166
rect 54835 2120 54905 2166
rect 54951 2120 55021 2166
rect 55067 2120 55137 2166
rect 55183 2120 55253 2166
rect 55299 2120 55369 2166
rect 55415 2120 55485 2166
rect 55531 2120 55601 2166
rect 55647 2120 55717 2166
rect 55763 2120 55833 2166
rect 55879 2120 55949 2166
rect 55995 2120 56065 2166
rect 56111 2120 56181 2166
rect 56227 2120 56297 2166
rect 56343 2120 56413 2166
rect 56459 2120 56529 2166
rect 56575 2120 56594 2166
rect 50826 2050 56594 2120
rect 50826 2004 50845 2050
rect 50891 2004 50961 2050
rect 51007 2004 51077 2050
rect 51123 2004 51193 2050
rect 51239 2004 51309 2050
rect 51355 2004 51425 2050
rect 51471 2004 51541 2050
rect 51587 2004 51657 2050
rect 51703 2004 51773 2050
rect 51819 2004 51889 2050
rect 51935 2004 52005 2050
rect 52051 2004 52121 2050
rect 52167 2004 52237 2050
rect 52283 2004 52353 2050
rect 52399 2004 52469 2050
rect 52515 2004 52585 2050
rect 52631 2004 52701 2050
rect 52747 2004 52817 2050
rect 52863 2004 52933 2050
rect 52979 2004 53049 2050
rect 53095 2004 53165 2050
rect 53211 2004 53281 2050
rect 53327 2004 53397 2050
rect 53443 2004 53513 2050
rect 53559 2004 53629 2050
rect 53675 2004 53745 2050
rect 53791 2004 53861 2050
rect 53907 2004 53977 2050
rect 54023 2004 54093 2050
rect 54139 2004 54209 2050
rect 54255 2004 54325 2050
rect 54371 2004 54441 2050
rect 54487 2004 54557 2050
rect 54603 2004 54673 2050
rect 54719 2004 54789 2050
rect 54835 2004 54905 2050
rect 54951 2004 55021 2050
rect 55067 2004 55137 2050
rect 55183 2004 55253 2050
rect 55299 2004 55369 2050
rect 55415 2004 55485 2050
rect 55531 2004 55601 2050
rect 55647 2004 55717 2050
rect 55763 2004 55833 2050
rect 55879 2004 55949 2050
rect 55995 2004 56065 2050
rect 56111 2004 56181 2050
rect 56227 2004 56297 2050
rect 56343 2004 56413 2050
rect 56459 2004 56529 2050
rect 56575 2004 56594 2050
rect 50826 1934 56594 2004
rect 50826 1888 50845 1934
rect 50891 1888 50961 1934
rect 51007 1888 51077 1934
rect 51123 1888 51193 1934
rect 51239 1888 51309 1934
rect 51355 1888 51425 1934
rect 51471 1888 51541 1934
rect 51587 1888 51657 1934
rect 51703 1888 51773 1934
rect 51819 1888 51889 1934
rect 51935 1888 52005 1934
rect 52051 1888 52121 1934
rect 52167 1888 52237 1934
rect 52283 1888 52353 1934
rect 52399 1888 52469 1934
rect 52515 1888 52585 1934
rect 52631 1888 52701 1934
rect 52747 1888 52817 1934
rect 52863 1888 52933 1934
rect 52979 1888 53049 1934
rect 53095 1888 53165 1934
rect 53211 1888 53281 1934
rect 53327 1888 53397 1934
rect 53443 1888 53513 1934
rect 53559 1888 53629 1934
rect 53675 1888 53745 1934
rect 53791 1888 53861 1934
rect 53907 1888 53977 1934
rect 54023 1888 54093 1934
rect 54139 1888 54209 1934
rect 54255 1888 54325 1934
rect 54371 1888 54441 1934
rect 54487 1888 54557 1934
rect 54603 1888 54673 1934
rect 54719 1888 54789 1934
rect 54835 1888 54905 1934
rect 54951 1888 55021 1934
rect 55067 1888 55137 1934
rect 55183 1888 55253 1934
rect 55299 1888 55369 1934
rect 55415 1888 55485 1934
rect 55531 1888 55601 1934
rect 55647 1888 55717 1934
rect 55763 1888 55833 1934
rect 55879 1888 55949 1934
rect 55995 1888 56065 1934
rect 56111 1888 56181 1934
rect 56227 1888 56297 1934
rect 56343 1888 56413 1934
rect 56459 1888 56529 1934
rect 56575 1888 56594 1934
rect 50826 1818 56594 1888
rect 50826 1772 50845 1818
rect 50891 1772 50961 1818
rect 51007 1772 51077 1818
rect 51123 1772 51193 1818
rect 51239 1772 51309 1818
rect 51355 1772 51425 1818
rect 51471 1772 51541 1818
rect 51587 1772 51657 1818
rect 51703 1772 51773 1818
rect 51819 1772 51889 1818
rect 51935 1772 52005 1818
rect 52051 1772 52121 1818
rect 52167 1772 52237 1818
rect 52283 1772 52353 1818
rect 52399 1772 52469 1818
rect 52515 1772 52585 1818
rect 52631 1772 52701 1818
rect 52747 1772 52817 1818
rect 52863 1772 52933 1818
rect 52979 1772 53049 1818
rect 53095 1772 53165 1818
rect 53211 1772 53281 1818
rect 53327 1772 53397 1818
rect 53443 1772 53513 1818
rect 53559 1772 53629 1818
rect 53675 1772 53745 1818
rect 53791 1772 53861 1818
rect 53907 1772 53977 1818
rect 54023 1772 54093 1818
rect 54139 1772 54209 1818
rect 54255 1772 54325 1818
rect 54371 1772 54441 1818
rect 54487 1772 54557 1818
rect 54603 1772 54673 1818
rect 54719 1772 54789 1818
rect 54835 1772 54905 1818
rect 54951 1772 55021 1818
rect 55067 1772 55137 1818
rect 55183 1772 55253 1818
rect 55299 1772 55369 1818
rect 55415 1772 55485 1818
rect 55531 1772 55601 1818
rect 55647 1772 55717 1818
rect 55763 1772 55833 1818
rect 55879 1772 55949 1818
rect 55995 1772 56065 1818
rect 56111 1772 56181 1818
rect 56227 1772 56297 1818
rect 56343 1772 56413 1818
rect 56459 1772 56529 1818
rect 56575 1772 56594 1818
rect 50826 1702 56594 1772
rect 50826 1656 50845 1702
rect 50891 1656 50961 1702
rect 51007 1656 51077 1702
rect 51123 1656 51193 1702
rect 51239 1656 51309 1702
rect 51355 1656 51425 1702
rect 51471 1656 51541 1702
rect 51587 1656 51657 1702
rect 51703 1656 51773 1702
rect 51819 1656 51889 1702
rect 51935 1656 52005 1702
rect 52051 1656 52121 1702
rect 52167 1656 52237 1702
rect 52283 1656 52353 1702
rect 52399 1656 52469 1702
rect 52515 1656 52585 1702
rect 52631 1656 52701 1702
rect 52747 1656 52817 1702
rect 52863 1656 52933 1702
rect 52979 1656 53049 1702
rect 53095 1656 53165 1702
rect 53211 1656 53281 1702
rect 53327 1656 53397 1702
rect 53443 1656 53513 1702
rect 53559 1656 53629 1702
rect 53675 1656 53745 1702
rect 53791 1656 53861 1702
rect 53907 1656 53977 1702
rect 54023 1656 54093 1702
rect 54139 1656 54209 1702
rect 54255 1656 54325 1702
rect 54371 1656 54441 1702
rect 54487 1656 54557 1702
rect 54603 1656 54673 1702
rect 54719 1656 54789 1702
rect 54835 1656 54905 1702
rect 54951 1656 55021 1702
rect 55067 1656 55137 1702
rect 55183 1656 55253 1702
rect 55299 1656 55369 1702
rect 55415 1656 55485 1702
rect 55531 1656 55601 1702
rect 55647 1656 55717 1702
rect 55763 1656 55833 1702
rect 55879 1656 55949 1702
rect 55995 1656 56065 1702
rect 56111 1656 56181 1702
rect 56227 1656 56297 1702
rect 56343 1656 56413 1702
rect 56459 1656 56529 1702
rect 56575 1656 56594 1702
rect 50826 1637 56594 1656
<< mvnsubdiff >>
rect 30583 65893 30802 65894
rect 30583 65836 32694 65893
rect 30583 65790 30854 65836
rect 30900 65790 31012 65836
rect 31058 65790 31170 65836
rect 31216 65790 31328 65836
rect 31374 65790 31487 65836
rect 31533 65790 31645 65836
rect 31691 65790 31803 65836
rect 31849 65790 31961 65836
rect 32007 65790 32119 65836
rect 32165 65790 32277 65836
rect 32323 65790 32435 65836
rect 32481 65790 32593 65836
rect 32639 65790 32694 65836
rect 30583 65722 32694 65790
rect 42662 65909 43608 65966
rect 42662 65863 42717 65909
rect 42763 65863 42875 65909
rect 42921 65863 43033 65909
rect 43079 65863 43191 65909
rect 43237 65863 43350 65909
rect 43396 65863 43508 65909
rect 43554 65863 43608 65909
rect 42662 65806 43608 65863
rect 30583 65676 30637 65722
rect 30683 65676 32694 65722
rect 30583 65673 32694 65676
rect 30583 65627 30854 65673
rect 30900 65627 31012 65673
rect 31058 65627 31170 65673
rect 31216 65627 31328 65673
rect 31374 65627 31487 65673
rect 31533 65627 31645 65673
rect 31691 65627 31803 65673
rect 31849 65627 31961 65673
rect 32007 65627 32119 65673
rect 32165 65627 32277 65673
rect 32323 65627 32435 65673
rect 32481 65627 32593 65673
rect 32639 65627 32694 65673
rect 30583 65558 32694 65627
rect 30583 65512 30637 65558
rect 30683 65512 32694 65558
rect 30583 65509 32694 65512
rect 30583 65463 30854 65509
rect 30900 65463 31012 65509
rect 31058 65463 31170 65509
rect 31216 65463 31328 65509
rect 31374 65463 31487 65509
rect 31533 65463 31645 65509
rect 31691 65463 31803 65509
rect 31849 65463 31961 65509
rect 32007 65463 32119 65509
rect 32165 65463 32277 65509
rect 32323 65463 32435 65509
rect 32481 65463 32593 65509
rect 32639 65463 32694 65509
rect 30583 65395 32694 65463
rect 54321 65893 54540 65894
rect 52428 65836 54540 65893
rect 52428 65790 52483 65836
rect 52529 65790 52641 65836
rect 52687 65790 52799 65836
rect 52845 65790 52957 65836
rect 53003 65790 53115 65836
rect 53161 65790 53273 65836
rect 53319 65790 53431 65836
rect 53477 65790 53589 65836
rect 53635 65790 53748 65836
rect 53794 65790 53906 65836
rect 53952 65790 54064 65836
rect 54110 65790 54222 65836
rect 54268 65790 54540 65836
rect 30583 65349 30637 65395
rect 30683 65349 32694 65395
rect 30583 65346 32694 65349
rect 30583 65300 30854 65346
rect 30900 65300 31012 65346
rect 31058 65300 31170 65346
rect 31216 65300 31328 65346
rect 31374 65300 31487 65346
rect 31533 65300 31645 65346
rect 31691 65300 31803 65346
rect 31849 65300 31961 65346
rect 32007 65300 32119 65346
rect 32165 65300 32277 65346
rect 32323 65300 32435 65346
rect 32481 65300 32593 65346
rect 32639 65300 32694 65346
rect 52428 65722 54540 65790
rect 52428 65676 54440 65722
rect 54486 65676 54540 65722
rect 52428 65673 54540 65676
rect 52428 65627 52483 65673
rect 52529 65627 52641 65673
rect 52687 65627 52799 65673
rect 52845 65627 52957 65673
rect 53003 65627 53115 65673
rect 53161 65627 53273 65673
rect 53319 65627 53431 65673
rect 53477 65627 53589 65673
rect 53635 65627 53748 65673
rect 53794 65627 53906 65673
rect 53952 65627 54064 65673
rect 54110 65627 54222 65673
rect 54268 65627 54540 65673
rect 52428 65558 54540 65627
rect 52428 65512 54440 65558
rect 54486 65512 54540 65558
rect 52428 65509 54540 65512
rect 52428 65463 52483 65509
rect 52529 65463 52641 65509
rect 52687 65463 52799 65509
rect 52845 65463 52957 65509
rect 53003 65463 53115 65509
rect 53161 65463 53273 65509
rect 53319 65463 53431 65509
rect 53477 65463 53589 65509
rect 53635 65463 53748 65509
rect 53794 65463 53906 65509
rect 53952 65463 54064 65509
rect 54110 65463 54222 65509
rect 54268 65463 54540 65509
rect 52428 65395 54540 65463
rect 52428 65349 54440 65395
rect 54486 65349 54540 65395
rect 52428 65346 54540 65349
rect 30583 65243 32694 65300
rect 52428 65300 52483 65346
rect 52529 65300 52641 65346
rect 52687 65300 52799 65346
rect 52845 65300 52957 65346
rect 53003 65300 53115 65346
rect 53161 65300 53273 65346
rect 53319 65300 53431 65346
rect 53477 65300 53589 65346
rect 53635 65300 53748 65346
rect 53794 65300 53906 65346
rect 53952 65300 54064 65346
rect 54110 65300 54222 65346
rect 54268 65300 54540 65346
rect 52428 65243 54540 65300
rect 30583 65232 30955 65243
rect 30583 65186 30637 65232
rect 30683 65186 30955 65232
rect 30583 65068 30955 65186
rect 30583 65022 30637 65068
rect 30683 65022 30955 65068
rect 30583 64989 30955 65022
rect 54167 65232 54540 65243
rect 54167 65186 54440 65232
rect 54486 65186 54540 65232
rect 54167 65068 54540 65186
rect 54167 65022 54440 65068
rect 54486 65022 54540 65068
rect 30583 64866 30956 64989
rect 36348 64950 36861 64996
rect 36348 64904 36489 64950
rect 36723 64904 36861 64950
rect 30583 64820 30637 64866
rect 30683 64826 30956 64866
rect 30683 64820 30855 64826
rect 30583 64780 30855 64820
rect 30901 64780 30956 64826
rect 30583 64703 30956 64780
rect 30583 64657 30637 64703
rect 30683 64662 30956 64703
rect 30683 64657 30855 64662
rect 30583 64616 30855 64657
rect 30901 64616 30956 64662
rect 30583 64540 30956 64616
rect 30583 64494 30637 64540
rect 30683 64499 30956 64540
rect 30683 64494 30855 64499
rect 30583 64453 30855 64494
rect 30901 64453 30956 64499
rect 30583 64377 30956 64453
rect 30583 64331 30637 64377
rect 30683 64336 30956 64377
rect 30683 64331 30855 64336
rect 30583 64290 30855 64331
rect 30901 64290 30956 64336
rect 36348 64858 36861 64904
rect 39007 64950 39321 65007
rect 39007 64904 39062 64950
rect 39108 64904 39220 64950
rect 39266 64904 39321 64950
rect 39007 64847 39321 64904
rect 45564 64996 48566 65007
rect 45564 64950 48766 64996
rect 54167 64987 54540 65022
rect 45564 64904 45619 64950
rect 45665 64904 45777 64950
rect 45823 64904 45935 64950
rect 45981 64904 46093 64950
rect 46139 64904 46251 64950
rect 46297 64904 46409 64950
rect 46455 64904 46568 64950
rect 46614 64904 46726 64950
rect 46772 64904 46884 64950
rect 46930 64904 47042 64950
rect 47088 64904 47200 64950
rect 47246 64904 47358 64950
rect 47404 64904 47516 64950
rect 47562 64904 47675 64950
rect 47721 64904 47833 64950
rect 47879 64904 47991 64950
rect 48037 64904 48149 64950
rect 48195 64904 48307 64950
rect 48353 64904 48465 64950
rect 48511 64904 48766 64950
rect 45564 64858 48766 64904
rect 45564 64786 48566 64858
rect 45564 64740 45619 64786
rect 45665 64740 45777 64786
rect 45823 64740 45935 64786
rect 45981 64740 46093 64786
rect 46139 64740 46251 64786
rect 46297 64740 46409 64786
rect 46455 64740 46568 64786
rect 46614 64740 46726 64786
rect 46772 64740 46884 64786
rect 46930 64740 47042 64786
rect 47088 64740 47200 64786
rect 47246 64740 47358 64786
rect 47404 64740 47516 64786
rect 47562 64740 47675 64786
rect 47721 64740 47833 64786
rect 47879 64740 47991 64786
rect 48037 64740 48149 64786
rect 48195 64740 48307 64786
rect 48353 64740 48465 64786
rect 48511 64740 48566 64786
rect 54168 64866 54540 64987
rect 54168 64826 54440 64866
rect 54168 64780 54223 64826
rect 54269 64820 54440 64826
rect 54486 64820 54540 64866
rect 54269 64780 54540 64820
rect 45564 64683 48566 64740
rect 30583 64213 30956 64290
rect 30583 64167 30637 64213
rect 30683 64173 30956 64213
rect 30683 64167 30855 64173
rect 30583 64127 30855 64167
rect 30901 64127 30956 64173
rect 54168 64703 54540 64780
rect 54168 64662 54440 64703
rect 54168 64616 54223 64662
rect 54269 64657 54440 64662
rect 54486 64657 54540 64703
rect 54269 64616 54540 64657
rect 54168 64540 54540 64616
rect 54168 64494 54440 64540
rect 54486 64494 54540 64540
rect 54168 64377 54540 64494
rect 54168 64331 54440 64377
rect 54486 64331 54540 64377
rect 54168 64213 54540 64331
rect 54168 64173 54440 64213
rect 30583 64050 30956 64127
rect 54168 64127 54223 64173
rect 54269 64167 54440 64173
rect 54486 64167 54540 64213
rect 54269 64127 54540 64167
rect 30583 64004 30637 64050
rect 30683 64004 30956 64050
rect 30583 63927 30956 64004
rect 54168 64050 54540 64127
rect 54168 64004 54440 64050
rect 54486 64004 54540 64050
rect 30583 63887 30855 63927
rect 30583 63841 30637 63887
rect 30683 63881 30855 63887
rect 30901 63881 30956 63927
rect 54168 63927 54540 64004
rect 30683 63841 30956 63881
rect 30583 63764 30956 63841
rect 30583 63723 30855 63764
rect 30583 63677 30637 63723
rect 30683 63718 30855 63723
rect 30901 63718 30956 63764
rect 30683 63677 30956 63718
rect 30583 63601 30956 63677
rect 30583 63560 30855 63601
rect 30583 63514 30637 63560
rect 30683 63555 30855 63560
rect 30901 63555 30956 63601
rect 30683 63514 30956 63555
rect 30583 63438 30956 63514
rect 30583 63397 30855 63438
rect 30583 63351 30637 63397
rect 30683 63392 30855 63397
rect 30901 63392 30956 63438
rect 30683 63351 30956 63392
rect 30583 63274 30956 63351
rect 30583 63234 30855 63274
rect 30583 63188 30637 63234
rect 30683 63228 30855 63234
rect 30901 63228 30956 63274
rect 30683 63188 30956 63228
rect 30583 63066 30956 63188
rect 54168 63881 54223 63927
rect 54269 63887 54540 63927
rect 54269 63881 54440 63887
rect 54168 63841 54440 63881
rect 54486 63841 54540 63887
rect 36348 63150 36861 63196
rect 36348 63104 36489 63150
rect 36723 63104 36861 63150
rect 30583 63020 30637 63066
rect 30683 63026 30956 63066
rect 30683 63020 30855 63026
rect 30583 62980 30855 63020
rect 30901 62980 30956 63026
rect 30583 62903 30956 62980
rect 30583 62857 30637 62903
rect 30683 62862 30956 62903
rect 30683 62857 30855 62862
rect 30583 62816 30855 62857
rect 30901 62816 30956 62862
rect 30583 62740 30956 62816
rect 30583 62694 30637 62740
rect 30683 62699 30956 62740
rect 30683 62694 30855 62699
rect 30583 62653 30855 62694
rect 30901 62653 30956 62699
rect 30583 62577 30956 62653
rect 30583 62531 30637 62577
rect 30683 62536 30956 62577
rect 30683 62531 30855 62536
rect 30583 62490 30855 62531
rect 30901 62490 30956 62536
rect 36348 63058 36861 63104
rect 39007 63150 39321 63207
rect 39007 63104 39062 63150
rect 39108 63104 39220 63150
rect 39266 63104 39321 63150
rect 39007 63047 39321 63104
rect 45564 63314 48566 63371
rect 45564 63268 45619 63314
rect 45665 63268 45777 63314
rect 45823 63268 45935 63314
rect 45981 63268 46093 63314
rect 46139 63268 46251 63314
rect 46297 63268 46409 63314
rect 46455 63268 46568 63314
rect 46614 63268 46726 63314
rect 46772 63268 46884 63314
rect 46930 63268 47042 63314
rect 47088 63268 47200 63314
rect 47246 63268 47358 63314
rect 47404 63268 47516 63314
rect 47562 63268 47675 63314
rect 47721 63268 47833 63314
rect 47879 63268 47991 63314
rect 48037 63268 48149 63314
rect 48195 63268 48307 63314
rect 48353 63268 48465 63314
rect 48511 63268 48566 63314
rect 54168 63723 54540 63841
rect 54168 63677 54440 63723
rect 54486 63677 54540 63723
rect 54168 63560 54540 63677
rect 54168 63514 54440 63560
rect 54486 63514 54540 63560
rect 54168 63438 54540 63514
rect 54168 63392 54223 63438
rect 54269 63397 54540 63438
rect 54269 63392 54440 63397
rect 54168 63351 54440 63392
rect 54486 63351 54540 63397
rect 45564 63196 48566 63268
rect 45564 63150 48766 63196
rect 54168 63274 54540 63351
rect 54168 63228 54223 63274
rect 54269 63234 54540 63274
rect 54269 63228 54440 63234
rect 54168 63188 54440 63228
rect 54486 63188 54540 63234
rect 45564 63104 45619 63150
rect 45665 63104 45777 63150
rect 45823 63104 45935 63150
rect 45981 63104 46093 63150
rect 46139 63104 46251 63150
rect 46297 63104 46409 63150
rect 46455 63104 46568 63150
rect 46614 63104 46726 63150
rect 46772 63104 46884 63150
rect 46930 63104 47042 63150
rect 47088 63104 47200 63150
rect 47246 63104 47358 63150
rect 47404 63104 47516 63150
rect 47562 63104 47675 63150
rect 47721 63104 47833 63150
rect 47879 63104 47991 63150
rect 48037 63104 48149 63150
rect 48195 63104 48307 63150
rect 48353 63104 48465 63150
rect 48511 63104 48766 63150
rect 45564 63058 48766 63104
rect 45564 62986 48566 63058
rect 45564 62940 45619 62986
rect 45665 62940 45777 62986
rect 45823 62940 45935 62986
rect 45981 62940 46093 62986
rect 46139 62940 46251 62986
rect 46297 62940 46409 62986
rect 46455 62940 46568 62986
rect 46614 62940 46726 62986
rect 46772 62940 46884 62986
rect 46930 62940 47042 62986
rect 47088 62940 47200 62986
rect 47246 62940 47358 62986
rect 47404 62940 47516 62986
rect 47562 62940 47675 62986
rect 47721 62940 47833 62986
rect 47879 62940 47991 62986
rect 48037 62940 48149 62986
rect 48195 62940 48307 62986
rect 48353 62940 48465 62986
rect 48511 62940 48566 62986
rect 54168 63066 54540 63188
rect 54168 63026 54440 63066
rect 54168 62980 54223 63026
rect 54269 63020 54440 63026
rect 54486 63020 54540 63066
rect 54269 62980 54540 63020
rect 45564 62883 48566 62940
rect 30583 62413 30956 62490
rect 30583 62367 30637 62413
rect 30683 62373 30956 62413
rect 30683 62367 30855 62373
rect 30583 62327 30855 62367
rect 30901 62327 30956 62373
rect 54168 62903 54540 62980
rect 54168 62862 54440 62903
rect 54168 62816 54223 62862
rect 54269 62857 54440 62862
rect 54486 62857 54540 62903
rect 54269 62816 54540 62857
rect 54168 62740 54540 62816
rect 54168 62694 54440 62740
rect 54486 62694 54540 62740
rect 54168 62577 54540 62694
rect 54168 62531 54440 62577
rect 54486 62531 54540 62577
rect 54168 62413 54540 62531
rect 54168 62373 54440 62413
rect 30583 62250 30956 62327
rect 54168 62327 54223 62373
rect 54269 62367 54440 62373
rect 54486 62367 54540 62413
rect 54269 62327 54540 62367
rect 30583 62204 30637 62250
rect 30683 62204 30956 62250
rect 30583 62127 30956 62204
rect 54168 62250 54540 62327
rect 54168 62204 54440 62250
rect 54486 62204 54540 62250
rect 30583 62087 30855 62127
rect 30583 62041 30637 62087
rect 30683 62081 30855 62087
rect 30901 62081 30956 62127
rect 54168 62127 54540 62204
rect 30683 62041 30956 62081
rect 30583 61964 30956 62041
rect 30583 61923 30855 61964
rect 30583 61877 30637 61923
rect 30683 61918 30855 61923
rect 30901 61918 30956 61964
rect 30683 61877 30956 61918
rect 30583 61801 30956 61877
rect 30583 61760 30855 61801
rect 30583 61714 30637 61760
rect 30683 61755 30855 61760
rect 30901 61755 30956 61801
rect 30683 61714 30956 61755
rect 30583 61638 30956 61714
rect 30583 61597 30855 61638
rect 30583 61551 30637 61597
rect 30683 61592 30855 61597
rect 30901 61592 30956 61638
rect 30683 61551 30956 61592
rect 30583 61474 30956 61551
rect 30583 61434 30855 61474
rect 30583 61388 30637 61434
rect 30683 61428 30855 61434
rect 30901 61428 30956 61474
rect 30683 61388 30956 61428
rect 30583 61266 30956 61388
rect 54168 62081 54223 62127
rect 54269 62087 54540 62127
rect 54269 62081 54440 62087
rect 54168 62041 54440 62081
rect 54486 62041 54540 62087
rect 36348 61350 36861 61396
rect 36348 61304 36489 61350
rect 36723 61304 36861 61350
rect 30583 61220 30637 61266
rect 30683 61226 30956 61266
rect 30683 61220 30855 61226
rect 30583 61180 30855 61220
rect 30901 61180 30956 61226
rect 30583 61103 30956 61180
rect 30583 61057 30637 61103
rect 30683 61062 30956 61103
rect 30683 61057 30855 61062
rect 30583 61016 30855 61057
rect 30901 61016 30956 61062
rect 30583 60940 30956 61016
rect 30583 60894 30637 60940
rect 30683 60899 30956 60940
rect 30683 60894 30855 60899
rect 30583 60853 30855 60894
rect 30901 60853 30956 60899
rect 30583 60777 30956 60853
rect 30583 60731 30637 60777
rect 30683 60736 30956 60777
rect 30683 60731 30855 60736
rect 30583 60690 30855 60731
rect 30901 60690 30956 60736
rect 36348 61258 36861 61304
rect 39007 61350 39321 61407
rect 39007 61304 39062 61350
rect 39108 61304 39220 61350
rect 39266 61304 39321 61350
rect 39007 61247 39321 61304
rect 45564 61514 48566 61571
rect 45564 61468 45619 61514
rect 45665 61468 45777 61514
rect 45823 61468 45935 61514
rect 45981 61468 46093 61514
rect 46139 61468 46251 61514
rect 46297 61468 46409 61514
rect 46455 61468 46568 61514
rect 46614 61468 46726 61514
rect 46772 61468 46884 61514
rect 46930 61468 47042 61514
rect 47088 61468 47200 61514
rect 47246 61468 47358 61514
rect 47404 61468 47516 61514
rect 47562 61468 47675 61514
rect 47721 61468 47833 61514
rect 47879 61468 47991 61514
rect 48037 61468 48149 61514
rect 48195 61468 48307 61514
rect 48353 61468 48465 61514
rect 48511 61468 48566 61514
rect 54168 61923 54540 62041
rect 54168 61877 54440 61923
rect 54486 61877 54540 61923
rect 54168 61760 54540 61877
rect 54168 61714 54440 61760
rect 54486 61714 54540 61760
rect 54168 61638 54540 61714
rect 54168 61592 54223 61638
rect 54269 61597 54540 61638
rect 54269 61592 54440 61597
rect 54168 61551 54440 61592
rect 54486 61551 54540 61597
rect 45564 61396 48566 61468
rect 45564 61350 48766 61396
rect 54168 61474 54540 61551
rect 54168 61428 54223 61474
rect 54269 61434 54540 61474
rect 54269 61428 54440 61434
rect 54168 61388 54440 61428
rect 54486 61388 54540 61434
rect 45564 61304 45619 61350
rect 45665 61304 45777 61350
rect 45823 61304 45935 61350
rect 45981 61304 46093 61350
rect 46139 61304 46251 61350
rect 46297 61304 46409 61350
rect 46455 61304 46568 61350
rect 46614 61304 46726 61350
rect 46772 61304 46884 61350
rect 46930 61304 47042 61350
rect 47088 61304 47200 61350
rect 47246 61304 47358 61350
rect 47404 61304 47516 61350
rect 47562 61304 47675 61350
rect 47721 61304 47833 61350
rect 47879 61304 47991 61350
rect 48037 61304 48149 61350
rect 48195 61304 48307 61350
rect 48353 61304 48465 61350
rect 48511 61304 48766 61350
rect 45564 61258 48766 61304
rect 45564 61186 48566 61258
rect 45564 61140 45619 61186
rect 45665 61140 45777 61186
rect 45823 61140 45935 61186
rect 45981 61140 46093 61186
rect 46139 61140 46251 61186
rect 46297 61140 46409 61186
rect 46455 61140 46568 61186
rect 46614 61140 46726 61186
rect 46772 61140 46884 61186
rect 46930 61140 47042 61186
rect 47088 61140 47200 61186
rect 47246 61140 47358 61186
rect 47404 61140 47516 61186
rect 47562 61140 47675 61186
rect 47721 61140 47833 61186
rect 47879 61140 47991 61186
rect 48037 61140 48149 61186
rect 48195 61140 48307 61186
rect 48353 61140 48465 61186
rect 48511 61140 48566 61186
rect 54168 61266 54540 61388
rect 54168 61226 54440 61266
rect 54168 61180 54223 61226
rect 54269 61220 54440 61226
rect 54486 61220 54540 61266
rect 54269 61180 54540 61220
rect 45564 61083 48566 61140
rect 30583 60613 30956 60690
rect 30583 60567 30637 60613
rect 30683 60573 30956 60613
rect 30683 60567 30855 60573
rect 30583 60527 30855 60567
rect 30901 60527 30956 60573
rect 54168 61103 54540 61180
rect 54168 61062 54440 61103
rect 54168 61016 54223 61062
rect 54269 61057 54440 61062
rect 54486 61057 54540 61103
rect 54269 61016 54540 61057
rect 54168 60940 54540 61016
rect 54168 60894 54440 60940
rect 54486 60894 54540 60940
rect 54168 60777 54540 60894
rect 54168 60731 54440 60777
rect 54486 60731 54540 60777
rect 54168 60613 54540 60731
rect 54168 60573 54440 60613
rect 30583 60450 30956 60527
rect 54168 60527 54223 60573
rect 54269 60567 54440 60573
rect 54486 60567 54540 60613
rect 54269 60527 54540 60567
rect 30583 60404 30637 60450
rect 30683 60404 30956 60450
rect 30583 60327 30956 60404
rect 54168 60450 54540 60527
rect 54168 60404 54440 60450
rect 54486 60404 54540 60450
rect 30583 60287 30855 60327
rect 30583 60241 30637 60287
rect 30683 60281 30855 60287
rect 30901 60281 30956 60327
rect 54168 60327 54540 60404
rect 30683 60241 30956 60281
rect 30583 60164 30956 60241
rect 30583 60123 30855 60164
rect 30583 60077 30637 60123
rect 30683 60118 30855 60123
rect 30901 60118 30956 60164
rect 30683 60077 30956 60118
rect 30583 60001 30956 60077
rect 30583 59960 30855 60001
rect 30583 59914 30637 59960
rect 30683 59955 30855 59960
rect 30901 59955 30956 60001
rect 30683 59914 30956 59955
rect 30583 59838 30956 59914
rect 30583 59797 30855 59838
rect 30583 59751 30637 59797
rect 30683 59792 30855 59797
rect 30901 59792 30956 59838
rect 30683 59751 30956 59792
rect 30583 59674 30956 59751
rect 30583 59634 30855 59674
rect 30583 59588 30637 59634
rect 30683 59628 30855 59634
rect 30901 59628 30956 59674
rect 30683 59588 30956 59628
rect 30583 59466 30956 59588
rect 54168 60281 54223 60327
rect 54269 60287 54540 60327
rect 54269 60281 54440 60287
rect 54168 60241 54440 60281
rect 54486 60241 54540 60287
rect 36348 59550 36861 59596
rect 36348 59504 36489 59550
rect 36723 59504 36861 59550
rect 30583 59420 30637 59466
rect 30683 59426 30956 59466
rect 30683 59420 30855 59426
rect 30583 59380 30855 59420
rect 30901 59380 30956 59426
rect 30583 59303 30956 59380
rect 30583 59257 30637 59303
rect 30683 59262 30956 59303
rect 30683 59257 30855 59262
rect 30583 59216 30855 59257
rect 30901 59216 30956 59262
rect 30583 59140 30956 59216
rect 30583 59094 30637 59140
rect 30683 59099 30956 59140
rect 30683 59094 30855 59099
rect 30583 59053 30855 59094
rect 30901 59053 30956 59099
rect 30583 58977 30956 59053
rect 30583 58931 30637 58977
rect 30683 58936 30956 58977
rect 30683 58931 30855 58936
rect 30583 58890 30855 58931
rect 30901 58890 30956 58936
rect 36348 59458 36861 59504
rect 39007 59550 39321 59607
rect 39007 59504 39062 59550
rect 39108 59504 39220 59550
rect 39266 59504 39321 59550
rect 39007 59447 39321 59504
rect 45564 59714 48566 59771
rect 45564 59668 45619 59714
rect 45665 59668 45777 59714
rect 45823 59668 45935 59714
rect 45981 59668 46093 59714
rect 46139 59668 46251 59714
rect 46297 59668 46409 59714
rect 46455 59668 46568 59714
rect 46614 59668 46726 59714
rect 46772 59668 46884 59714
rect 46930 59668 47042 59714
rect 47088 59668 47200 59714
rect 47246 59668 47358 59714
rect 47404 59668 47516 59714
rect 47562 59668 47675 59714
rect 47721 59668 47833 59714
rect 47879 59668 47991 59714
rect 48037 59668 48149 59714
rect 48195 59668 48307 59714
rect 48353 59668 48465 59714
rect 48511 59668 48566 59714
rect 54168 60123 54540 60241
rect 54168 60077 54440 60123
rect 54486 60077 54540 60123
rect 54168 59960 54540 60077
rect 54168 59914 54440 59960
rect 54486 59914 54540 59960
rect 54168 59838 54540 59914
rect 54168 59792 54223 59838
rect 54269 59797 54540 59838
rect 54269 59792 54440 59797
rect 54168 59751 54440 59792
rect 54486 59751 54540 59797
rect 45564 59596 48566 59668
rect 45564 59550 48766 59596
rect 54168 59674 54540 59751
rect 54168 59628 54223 59674
rect 54269 59634 54540 59674
rect 54269 59628 54440 59634
rect 54168 59588 54440 59628
rect 54486 59588 54540 59634
rect 45564 59504 45619 59550
rect 45665 59504 45777 59550
rect 45823 59504 45935 59550
rect 45981 59504 46093 59550
rect 46139 59504 46251 59550
rect 46297 59504 46409 59550
rect 46455 59504 46568 59550
rect 46614 59504 46726 59550
rect 46772 59504 46884 59550
rect 46930 59504 47042 59550
rect 47088 59504 47200 59550
rect 47246 59504 47358 59550
rect 47404 59504 47516 59550
rect 47562 59504 47675 59550
rect 47721 59504 47833 59550
rect 47879 59504 47991 59550
rect 48037 59504 48149 59550
rect 48195 59504 48307 59550
rect 48353 59504 48465 59550
rect 48511 59504 48766 59550
rect 45564 59458 48766 59504
rect 45564 59386 48566 59458
rect 45564 59340 45619 59386
rect 45665 59340 45777 59386
rect 45823 59340 45935 59386
rect 45981 59340 46093 59386
rect 46139 59340 46251 59386
rect 46297 59340 46409 59386
rect 46455 59340 46568 59386
rect 46614 59340 46726 59386
rect 46772 59340 46884 59386
rect 46930 59340 47042 59386
rect 47088 59340 47200 59386
rect 47246 59340 47358 59386
rect 47404 59340 47516 59386
rect 47562 59340 47675 59386
rect 47721 59340 47833 59386
rect 47879 59340 47991 59386
rect 48037 59340 48149 59386
rect 48195 59340 48307 59386
rect 48353 59340 48465 59386
rect 48511 59340 48566 59386
rect 54168 59466 54540 59588
rect 54168 59426 54440 59466
rect 54168 59380 54223 59426
rect 54269 59420 54440 59426
rect 54486 59420 54540 59466
rect 54269 59380 54540 59420
rect 45564 59283 48566 59340
rect 30583 58813 30956 58890
rect 30583 58767 30637 58813
rect 30683 58773 30956 58813
rect 30683 58767 30855 58773
rect 30583 58727 30855 58767
rect 30901 58727 30956 58773
rect 54168 59303 54540 59380
rect 54168 59262 54440 59303
rect 54168 59216 54223 59262
rect 54269 59257 54440 59262
rect 54486 59257 54540 59303
rect 54269 59216 54540 59257
rect 54168 59140 54540 59216
rect 54168 59094 54440 59140
rect 54486 59094 54540 59140
rect 54168 58977 54540 59094
rect 54168 58931 54440 58977
rect 54486 58931 54540 58977
rect 54168 58813 54540 58931
rect 54168 58773 54440 58813
rect 30583 58650 30956 58727
rect 54168 58727 54223 58773
rect 54269 58767 54440 58773
rect 54486 58767 54540 58813
rect 54269 58727 54540 58767
rect 30583 58604 30637 58650
rect 30683 58604 30956 58650
rect 30583 58527 30956 58604
rect 54168 58650 54540 58727
rect 54168 58604 54440 58650
rect 54486 58604 54540 58650
rect 30583 58487 30855 58527
rect 30583 58441 30637 58487
rect 30683 58481 30855 58487
rect 30901 58481 30956 58527
rect 54168 58527 54540 58604
rect 30683 58441 30956 58481
rect 30583 58364 30956 58441
rect 30583 58323 30855 58364
rect 30583 58277 30637 58323
rect 30683 58318 30855 58323
rect 30901 58318 30956 58364
rect 30683 58277 30956 58318
rect 30583 58201 30956 58277
rect 30583 58160 30855 58201
rect 30583 58114 30637 58160
rect 30683 58155 30855 58160
rect 30901 58155 30956 58201
rect 30683 58114 30956 58155
rect 30583 58038 30956 58114
rect 30583 57997 30855 58038
rect 30583 57951 30637 57997
rect 30683 57992 30855 57997
rect 30901 57992 30956 58038
rect 30683 57951 30956 57992
rect 30583 57874 30956 57951
rect 30583 57834 30855 57874
rect 30583 57788 30637 57834
rect 30683 57828 30855 57834
rect 30901 57828 30956 57874
rect 30683 57788 30956 57828
rect 30583 57666 30956 57788
rect 54168 58481 54223 58527
rect 54269 58487 54540 58527
rect 54269 58481 54440 58487
rect 54168 58441 54440 58481
rect 54486 58441 54540 58487
rect 36348 57750 36861 57796
rect 36348 57704 36489 57750
rect 36723 57704 36861 57750
rect 30583 57620 30637 57666
rect 30683 57626 30956 57666
rect 30683 57620 30855 57626
rect 30583 57580 30855 57620
rect 30901 57580 30956 57626
rect 30583 57503 30956 57580
rect 30583 57457 30637 57503
rect 30683 57462 30956 57503
rect 30683 57457 30855 57462
rect 30583 57416 30855 57457
rect 30901 57416 30956 57462
rect 30583 57340 30956 57416
rect 30583 57294 30637 57340
rect 30683 57299 30956 57340
rect 30683 57294 30855 57299
rect 30583 57253 30855 57294
rect 30901 57253 30956 57299
rect 30583 57177 30956 57253
rect 30583 57131 30637 57177
rect 30683 57136 30956 57177
rect 30683 57131 30855 57136
rect 30583 57090 30855 57131
rect 30901 57090 30956 57136
rect 36348 57658 36861 57704
rect 39007 57750 39321 57807
rect 39007 57704 39062 57750
rect 39108 57704 39220 57750
rect 39266 57704 39321 57750
rect 39007 57647 39321 57704
rect 45564 57914 48566 57971
rect 45564 57868 45619 57914
rect 45665 57868 45777 57914
rect 45823 57868 45935 57914
rect 45981 57868 46093 57914
rect 46139 57868 46251 57914
rect 46297 57868 46409 57914
rect 46455 57868 46568 57914
rect 46614 57868 46726 57914
rect 46772 57868 46884 57914
rect 46930 57868 47042 57914
rect 47088 57868 47200 57914
rect 47246 57868 47358 57914
rect 47404 57868 47516 57914
rect 47562 57868 47675 57914
rect 47721 57868 47833 57914
rect 47879 57868 47991 57914
rect 48037 57868 48149 57914
rect 48195 57868 48307 57914
rect 48353 57868 48465 57914
rect 48511 57868 48566 57914
rect 54168 58323 54540 58441
rect 54168 58277 54440 58323
rect 54486 58277 54540 58323
rect 54168 58160 54540 58277
rect 54168 58114 54440 58160
rect 54486 58114 54540 58160
rect 54168 58038 54540 58114
rect 54168 57992 54223 58038
rect 54269 57997 54540 58038
rect 54269 57992 54440 57997
rect 54168 57951 54440 57992
rect 54486 57951 54540 57997
rect 45564 57796 48566 57868
rect 45564 57750 48766 57796
rect 54168 57874 54540 57951
rect 54168 57828 54223 57874
rect 54269 57834 54540 57874
rect 54269 57828 54440 57834
rect 54168 57788 54440 57828
rect 54486 57788 54540 57834
rect 45564 57704 45619 57750
rect 45665 57704 45777 57750
rect 45823 57704 45935 57750
rect 45981 57704 46093 57750
rect 46139 57704 46251 57750
rect 46297 57704 46409 57750
rect 46455 57704 46568 57750
rect 46614 57704 46726 57750
rect 46772 57704 46884 57750
rect 46930 57704 47042 57750
rect 47088 57704 47200 57750
rect 47246 57704 47358 57750
rect 47404 57704 47516 57750
rect 47562 57704 47675 57750
rect 47721 57704 47833 57750
rect 47879 57704 47991 57750
rect 48037 57704 48149 57750
rect 48195 57704 48307 57750
rect 48353 57704 48465 57750
rect 48511 57704 48766 57750
rect 45564 57658 48766 57704
rect 45564 57586 48566 57658
rect 45564 57540 45619 57586
rect 45665 57540 45777 57586
rect 45823 57540 45935 57586
rect 45981 57540 46093 57586
rect 46139 57540 46251 57586
rect 46297 57540 46409 57586
rect 46455 57540 46568 57586
rect 46614 57540 46726 57586
rect 46772 57540 46884 57586
rect 46930 57540 47042 57586
rect 47088 57540 47200 57586
rect 47246 57540 47358 57586
rect 47404 57540 47516 57586
rect 47562 57540 47675 57586
rect 47721 57540 47833 57586
rect 47879 57540 47991 57586
rect 48037 57540 48149 57586
rect 48195 57540 48307 57586
rect 48353 57540 48465 57586
rect 48511 57540 48566 57586
rect 54168 57666 54540 57788
rect 54168 57626 54440 57666
rect 54168 57580 54223 57626
rect 54269 57620 54440 57626
rect 54486 57620 54540 57666
rect 54269 57580 54540 57620
rect 45564 57483 48566 57540
rect 30583 57013 30956 57090
rect 30583 56967 30637 57013
rect 30683 56973 30956 57013
rect 30683 56967 30855 56973
rect 30583 56927 30855 56967
rect 30901 56927 30956 56973
rect 54168 57503 54540 57580
rect 54168 57462 54440 57503
rect 54168 57416 54223 57462
rect 54269 57457 54440 57462
rect 54486 57457 54540 57503
rect 54269 57416 54540 57457
rect 54168 57340 54540 57416
rect 54168 57294 54440 57340
rect 54486 57294 54540 57340
rect 54168 57177 54540 57294
rect 54168 57131 54440 57177
rect 54486 57131 54540 57177
rect 54168 57013 54540 57131
rect 54168 56973 54440 57013
rect 30583 56850 30956 56927
rect 54168 56927 54223 56973
rect 54269 56967 54440 56973
rect 54486 56967 54540 57013
rect 54269 56927 54540 56967
rect 30583 56804 30637 56850
rect 30683 56804 30956 56850
rect 30583 56727 30956 56804
rect 54168 56850 54540 56927
rect 54168 56804 54440 56850
rect 54486 56804 54540 56850
rect 30583 56687 30855 56727
rect 30583 56641 30637 56687
rect 30683 56681 30855 56687
rect 30901 56681 30956 56727
rect 54168 56727 54540 56804
rect 30683 56641 30956 56681
rect 30583 56564 30956 56641
rect 30583 56523 30855 56564
rect 30583 56477 30637 56523
rect 30683 56518 30855 56523
rect 30901 56518 30956 56564
rect 30683 56477 30956 56518
rect 30583 56401 30956 56477
rect 30583 56360 30855 56401
rect 30583 56314 30637 56360
rect 30683 56355 30855 56360
rect 30901 56355 30956 56401
rect 30683 56314 30956 56355
rect 30583 56238 30956 56314
rect 30583 56197 30855 56238
rect 30583 56151 30637 56197
rect 30683 56192 30855 56197
rect 30901 56192 30956 56238
rect 30683 56151 30956 56192
rect 30583 56074 30956 56151
rect 30583 56034 30855 56074
rect 30583 55988 30637 56034
rect 30683 56028 30855 56034
rect 30901 56028 30956 56074
rect 30683 55988 30956 56028
rect 30583 55866 30956 55988
rect 54168 56681 54223 56727
rect 54269 56687 54540 56727
rect 54269 56681 54440 56687
rect 54168 56641 54440 56681
rect 54486 56641 54540 56687
rect 36348 55950 36861 55996
rect 36348 55904 36489 55950
rect 36723 55904 36861 55950
rect 30583 55820 30637 55866
rect 30683 55826 30956 55866
rect 30683 55820 30855 55826
rect 30583 55780 30855 55820
rect 30901 55780 30956 55826
rect 30583 55703 30956 55780
rect 30583 55657 30637 55703
rect 30683 55662 30956 55703
rect 30683 55657 30855 55662
rect 30583 55616 30855 55657
rect 30901 55616 30956 55662
rect 30583 55540 30956 55616
rect 30583 55494 30637 55540
rect 30683 55499 30956 55540
rect 30683 55494 30855 55499
rect 30583 55453 30855 55494
rect 30901 55453 30956 55499
rect 30583 55377 30956 55453
rect 30583 55331 30637 55377
rect 30683 55336 30956 55377
rect 30683 55331 30855 55336
rect 30583 55290 30855 55331
rect 30901 55290 30956 55336
rect 36348 55858 36861 55904
rect 39007 55950 39321 56007
rect 39007 55904 39062 55950
rect 39108 55904 39220 55950
rect 39266 55904 39321 55950
rect 39007 55847 39321 55904
rect 45564 56114 48566 56171
rect 45564 56068 45619 56114
rect 45665 56068 45777 56114
rect 45823 56068 45935 56114
rect 45981 56068 46093 56114
rect 46139 56068 46251 56114
rect 46297 56068 46409 56114
rect 46455 56068 46568 56114
rect 46614 56068 46726 56114
rect 46772 56068 46884 56114
rect 46930 56068 47042 56114
rect 47088 56068 47200 56114
rect 47246 56068 47358 56114
rect 47404 56068 47516 56114
rect 47562 56068 47675 56114
rect 47721 56068 47833 56114
rect 47879 56068 47991 56114
rect 48037 56068 48149 56114
rect 48195 56068 48307 56114
rect 48353 56068 48465 56114
rect 48511 56068 48566 56114
rect 54168 56523 54540 56641
rect 54168 56477 54440 56523
rect 54486 56477 54540 56523
rect 54168 56360 54540 56477
rect 54168 56314 54440 56360
rect 54486 56314 54540 56360
rect 54168 56238 54540 56314
rect 54168 56192 54223 56238
rect 54269 56197 54540 56238
rect 54269 56192 54440 56197
rect 54168 56151 54440 56192
rect 54486 56151 54540 56197
rect 45564 55996 48566 56068
rect 45564 55950 48766 55996
rect 54168 56074 54540 56151
rect 54168 56028 54223 56074
rect 54269 56034 54540 56074
rect 54269 56028 54440 56034
rect 54168 55988 54440 56028
rect 54486 55988 54540 56034
rect 45564 55904 45619 55950
rect 45665 55904 45777 55950
rect 45823 55904 45935 55950
rect 45981 55904 46093 55950
rect 46139 55904 46251 55950
rect 46297 55904 46409 55950
rect 46455 55904 46568 55950
rect 46614 55904 46726 55950
rect 46772 55904 46884 55950
rect 46930 55904 47042 55950
rect 47088 55904 47200 55950
rect 47246 55904 47358 55950
rect 47404 55904 47516 55950
rect 47562 55904 47675 55950
rect 47721 55904 47833 55950
rect 47879 55904 47991 55950
rect 48037 55904 48149 55950
rect 48195 55904 48307 55950
rect 48353 55904 48465 55950
rect 48511 55904 48766 55950
rect 45564 55858 48766 55904
rect 45564 55786 48566 55858
rect 45564 55740 45619 55786
rect 45665 55740 45777 55786
rect 45823 55740 45935 55786
rect 45981 55740 46093 55786
rect 46139 55740 46251 55786
rect 46297 55740 46409 55786
rect 46455 55740 46568 55786
rect 46614 55740 46726 55786
rect 46772 55740 46884 55786
rect 46930 55740 47042 55786
rect 47088 55740 47200 55786
rect 47246 55740 47358 55786
rect 47404 55740 47516 55786
rect 47562 55740 47675 55786
rect 47721 55740 47833 55786
rect 47879 55740 47991 55786
rect 48037 55740 48149 55786
rect 48195 55740 48307 55786
rect 48353 55740 48465 55786
rect 48511 55740 48566 55786
rect 54168 55866 54540 55988
rect 54168 55826 54440 55866
rect 54168 55780 54223 55826
rect 54269 55820 54440 55826
rect 54486 55820 54540 55866
rect 54269 55780 54540 55820
rect 45564 55683 48566 55740
rect 30583 55213 30956 55290
rect 30583 55167 30637 55213
rect 30683 55173 30956 55213
rect 30683 55167 30855 55173
rect 30583 55127 30855 55167
rect 30901 55127 30956 55173
rect 54168 55703 54540 55780
rect 54168 55662 54440 55703
rect 54168 55616 54223 55662
rect 54269 55657 54440 55662
rect 54486 55657 54540 55703
rect 54269 55616 54540 55657
rect 54168 55540 54540 55616
rect 54168 55494 54440 55540
rect 54486 55494 54540 55540
rect 54168 55377 54540 55494
rect 54168 55331 54440 55377
rect 54486 55331 54540 55377
rect 54168 55213 54540 55331
rect 54168 55173 54440 55213
rect 30583 55050 30956 55127
rect 54168 55127 54223 55173
rect 54269 55167 54440 55173
rect 54486 55167 54540 55213
rect 54269 55127 54540 55167
rect 30583 55004 30637 55050
rect 30683 55004 30956 55050
rect 30583 54927 30956 55004
rect 54168 55050 54540 55127
rect 54168 55004 54440 55050
rect 54486 55004 54540 55050
rect 30583 54887 30855 54927
rect 30583 54841 30637 54887
rect 30683 54881 30855 54887
rect 30901 54881 30956 54927
rect 54168 54927 54540 55004
rect 30683 54841 30956 54881
rect 30583 54764 30956 54841
rect 30583 54723 30855 54764
rect 30583 54677 30637 54723
rect 30683 54718 30855 54723
rect 30901 54718 30956 54764
rect 30683 54677 30956 54718
rect 30583 54601 30956 54677
rect 30583 54560 30855 54601
rect 30583 54514 30637 54560
rect 30683 54555 30855 54560
rect 30901 54555 30956 54601
rect 30683 54514 30956 54555
rect 30583 54438 30956 54514
rect 30583 54397 30855 54438
rect 30583 54351 30637 54397
rect 30683 54392 30855 54397
rect 30901 54392 30956 54438
rect 30683 54351 30956 54392
rect 30583 54274 30956 54351
rect 30583 54234 30855 54274
rect 30583 54188 30637 54234
rect 30683 54228 30855 54234
rect 30901 54228 30956 54274
rect 30683 54188 30956 54228
rect 30583 54066 30956 54188
rect 54168 54881 54223 54927
rect 54269 54887 54540 54927
rect 54269 54881 54440 54887
rect 54168 54841 54440 54881
rect 54486 54841 54540 54887
rect 36348 54150 36861 54196
rect 36348 54104 36489 54150
rect 36723 54104 36861 54150
rect 30583 54020 30637 54066
rect 30683 54026 30956 54066
rect 30683 54020 30855 54026
rect 30583 53980 30855 54020
rect 30901 53980 30956 54026
rect 30583 53903 30956 53980
rect 30583 53857 30637 53903
rect 30683 53862 30956 53903
rect 30683 53857 30855 53862
rect 30583 53816 30855 53857
rect 30901 53816 30956 53862
rect 30583 53740 30956 53816
rect 30583 53694 30637 53740
rect 30683 53699 30956 53740
rect 30683 53694 30855 53699
rect 30583 53653 30855 53694
rect 30901 53653 30956 53699
rect 30583 53577 30956 53653
rect 30583 53531 30637 53577
rect 30683 53536 30956 53577
rect 30683 53531 30855 53536
rect 30583 53490 30855 53531
rect 30901 53490 30956 53536
rect 36348 54058 36861 54104
rect 39007 54150 39321 54207
rect 39007 54104 39062 54150
rect 39108 54104 39220 54150
rect 39266 54104 39321 54150
rect 39007 54047 39321 54104
rect 45564 54314 48566 54371
rect 45564 54268 45619 54314
rect 45665 54268 45777 54314
rect 45823 54268 45935 54314
rect 45981 54268 46093 54314
rect 46139 54268 46251 54314
rect 46297 54268 46409 54314
rect 46455 54268 46568 54314
rect 46614 54268 46726 54314
rect 46772 54268 46884 54314
rect 46930 54268 47042 54314
rect 47088 54268 47200 54314
rect 47246 54268 47358 54314
rect 47404 54268 47516 54314
rect 47562 54268 47675 54314
rect 47721 54268 47833 54314
rect 47879 54268 47991 54314
rect 48037 54268 48149 54314
rect 48195 54268 48307 54314
rect 48353 54268 48465 54314
rect 48511 54268 48566 54314
rect 54168 54723 54540 54841
rect 54168 54677 54440 54723
rect 54486 54677 54540 54723
rect 54168 54560 54540 54677
rect 54168 54514 54440 54560
rect 54486 54514 54540 54560
rect 54168 54438 54540 54514
rect 54168 54392 54223 54438
rect 54269 54397 54540 54438
rect 54269 54392 54440 54397
rect 54168 54351 54440 54392
rect 54486 54351 54540 54397
rect 45564 54196 48566 54268
rect 45564 54150 48766 54196
rect 54168 54274 54540 54351
rect 54168 54228 54223 54274
rect 54269 54234 54540 54274
rect 54269 54228 54440 54234
rect 54168 54188 54440 54228
rect 54486 54188 54540 54234
rect 45564 54104 45619 54150
rect 45665 54104 45777 54150
rect 45823 54104 45935 54150
rect 45981 54104 46093 54150
rect 46139 54104 46251 54150
rect 46297 54104 46409 54150
rect 46455 54104 46568 54150
rect 46614 54104 46726 54150
rect 46772 54104 46884 54150
rect 46930 54104 47042 54150
rect 47088 54104 47200 54150
rect 47246 54104 47358 54150
rect 47404 54104 47516 54150
rect 47562 54104 47675 54150
rect 47721 54104 47833 54150
rect 47879 54104 47991 54150
rect 48037 54104 48149 54150
rect 48195 54104 48307 54150
rect 48353 54104 48465 54150
rect 48511 54104 48766 54150
rect 45564 54058 48766 54104
rect 45564 53986 48566 54058
rect 45564 53940 45619 53986
rect 45665 53940 45777 53986
rect 45823 53940 45935 53986
rect 45981 53940 46093 53986
rect 46139 53940 46251 53986
rect 46297 53940 46409 53986
rect 46455 53940 46568 53986
rect 46614 53940 46726 53986
rect 46772 53940 46884 53986
rect 46930 53940 47042 53986
rect 47088 53940 47200 53986
rect 47246 53940 47358 53986
rect 47404 53940 47516 53986
rect 47562 53940 47675 53986
rect 47721 53940 47833 53986
rect 47879 53940 47991 53986
rect 48037 53940 48149 53986
rect 48195 53940 48307 53986
rect 48353 53940 48465 53986
rect 48511 53940 48566 53986
rect 54168 54066 54540 54188
rect 54168 54026 54440 54066
rect 54168 53980 54223 54026
rect 54269 54020 54440 54026
rect 54486 54020 54540 54066
rect 54269 53980 54540 54020
rect 45564 53883 48566 53940
rect 30583 53413 30956 53490
rect 30583 53367 30637 53413
rect 30683 53373 30956 53413
rect 30683 53367 30855 53373
rect 30583 53327 30855 53367
rect 30901 53327 30956 53373
rect 54168 53903 54540 53980
rect 54168 53862 54440 53903
rect 54168 53816 54223 53862
rect 54269 53857 54440 53862
rect 54486 53857 54540 53903
rect 54269 53816 54540 53857
rect 54168 53740 54540 53816
rect 54168 53694 54440 53740
rect 54486 53694 54540 53740
rect 54168 53577 54540 53694
rect 54168 53531 54440 53577
rect 54486 53531 54540 53577
rect 54168 53413 54540 53531
rect 54168 53373 54440 53413
rect 30583 53250 30956 53327
rect 54168 53327 54223 53373
rect 54269 53367 54440 53373
rect 54486 53367 54540 53413
rect 54269 53327 54540 53367
rect 30583 53204 30637 53250
rect 30683 53204 30956 53250
rect 30583 53127 30956 53204
rect 54168 53250 54540 53327
rect 54168 53204 54440 53250
rect 54486 53204 54540 53250
rect 30583 53087 30855 53127
rect 30583 53041 30637 53087
rect 30683 53081 30855 53087
rect 30901 53081 30956 53127
rect 54168 53127 54540 53204
rect 30683 53041 30956 53081
rect 30583 52964 30956 53041
rect 30583 52923 30855 52964
rect 30583 52877 30637 52923
rect 30683 52918 30855 52923
rect 30901 52918 30956 52964
rect 30683 52877 30956 52918
rect 30583 52801 30956 52877
rect 30583 52760 30855 52801
rect 30583 52714 30637 52760
rect 30683 52755 30855 52760
rect 30901 52755 30956 52801
rect 30683 52714 30956 52755
rect 30583 52638 30956 52714
rect 30583 52597 30855 52638
rect 30583 52551 30637 52597
rect 30683 52592 30855 52597
rect 30901 52592 30956 52638
rect 30683 52551 30956 52592
rect 30583 52474 30956 52551
rect 30583 52434 30855 52474
rect 30583 52388 30637 52434
rect 30683 52428 30855 52434
rect 30901 52428 30956 52474
rect 30683 52388 30956 52428
rect 30583 52266 30956 52388
rect 54168 53081 54223 53127
rect 54269 53087 54540 53127
rect 54269 53081 54440 53087
rect 54168 53041 54440 53081
rect 54486 53041 54540 53087
rect 36348 52350 36861 52396
rect 36348 52304 36489 52350
rect 36723 52304 36861 52350
rect 30583 52220 30637 52266
rect 30683 52226 30956 52266
rect 30683 52220 30855 52226
rect 30583 52180 30855 52220
rect 30901 52180 30956 52226
rect 30583 52103 30956 52180
rect 30583 52057 30637 52103
rect 30683 52062 30956 52103
rect 30683 52057 30855 52062
rect 30583 52016 30855 52057
rect 30901 52016 30956 52062
rect 30583 51940 30956 52016
rect 30583 51894 30637 51940
rect 30683 51899 30956 51940
rect 30683 51894 30855 51899
rect 30583 51853 30855 51894
rect 30901 51853 30956 51899
rect 30583 51777 30956 51853
rect 30583 51731 30637 51777
rect 30683 51736 30956 51777
rect 30683 51731 30855 51736
rect 30583 51690 30855 51731
rect 30901 51690 30956 51736
rect 36348 52258 36861 52304
rect 39007 52350 39321 52407
rect 39007 52304 39062 52350
rect 39108 52304 39220 52350
rect 39266 52304 39321 52350
rect 39007 52247 39321 52304
rect 45564 52514 48566 52571
rect 45564 52468 45619 52514
rect 45665 52468 45777 52514
rect 45823 52468 45935 52514
rect 45981 52468 46093 52514
rect 46139 52468 46251 52514
rect 46297 52468 46409 52514
rect 46455 52468 46568 52514
rect 46614 52468 46726 52514
rect 46772 52468 46884 52514
rect 46930 52468 47042 52514
rect 47088 52468 47200 52514
rect 47246 52468 47358 52514
rect 47404 52468 47516 52514
rect 47562 52468 47675 52514
rect 47721 52468 47833 52514
rect 47879 52468 47991 52514
rect 48037 52468 48149 52514
rect 48195 52468 48307 52514
rect 48353 52468 48465 52514
rect 48511 52468 48566 52514
rect 54168 52923 54540 53041
rect 54168 52877 54440 52923
rect 54486 52877 54540 52923
rect 54168 52760 54540 52877
rect 54168 52714 54440 52760
rect 54486 52714 54540 52760
rect 54168 52638 54540 52714
rect 54168 52592 54223 52638
rect 54269 52597 54540 52638
rect 54269 52592 54440 52597
rect 54168 52551 54440 52592
rect 54486 52551 54540 52597
rect 45564 52396 48566 52468
rect 45564 52350 48766 52396
rect 54168 52474 54540 52551
rect 54168 52428 54223 52474
rect 54269 52434 54540 52474
rect 54269 52428 54440 52434
rect 54168 52388 54440 52428
rect 54486 52388 54540 52434
rect 45564 52304 45619 52350
rect 45665 52304 45777 52350
rect 45823 52304 45935 52350
rect 45981 52304 46093 52350
rect 46139 52304 46251 52350
rect 46297 52304 46409 52350
rect 46455 52304 46568 52350
rect 46614 52304 46726 52350
rect 46772 52304 46884 52350
rect 46930 52304 47042 52350
rect 47088 52304 47200 52350
rect 47246 52304 47358 52350
rect 47404 52304 47516 52350
rect 47562 52304 47675 52350
rect 47721 52304 47833 52350
rect 47879 52304 47991 52350
rect 48037 52304 48149 52350
rect 48195 52304 48307 52350
rect 48353 52304 48465 52350
rect 48511 52304 48766 52350
rect 45564 52258 48766 52304
rect 45564 52186 48566 52258
rect 45564 52140 45619 52186
rect 45665 52140 45777 52186
rect 45823 52140 45935 52186
rect 45981 52140 46093 52186
rect 46139 52140 46251 52186
rect 46297 52140 46409 52186
rect 46455 52140 46568 52186
rect 46614 52140 46726 52186
rect 46772 52140 46884 52186
rect 46930 52140 47042 52186
rect 47088 52140 47200 52186
rect 47246 52140 47358 52186
rect 47404 52140 47516 52186
rect 47562 52140 47675 52186
rect 47721 52140 47833 52186
rect 47879 52140 47991 52186
rect 48037 52140 48149 52186
rect 48195 52140 48307 52186
rect 48353 52140 48465 52186
rect 48511 52140 48566 52186
rect 54168 52266 54540 52388
rect 54168 52226 54440 52266
rect 54168 52180 54223 52226
rect 54269 52220 54440 52226
rect 54486 52220 54540 52266
rect 54269 52180 54540 52220
rect 45564 52083 48566 52140
rect 30583 51613 30956 51690
rect 30583 51567 30637 51613
rect 30683 51573 30956 51613
rect 30683 51567 30855 51573
rect 30583 51527 30855 51567
rect 30901 51527 30956 51573
rect 54168 52103 54540 52180
rect 54168 52062 54440 52103
rect 54168 52016 54223 52062
rect 54269 52057 54440 52062
rect 54486 52057 54540 52103
rect 54269 52016 54540 52057
rect 54168 51940 54540 52016
rect 54168 51894 54440 51940
rect 54486 51894 54540 51940
rect 54168 51777 54540 51894
rect 54168 51731 54440 51777
rect 54486 51731 54540 51777
rect 54168 51613 54540 51731
rect 54168 51573 54440 51613
rect 30583 51450 30956 51527
rect 54168 51527 54223 51573
rect 54269 51567 54440 51573
rect 54486 51567 54540 51613
rect 54269 51527 54540 51567
rect 30583 51404 30637 51450
rect 30683 51404 30956 51450
rect 30583 51327 30956 51404
rect 54168 51450 54540 51527
rect 54168 51404 54440 51450
rect 54486 51404 54540 51450
rect 30583 51287 30855 51327
rect 30583 51241 30637 51287
rect 30683 51281 30855 51287
rect 30901 51281 30956 51327
rect 54168 51327 54540 51404
rect 30683 51241 30956 51281
rect 30583 51164 30956 51241
rect 30583 51123 30855 51164
rect 30583 51077 30637 51123
rect 30683 51118 30855 51123
rect 30901 51118 30956 51164
rect 30683 51077 30956 51118
rect 30583 51001 30956 51077
rect 30583 50960 30855 51001
rect 30583 50914 30637 50960
rect 30683 50955 30855 50960
rect 30901 50955 30956 51001
rect 30683 50914 30956 50955
rect 30583 50838 30956 50914
rect 30583 50797 30855 50838
rect 30583 50751 30637 50797
rect 30683 50792 30855 50797
rect 30901 50792 30956 50838
rect 30683 50751 30956 50792
rect 30583 50674 30956 50751
rect 30583 50634 30855 50674
rect 30583 50588 30637 50634
rect 30683 50628 30855 50634
rect 30901 50628 30956 50674
rect 30683 50588 30956 50628
rect 30583 50466 30956 50588
rect 54168 51281 54223 51327
rect 54269 51287 54540 51327
rect 54269 51281 54440 51287
rect 54168 51241 54440 51281
rect 54486 51241 54540 51287
rect 36348 50550 36861 50596
rect 36348 50504 36489 50550
rect 36723 50504 36861 50550
rect 30583 50420 30637 50466
rect 30683 50426 30956 50466
rect 30683 50420 30855 50426
rect 30583 50380 30855 50420
rect 30901 50380 30956 50426
rect 30583 50303 30956 50380
rect 30583 50257 30637 50303
rect 30683 50262 30956 50303
rect 30683 50257 30855 50262
rect 30583 50216 30855 50257
rect 30901 50216 30956 50262
rect 30583 50140 30956 50216
rect 30583 50094 30637 50140
rect 30683 50099 30956 50140
rect 30683 50094 30855 50099
rect 30583 50053 30855 50094
rect 30901 50053 30956 50099
rect 30583 49977 30956 50053
rect 30583 49931 30637 49977
rect 30683 49936 30956 49977
rect 30683 49931 30855 49936
rect 30583 49890 30855 49931
rect 30901 49890 30956 49936
rect 36348 50458 36861 50504
rect 39007 50550 39321 50607
rect 39007 50504 39062 50550
rect 39108 50504 39220 50550
rect 39266 50504 39321 50550
rect 39007 50447 39321 50504
rect 45564 50714 48566 50771
rect 45564 50668 45619 50714
rect 45665 50668 45777 50714
rect 45823 50668 45935 50714
rect 45981 50668 46093 50714
rect 46139 50668 46251 50714
rect 46297 50668 46409 50714
rect 46455 50668 46568 50714
rect 46614 50668 46726 50714
rect 46772 50668 46884 50714
rect 46930 50668 47042 50714
rect 47088 50668 47200 50714
rect 47246 50668 47358 50714
rect 47404 50668 47516 50714
rect 47562 50668 47675 50714
rect 47721 50668 47833 50714
rect 47879 50668 47991 50714
rect 48037 50668 48149 50714
rect 48195 50668 48307 50714
rect 48353 50668 48465 50714
rect 48511 50668 48566 50714
rect 54168 51123 54540 51241
rect 54168 51077 54440 51123
rect 54486 51077 54540 51123
rect 54168 50960 54540 51077
rect 54168 50914 54440 50960
rect 54486 50914 54540 50960
rect 54168 50838 54540 50914
rect 54168 50792 54223 50838
rect 54269 50797 54540 50838
rect 54269 50792 54440 50797
rect 54168 50751 54440 50792
rect 54486 50751 54540 50797
rect 45564 50596 48566 50668
rect 45564 50550 48766 50596
rect 54168 50674 54540 50751
rect 54168 50628 54223 50674
rect 54269 50634 54540 50674
rect 54269 50628 54440 50634
rect 54168 50588 54440 50628
rect 54486 50588 54540 50634
rect 45564 50504 45619 50550
rect 45665 50504 45777 50550
rect 45823 50504 45935 50550
rect 45981 50504 46093 50550
rect 46139 50504 46251 50550
rect 46297 50504 46409 50550
rect 46455 50504 46568 50550
rect 46614 50504 46726 50550
rect 46772 50504 46884 50550
rect 46930 50504 47042 50550
rect 47088 50504 47200 50550
rect 47246 50504 47358 50550
rect 47404 50504 47516 50550
rect 47562 50504 47675 50550
rect 47721 50504 47833 50550
rect 47879 50504 47991 50550
rect 48037 50504 48149 50550
rect 48195 50504 48307 50550
rect 48353 50504 48465 50550
rect 48511 50504 48766 50550
rect 45564 50458 48766 50504
rect 45564 50386 48566 50458
rect 45564 50340 45619 50386
rect 45665 50340 45777 50386
rect 45823 50340 45935 50386
rect 45981 50340 46093 50386
rect 46139 50340 46251 50386
rect 46297 50340 46409 50386
rect 46455 50340 46568 50386
rect 46614 50340 46726 50386
rect 46772 50340 46884 50386
rect 46930 50340 47042 50386
rect 47088 50340 47200 50386
rect 47246 50340 47358 50386
rect 47404 50340 47516 50386
rect 47562 50340 47675 50386
rect 47721 50340 47833 50386
rect 47879 50340 47991 50386
rect 48037 50340 48149 50386
rect 48195 50340 48307 50386
rect 48353 50340 48465 50386
rect 48511 50340 48566 50386
rect 54168 50466 54540 50588
rect 54168 50426 54440 50466
rect 54168 50380 54223 50426
rect 54269 50420 54440 50426
rect 54486 50420 54540 50466
rect 54269 50380 54540 50420
rect 45564 50283 48566 50340
rect 30583 49813 30956 49890
rect 30583 49767 30637 49813
rect 30683 49773 30956 49813
rect 30683 49767 30855 49773
rect 30583 49727 30855 49767
rect 30901 49727 30956 49773
rect 54168 50303 54540 50380
rect 54168 50262 54440 50303
rect 54168 50216 54223 50262
rect 54269 50257 54440 50262
rect 54486 50257 54540 50303
rect 54269 50216 54540 50257
rect 54168 50140 54540 50216
rect 54168 50094 54440 50140
rect 54486 50094 54540 50140
rect 54168 49977 54540 50094
rect 54168 49931 54440 49977
rect 54486 49931 54540 49977
rect 54168 49813 54540 49931
rect 54168 49773 54440 49813
rect 30583 49650 30956 49727
rect 54168 49727 54223 49773
rect 54269 49767 54440 49773
rect 54486 49767 54540 49813
rect 54269 49727 54540 49767
rect 30583 49604 30637 49650
rect 30683 49604 30956 49650
rect 30583 49527 30956 49604
rect 54168 49650 54540 49727
rect 54168 49604 54440 49650
rect 54486 49604 54540 49650
rect 30583 49487 30855 49527
rect 30583 49441 30637 49487
rect 30683 49481 30855 49487
rect 30901 49481 30956 49527
rect 54168 49527 54540 49604
rect 30683 49441 30956 49481
rect 30583 49364 30956 49441
rect 30583 49323 30855 49364
rect 30583 49277 30637 49323
rect 30683 49318 30855 49323
rect 30901 49318 30956 49364
rect 30683 49277 30956 49318
rect 30583 49201 30956 49277
rect 30583 49160 30855 49201
rect 30583 49114 30637 49160
rect 30683 49155 30855 49160
rect 30901 49155 30956 49201
rect 30683 49114 30956 49155
rect 30583 49038 30956 49114
rect 30583 48997 30855 49038
rect 30583 48951 30637 48997
rect 30683 48992 30855 48997
rect 30901 48992 30956 49038
rect 30683 48951 30956 48992
rect 30583 48874 30956 48951
rect 30583 48834 30855 48874
rect 30583 48788 30637 48834
rect 30683 48828 30855 48834
rect 30901 48828 30956 48874
rect 30683 48788 30956 48828
rect 30583 48666 30956 48788
rect 54168 49481 54223 49527
rect 54269 49487 54540 49527
rect 54269 49481 54440 49487
rect 54168 49441 54440 49481
rect 54486 49441 54540 49487
rect 36348 48750 36861 48796
rect 36348 48704 36489 48750
rect 36723 48704 36861 48750
rect 30583 48620 30637 48666
rect 30683 48626 30956 48666
rect 30683 48620 30855 48626
rect 30583 48580 30855 48620
rect 30901 48580 30956 48626
rect 30583 48503 30956 48580
rect 30583 48457 30637 48503
rect 30683 48462 30956 48503
rect 30683 48457 30855 48462
rect 30583 48416 30855 48457
rect 30901 48416 30956 48462
rect 30583 48340 30956 48416
rect 30583 48294 30637 48340
rect 30683 48299 30956 48340
rect 30683 48294 30855 48299
rect 30583 48253 30855 48294
rect 30901 48253 30956 48299
rect 30583 48177 30956 48253
rect 30583 48131 30637 48177
rect 30683 48136 30956 48177
rect 30683 48131 30855 48136
rect 30583 48090 30855 48131
rect 30901 48090 30956 48136
rect 36348 48658 36861 48704
rect 39007 48750 39321 48807
rect 39007 48704 39062 48750
rect 39108 48704 39220 48750
rect 39266 48704 39321 48750
rect 39007 48647 39321 48704
rect 45564 48914 48566 48971
rect 45564 48868 45619 48914
rect 45665 48868 45777 48914
rect 45823 48868 45935 48914
rect 45981 48868 46093 48914
rect 46139 48868 46251 48914
rect 46297 48868 46409 48914
rect 46455 48868 46568 48914
rect 46614 48868 46726 48914
rect 46772 48868 46884 48914
rect 46930 48868 47042 48914
rect 47088 48868 47200 48914
rect 47246 48868 47358 48914
rect 47404 48868 47516 48914
rect 47562 48868 47675 48914
rect 47721 48868 47833 48914
rect 47879 48868 47991 48914
rect 48037 48868 48149 48914
rect 48195 48868 48307 48914
rect 48353 48868 48465 48914
rect 48511 48868 48566 48914
rect 54168 49323 54540 49441
rect 54168 49277 54440 49323
rect 54486 49277 54540 49323
rect 54168 49160 54540 49277
rect 54168 49114 54440 49160
rect 54486 49114 54540 49160
rect 54168 49038 54540 49114
rect 54168 48992 54223 49038
rect 54269 48997 54540 49038
rect 54269 48992 54440 48997
rect 54168 48951 54440 48992
rect 54486 48951 54540 48997
rect 45564 48796 48566 48868
rect 45564 48750 48766 48796
rect 54168 48874 54540 48951
rect 54168 48828 54223 48874
rect 54269 48834 54540 48874
rect 54269 48828 54440 48834
rect 54168 48788 54440 48828
rect 54486 48788 54540 48834
rect 45564 48704 45619 48750
rect 45665 48704 45777 48750
rect 45823 48704 45935 48750
rect 45981 48704 46093 48750
rect 46139 48704 46251 48750
rect 46297 48704 46409 48750
rect 46455 48704 46568 48750
rect 46614 48704 46726 48750
rect 46772 48704 46884 48750
rect 46930 48704 47042 48750
rect 47088 48704 47200 48750
rect 47246 48704 47358 48750
rect 47404 48704 47516 48750
rect 47562 48704 47675 48750
rect 47721 48704 47833 48750
rect 47879 48704 47991 48750
rect 48037 48704 48149 48750
rect 48195 48704 48307 48750
rect 48353 48704 48465 48750
rect 48511 48704 48766 48750
rect 45564 48658 48766 48704
rect 45564 48586 48566 48658
rect 45564 48540 45619 48586
rect 45665 48540 45777 48586
rect 45823 48540 45935 48586
rect 45981 48540 46093 48586
rect 46139 48540 46251 48586
rect 46297 48540 46409 48586
rect 46455 48540 46568 48586
rect 46614 48540 46726 48586
rect 46772 48540 46884 48586
rect 46930 48540 47042 48586
rect 47088 48540 47200 48586
rect 47246 48540 47358 48586
rect 47404 48540 47516 48586
rect 47562 48540 47675 48586
rect 47721 48540 47833 48586
rect 47879 48540 47991 48586
rect 48037 48540 48149 48586
rect 48195 48540 48307 48586
rect 48353 48540 48465 48586
rect 48511 48540 48566 48586
rect 54168 48666 54540 48788
rect 54168 48626 54440 48666
rect 54168 48580 54223 48626
rect 54269 48620 54440 48626
rect 54486 48620 54540 48666
rect 54269 48580 54540 48620
rect 45564 48483 48566 48540
rect 30583 48013 30956 48090
rect 30583 47967 30637 48013
rect 30683 47973 30956 48013
rect 30683 47967 30855 47973
rect 30583 47927 30855 47967
rect 30901 47927 30956 47973
rect 54168 48503 54540 48580
rect 54168 48462 54440 48503
rect 54168 48416 54223 48462
rect 54269 48457 54440 48462
rect 54486 48457 54540 48503
rect 54269 48416 54540 48457
rect 54168 48340 54540 48416
rect 54168 48294 54440 48340
rect 54486 48294 54540 48340
rect 54168 48177 54540 48294
rect 54168 48131 54440 48177
rect 54486 48131 54540 48177
rect 54168 48013 54540 48131
rect 54168 47973 54440 48013
rect 30583 47850 30956 47927
rect 54168 47927 54223 47973
rect 54269 47967 54440 47973
rect 54486 47967 54540 48013
rect 54269 47927 54540 47967
rect 30583 47804 30637 47850
rect 30683 47804 30956 47850
rect 30583 47727 30956 47804
rect 54168 47850 54540 47927
rect 54168 47804 54440 47850
rect 54486 47804 54540 47850
rect 30583 47687 30855 47727
rect 30583 47641 30637 47687
rect 30683 47681 30855 47687
rect 30901 47681 30956 47727
rect 54168 47727 54540 47804
rect 30683 47641 30956 47681
rect 30583 47564 30956 47641
rect 30583 47523 30855 47564
rect 30583 47477 30637 47523
rect 30683 47518 30855 47523
rect 30901 47518 30956 47564
rect 30683 47477 30956 47518
rect 30583 47401 30956 47477
rect 30583 47360 30855 47401
rect 30583 47314 30637 47360
rect 30683 47355 30855 47360
rect 30901 47355 30956 47401
rect 30683 47314 30956 47355
rect 30583 47238 30956 47314
rect 30583 47197 30855 47238
rect 30583 47151 30637 47197
rect 30683 47192 30855 47197
rect 30901 47192 30956 47238
rect 30683 47151 30956 47192
rect 30583 47074 30956 47151
rect 30583 47034 30855 47074
rect 30583 46988 30637 47034
rect 30683 47028 30855 47034
rect 30901 47028 30956 47074
rect 30683 46988 30956 47028
rect 30583 46866 30956 46988
rect 54168 47681 54223 47727
rect 54269 47687 54540 47727
rect 54269 47681 54440 47687
rect 54168 47641 54440 47681
rect 54486 47641 54540 47687
rect 36348 46950 36861 46996
rect 36348 46904 36489 46950
rect 36723 46904 36861 46950
rect 30583 46820 30637 46866
rect 30683 46826 30956 46866
rect 30683 46820 30855 46826
rect 30583 46780 30855 46820
rect 30901 46780 30956 46826
rect 30583 46703 30956 46780
rect 30583 46657 30637 46703
rect 30683 46662 30956 46703
rect 30683 46657 30855 46662
rect 30583 46616 30855 46657
rect 30901 46616 30956 46662
rect 30583 46540 30956 46616
rect 30583 46494 30637 46540
rect 30683 46499 30956 46540
rect 30683 46494 30855 46499
rect 30583 46453 30855 46494
rect 30901 46453 30956 46499
rect 30583 46377 30956 46453
rect 30583 46331 30637 46377
rect 30683 46336 30956 46377
rect 30683 46331 30855 46336
rect 30583 46290 30855 46331
rect 30901 46290 30956 46336
rect 36348 46858 36861 46904
rect 39007 46950 39321 47007
rect 39007 46904 39062 46950
rect 39108 46904 39220 46950
rect 39266 46904 39321 46950
rect 39007 46847 39321 46904
rect 45564 47114 48566 47171
rect 45564 47068 45619 47114
rect 45665 47068 45777 47114
rect 45823 47068 45935 47114
rect 45981 47068 46093 47114
rect 46139 47068 46251 47114
rect 46297 47068 46409 47114
rect 46455 47068 46568 47114
rect 46614 47068 46726 47114
rect 46772 47068 46884 47114
rect 46930 47068 47042 47114
rect 47088 47068 47200 47114
rect 47246 47068 47358 47114
rect 47404 47068 47516 47114
rect 47562 47068 47675 47114
rect 47721 47068 47833 47114
rect 47879 47068 47991 47114
rect 48037 47068 48149 47114
rect 48195 47068 48307 47114
rect 48353 47068 48465 47114
rect 48511 47068 48566 47114
rect 54168 47523 54540 47641
rect 54168 47477 54440 47523
rect 54486 47477 54540 47523
rect 54168 47360 54540 47477
rect 54168 47314 54440 47360
rect 54486 47314 54540 47360
rect 54168 47238 54540 47314
rect 54168 47192 54223 47238
rect 54269 47197 54540 47238
rect 54269 47192 54440 47197
rect 54168 47151 54440 47192
rect 54486 47151 54540 47197
rect 45564 46996 48566 47068
rect 45564 46950 48766 46996
rect 54168 47074 54540 47151
rect 54168 47028 54223 47074
rect 54269 47034 54540 47074
rect 54269 47028 54440 47034
rect 54168 46988 54440 47028
rect 54486 46988 54540 47034
rect 45564 46904 45619 46950
rect 45665 46904 45777 46950
rect 45823 46904 45935 46950
rect 45981 46904 46093 46950
rect 46139 46904 46251 46950
rect 46297 46904 46409 46950
rect 46455 46904 46568 46950
rect 46614 46904 46726 46950
rect 46772 46904 46884 46950
rect 46930 46904 47042 46950
rect 47088 46904 47200 46950
rect 47246 46904 47358 46950
rect 47404 46904 47516 46950
rect 47562 46904 47675 46950
rect 47721 46904 47833 46950
rect 47879 46904 47991 46950
rect 48037 46904 48149 46950
rect 48195 46904 48307 46950
rect 48353 46904 48465 46950
rect 48511 46904 48766 46950
rect 45564 46858 48766 46904
rect 45564 46786 48566 46858
rect 45564 46740 45619 46786
rect 45665 46740 45777 46786
rect 45823 46740 45935 46786
rect 45981 46740 46093 46786
rect 46139 46740 46251 46786
rect 46297 46740 46409 46786
rect 46455 46740 46568 46786
rect 46614 46740 46726 46786
rect 46772 46740 46884 46786
rect 46930 46740 47042 46786
rect 47088 46740 47200 46786
rect 47246 46740 47358 46786
rect 47404 46740 47516 46786
rect 47562 46740 47675 46786
rect 47721 46740 47833 46786
rect 47879 46740 47991 46786
rect 48037 46740 48149 46786
rect 48195 46740 48307 46786
rect 48353 46740 48465 46786
rect 48511 46740 48566 46786
rect 54168 46866 54540 46988
rect 54168 46826 54440 46866
rect 54168 46780 54223 46826
rect 54269 46820 54440 46826
rect 54486 46820 54540 46866
rect 54269 46780 54540 46820
rect 45564 46683 48566 46740
rect 30583 46213 30956 46290
rect 30583 46167 30637 46213
rect 30683 46173 30956 46213
rect 30683 46167 30855 46173
rect 30583 46127 30855 46167
rect 30901 46127 30956 46173
rect 54168 46703 54540 46780
rect 54168 46662 54440 46703
rect 54168 46616 54223 46662
rect 54269 46657 54440 46662
rect 54486 46657 54540 46703
rect 54269 46616 54540 46657
rect 54168 46540 54540 46616
rect 54168 46494 54440 46540
rect 54486 46494 54540 46540
rect 54168 46377 54540 46494
rect 54168 46331 54440 46377
rect 54486 46331 54540 46377
rect 54168 46213 54540 46331
rect 54168 46173 54440 46213
rect 30583 46050 30956 46127
rect 54168 46127 54223 46173
rect 54269 46167 54440 46173
rect 54486 46167 54540 46213
rect 54269 46127 54540 46167
rect 30583 46004 30637 46050
rect 30683 46004 30956 46050
rect 30583 45927 30956 46004
rect 54168 46050 54540 46127
rect 54168 46004 54440 46050
rect 54486 46004 54540 46050
rect 30583 45887 30855 45927
rect 30583 45841 30637 45887
rect 30683 45881 30855 45887
rect 30901 45881 30956 45927
rect 54168 45927 54540 46004
rect 30683 45841 30956 45881
rect 30583 45764 30956 45841
rect 30583 45723 30855 45764
rect 30583 45677 30637 45723
rect 30683 45718 30855 45723
rect 30901 45718 30956 45764
rect 30683 45677 30956 45718
rect 30583 45601 30956 45677
rect 30583 45560 30855 45601
rect 30583 45514 30637 45560
rect 30683 45555 30855 45560
rect 30901 45555 30956 45601
rect 30683 45514 30956 45555
rect 30583 45438 30956 45514
rect 30583 45397 30855 45438
rect 30583 45351 30637 45397
rect 30683 45392 30855 45397
rect 30901 45392 30956 45438
rect 30683 45351 30956 45392
rect 30583 45274 30956 45351
rect 30583 45234 30855 45274
rect 30583 45188 30637 45234
rect 30683 45228 30855 45234
rect 30901 45228 30956 45274
rect 30683 45188 30956 45228
rect 30583 45066 30956 45188
rect 54168 45881 54223 45927
rect 54269 45887 54540 45927
rect 54269 45881 54440 45887
rect 54168 45841 54440 45881
rect 54486 45841 54540 45887
rect 36348 45150 36861 45196
rect 36348 45104 36489 45150
rect 36723 45104 36861 45150
rect 30583 45020 30637 45066
rect 30683 45026 30956 45066
rect 30683 45020 30855 45026
rect 30583 44980 30855 45020
rect 30901 44980 30956 45026
rect 30583 44903 30956 44980
rect 30583 44857 30637 44903
rect 30683 44862 30956 44903
rect 30683 44857 30855 44862
rect 30583 44816 30855 44857
rect 30901 44816 30956 44862
rect 30583 44740 30956 44816
rect 30583 44694 30637 44740
rect 30683 44699 30956 44740
rect 30683 44694 30855 44699
rect 30583 44653 30855 44694
rect 30901 44653 30956 44699
rect 30583 44577 30956 44653
rect 30583 44531 30637 44577
rect 30683 44536 30956 44577
rect 30683 44531 30855 44536
rect 30583 44490 30855 44531
rect 30901 44490 30956 44536
rect 36348 45058 36861 45104
rect 39007 45150 39321 45207
rect 39007 45104 39062 45150
rect 39108 45104 39220 45150
rect 39266 45104 39321 45150
rect 39007 45047 39321 45104
rect 45564 45314 48566 45371
rect 45564 45268 45619 45314
rect 45665 45268 45777 45314
rect 45823 45268 45935 45314
rect 45981 45268 46093 45314
rect 46139 45268 46251 45314
rect 46297 45268 46409 45314
rect 46455 45268 46568 45314
rect 46614 45268 46726 45314
rect 46772 45268 46884 45314
rect 46930 45268 47042 45314
rect 47088 45268 47200 45314
rect 47246 45268 47358 45314
rect 47404 45268 47516 45314
rect 47562 45268 47675 45314
rect 47721 45268 47833 45314
rect 47879 45268 47991 45314
rect 48037 45268 48149 45314
rect 48195 45268 48307 45314
rect 48353 45268 48465 45314
rect 48511 45268 48566 45314
rect 54168 45723 54540 45841
rect 54168 45677 54440 45723
rect 54486 45677 54540 45723
rect 54168 45560 54540 45677
rect 54168 45514 54440 45560
rect 54486 45514 54540 45560
rect 54168 45438 54540 45514
rect 54168 45392 54223 45438
rect 54269 45397 54540 45438
rect 54269 45392 54440 45397
rect 54168 45351 54440 45392
rect 54486 45351 54540 45397
rect 45564 45196 48566 45268
rect 45564 45150 48766 45196
rect 54168 45274 54540 45351
rect 54168 45228 54223 45274
rect 54269 45234 54540 45274
rect 54269 45228 54440 45234
rect 54168 45188 54440 45228
rect 54486 45188 54540 45234
rect 45564 45104 45619 45150
rect 45665 45104 45777 45150
rect 45823 45104 45935 45150
rect 45981 45104 46093 45150
rect 46139 45104 46251 45150
rect 46297 45104 46409 45150
rect 46455 45104 46568 45150
rect 46614 45104 46726 45150
rect 46772 45104 46884 45150
rect 46930 45104 47042 45150
rect 47088 45104 47200 45150
rect 47246 45104 47358 45150
rect 47404 45104 47516 45150
rect 47562 45104 47675 45150
rect 47721 45104 47833 45150
rect 47879 45104 47991 45150
rect 48037 45104 48149 45150
rect 48195 45104 48307 45150
rect 48353 45104 48465 45150
rect 48511 45104 48766 45150
rect 45564 45058 48766 45104
rect 45564 44986 48566 45058
rect 45564 44940 45619 44986
rect 45665 44940 45777 44986
rect 45823 44940 45935 44986
rect 45981 44940 46093 44986
rect 46139 44940 46251 44986
rect 46297 44940 46409 44986
rect 46455 44940 46568 44986
rect 46614 44940 46726 44986
rect 46772 44940 46884 44986
rect 46930 44940 47042 44986
rect 47088 44940 47200 44986
rect 47246 44940 47358 44986
rect 47404 44940 47516 44986
rect 47562 44940 47675 44986
rect 47721 44940 47833 44986
rect 47879 44940 47991 44986
rect 48037 44940 48149 44986
rect 48195 44940 48307 44986
rect 48353 44940 48465 44986
rect 48511 44940 48566 44986
rect 54168 45066 54540 45188
rect 54168 45026 54440 45066
rect 54168 44980 54223 45026
rect 54269 45020 54440 45026
rect 54486 45020 54540 45066
rect 54269 44980 54540 45020
rect 45564 44883 48566 44940
rect 30583 44413 30956 44490
rect 30583 44367 30637 44413
rect 30683 44373 30956 44413
rect 30683 44367 30855 44373
rect 30583 44327 30855 44367
rect 30901 44327 30956 44373
rect 54168 44903 54540 44980
rect 54168 44862 54440 44903
rect 54168 44816 54223 44862
rect 54269 44857 54440 44862
rect 54486 44857 54540 44903
rect 54269 44816 54540 44857
rect 54168 44740 54540 44816
rect 54168 44694 54440 44740
rect 54486 44694 54540 44740
rect 54168 44577 54540 44694
rect 54168 44531 54440 44577
rect 54486 44531 54540 44577
rect 54168 44413 54540 44531
rect 54168 44373 54440 44413
rect 30583 44250 30956 44327
rect 54168 44327 54223 44373
rect 54269 44367 54440 44373
rect 54486 44367 54540 44413
rect 54269 44327 54540 44367
rect 30583 44204 30637 44250
rect 30683 44204 30956 44250
rect 30583 44127 30956 44204
rect 54168 44250 54540 44327
rect 54168 44204 54440 44250
rect 54486 44204 54540 44250
rect 30583 44087 30855 44127
rect 30583 44041 30637 44087
rect 30683 44081 30855 44087
rect 30901 44081 30956 44127
rect 54168 44127 54540 44204
rect 30683 44041 30956 44081
rect 30583 43964 30956 44041
rect 30583 43923 30855 43964
rect 30583 43877 30637 43923
rect 30683 43918 30855 43923
rect 30901 43918 30956 43964
rect 30683 43877 30956 43918
rect 30583 43801 30956 43877
rect 30583 43760 30855 43801
rect 30583 43714 30637 43760
rect 30683 43755 30855 43760
rect 30901 43755 30956 43801
rect 30683 43714 30956 43755
rect 30583 43638 30956 43714
rect 30583 43597 30855 43638
rect 30583 43551 30637 43597
rect 30683 43592 30855 43597
rect 30901 43592 30956 43638
rect 30683 43551 30956 43592
rect 30583 43474 30956 43551
rect 30583 43434 30855 43474
rect 30583 43388 30637 43434
rect 30683 43428 30855 43434
rect 30901 43428 30956 43474
rect 30683 43388 30956 43428
rect 30583 43266 30956 43388
rect 54168 44081 54223 44127
rect 54269 44087 54540 44127
rect 54269 44081 54440 44087
rect 54168 44041 54440 44081
rect 54486 44041 54540 44087
rect 36348 43350 36861 43396
rect 36348 43304 36489 43350
rect 36723 43304 36861 43350
rect 30583 43220 30637 43266
rect 30683 43226 30956 43266
rect 30683 43220 30855 43226
rect 30583 43180 30855 43220
rect 30901 43180 30956 43226
rect 30583 43103 30956 43180
rect 30583 43057 30637 43103
rect 30683 43062 30956 43103
rect 30683 43057 30855 43062
rect 30583 43016 30855 43057
rect 30901 43016 30956 43062
rect 30583 42940 30956 43016
rect 30583 42894 30637 42940
rect 30683 42899 30956 42940
rect 30683 42894 30855 42899
rect 30583 42853 30855 42894
rect 30901 42853 30956 42899
rect 30583 42777 30956 42853
rect 30583 42731 30637 42777
rect 30683 42736 30956 42777
rect 30683 42731 30855 42736
rect 30583 42690 30855 42731
rect 30901 42690 30956 42736
rect 36348 43258 36861 43304
rect 39007 43350 39321 43407
rect 39007 43304 39062 43350
rect 39108 43304 39220 43350
rect 39266 43304 39321 43350
rect 39007 43247 39321 43304
rect 45564 43514 48566 43571
rect 45564 43468 45619 43514
rect 45665 43468 45777 43514
rect 45823 43468 45935 43514
rect 45981 43468 46093 43514
rect 46139 43468 46251 43514
rect 46297 43468 46409 43514
rect 46455 43468 46568 43514
rect 46614 43468 46726 43514
rect 46772 43468 46884 43514
rect 46930 43468 47042 43514
rect 47088 43468 47200 43514
rect 47246 43468 47358 43514
rect 47404 43468 47516 43514
rect 47562 43468 47675 43514
rect 47721 43468 47833 43514
rect 47879 43468 47991 43514
rect 48037 43468 48149 43514
rect 48195 43468 48307 43514
rect 48353 43468 48465 43514
rect 48511 43468 48566 43514
rect 54168 43923 54540 44041
rect 54168 43877 54440 43923
rect 54486 43877 54540 43923
rect 54168 43760 54540 43877
rect 54168 43714 54440 43760
rect 54486 43714 54540 43760
rect 54168 43638 54540 43714
rect 54168 43592 54223 43638
rect 54269 43597 54540 43638
rect 54269 43592 54440 43597
rect 54168 43551 54440 43592
rect 54486 43551 54540 43597
rect 45564 43396 48566 43468
rect 45564 43350 48766 43396
rect 54168 43474 54540 43551
rect 54168 43428 54223 43474
rect 54269 43434 54540 43474
rect 54269 43428 54440 43434
rect 54168 43388 54440 43428
rect 54486 43388 54540 43434
rect 45564 43304 45619 43350
rect 45665 43304 45777 43350
rect 45823 43304 45935 43350
rect 45981 43304 46093 43350
rect 46139 43304 46251 43350
rect 46297 43304 46409 43350
rect 46455 43304 46568 43350
rect 46614 43304 46726 43350
rect 46772 43304 46884 43350
rect 46930 43304 47042 43350
rect 47088 43304 47200 43350
rect 47246 43304 47358 43350
rect 47404 43304 47516 43350
rect 47562 43304 47675 43350
rect 47721 43304 47833 43350
rect 47879 43304 47991 43350
rect 48037 43304 48149 43350
rect 48195 43304 48307 43350
rect 48353 43304 48465 43350
rect 48511 43304 48766 43350
rect 45564 43258 48766 43304
rect 45564 43186 48566 43258
rect 45564 43140 45619 43186
rect 45665 43140 45777 43186
rect 45823 43140 45935 43186
rect 45981 43140 46093 43186
rect 46139 43140 46251 43186
rect 46297 43140 46409 43186
rect 46455 43140 46568 43186
rect 46614 43140 46726 43186
rect 46772 43140 46884 43186
rect 46930 43140 47042 43186
rect 47088 43140 47200 43186
rect 47246 43140 47358 43186
rect 47404 43140 47516 43186
rect 47562 43140 47675 43186
rect 47721 43140 47833 43186
rect 47879 43140 47991 43186
rect 48037 43140 48149 43186
rect 48195 43140 48307 43186
rect 48353 43140 48465 43186
rect 48511 43140 48566 43186
rect 54168 43266 54540 43388
rect 54168 43226 54440 43266
rect 54168 43180 54223 43226
rect 54269 43220 54440 43226
rect 54486 43220 54540 43266
rect 54269 43180 54540 43220
rect 45564 43083 48566 43140
rect 30583 42613 30956 42690
rect 30583 42567 30637 42613
rect 30683 42573 30956 42613
rect 30683 42567 30855 42573
rect 30583 42527 30855 42567
rect 30901 42527 30956 42573
rect 54168 43103 54540 43180
rect 54168 43062 54440 43103
rect 54168 43016 54223 43062
rect 54269 43057 54440 43062
rect 54486 43057 54540 43103
rect 54269 43016 54540 43057
rect 54168 42940 54540 43016
rect 54168 42894 54440 42940
rect 54486 42894 54540 42940
rect 54168 42777 54540 42894
rect 54168 42731 54440 42777
rect 54486 42731 54540 42777
rect 54168 42613 54540 42731
rect 54168 42573 54440 42613
rect 30583 42450 30956 42527
rect 54168 42527 54223 42573
rect 54269 42567 54440 42573
rect 54486 42567 54540 42613
rect 54269 42527 54540 42567
rect 30583 42404 30637 42450
rect 30683 42404 30956 42450
rect 30583 42327 30956 42404
rect 54168 42450 54540 42527
rect 54168 42404 54440 42450
rect 54486 42404 54540 42450
rect 30583 42287 30855 42327
rect 30583 42241 30637 42287
rect 30683 42281 30855 42287
rect 30901 42281 30956 42327
rect 54168 42327 54540 42404
rect 30683 42241 30956 42281
rect 30583 42164 30956 42241
rect 30583 42123 30855 42164
rect 30583 42077 30637 42123
rect 30683 42118 30855 42123
rect 30901 42118 30956 42164
rect 30683 42077 30956 42118
rect 30583 42001 30956 42077
rect 30583 41960 30855 42001
rect 30583 41914 30637 41960
rect 30683 41955 30855 41960
rect 30901 41955 30956 42001
rect 30683 41914 30956 41955
rect 30583 41838 30956 41914
rect 30583 41797 30855 41838
rect 30583 41751 30637 41797
rect 30683 41792 30855 41797
rect 30901 41792 30956 41838
rect 30683 41751 30956 41792
rect 30583 41674 30956 41751
rect 30583 41634 30855 41674
rect 30583 41588 30637 41634
rect 30683 41628 30855 41634
rect 30901 41628 30956 41674
rect 30683 41588 30956 41628
rect 30583 41466 30956 41588
rect 54168 42281 54223 42327
rect 54269 42287 54540 42327
rect 54269 42281 54440 42287
rect 54168 42241 54440 42281
rect 54486 42241 54540 42287
rect 36348 41550 36861 41596
rect 36348 41504 36489 41550
rect 36723 41504 36861 41550
rect 30583 41420 30637 41466
rect 30683 41426 30956 41466
rect 30683 41420 30855 41426
rect 30583 41380 30855 41420
rect 30901 41380 30956 41426
rect 30583 41303 30956 41380
rect 30583 41257 30637 41303
rect 30683 41262 30956 41303
rect 30683 41257 30855 41262
rect 30583 41216 30855 41257
rect 30901 41216 30956 41262
rect 30583 41140 30956 41216
rect 30583 41094 30637 41140
rect 30683 41099 30956 41140
rect 30683 41094 30855 41099
rect 30583 41053 30855 41094
rect 30901 41053 30956 41099
rect 30583 40977 30956 41053
rect 30583 40931 30637 40977
rect 30683 40936 30956 40977
rect 30683 40931 30855 40936
rect 30583 40890 30855 40931
rect 30901 40890 30956 40936
rect 36348 41458 36861 41504
rect 39007 41550 39321 41607
rect 39007 41504 39062 41550
rect 39108 41504 39220 41550
rect 39266 41504 39321 41550
rect 39007 41447 39321 41504
rect 45564 41714 48566 41771
rect 45564 41668 45619 41714
rect 45665 41668 45777 41714
rect 45823 41668 45935 41714
rect 45981 41668 46093 41714
rect 46139 41668 46251 41714
rect 46297 41668 46409 41714
rect 46455 41668 46568 41714
rect 46614 41668 46726 41714
rect 46772 41668 46884 41714
rect 46930 41668 47042 41714
rect 47088 41668 47200 41714
rect 47246 41668 47358 41714
rect 47404 41668 47516 41714
rect 47562 41668 47675 41714
rect 47721 41668 47833 41714
rect 47879 41668 47991 41714
rect 48037 41668 48149 41714
rect 48195 41668 48307 41714
rect 48353 41668 48465 41714
rect 48511 41668 48566 41714
rect 54168 42123 54540 42241
rect 54168 42077 54440 42123
rect 54486 42077 54540 42123
rect 54168 41960 54540 42077
rect 54168 41914 54440 41960
rect 54486 41914 54540 41960
rect 54168 41838 54540 41914
rect 54168 41792 54223 41838
rect 54269 41797 54540 41838
rect 54269 41792 54440 41797
rect 54168 41751 54440 41792
rect 54486 41751 54540 41797
rect 45564 41596 48566 41668
rect 45564 41550 48766 41596
rect 54168 41674 54540 41751
rect 54168 41628 54223 41674
rect 54269 41634 54540 41674
rect 54269 41628 54440 41634
rect 54168 41588 54440 41628
rect 54486 41588 54540 41634
rect 45564 41504 45619 41550
rect 45665 41504 45777 41550
rect 45823 41504 45935 41550
rect 45981 41504 46093 41550
rect 46139 41504 46251 41550
rect 46297 41504 46409 41550
rect 46455 41504 46568 41550
rect 46614 41504 46726 41550
rect 46772 41504 46884 41550
rect 46930 41504 47042 41550
rect 47088 41504 47200 41550
rect 47246 41504 47358 41550
rect 47404 41504 47516 41550
rect 47562 41504 47675 41550
rect 47721 41504 47833 41550
rect 47879 41504 47991 41550
rect 48037 41504 48149 41550
rect 48195 41504 48307 41550
rect 48353 41504 48465 41550
rect 48511 41504 48766 41550
rect 45564 41458 48766 41504
rect 45564 41386 48566 41458
rect 45564 41340 45619 41386
rect 45665 41340 45777 41386
rect 45823 41340 45935 41386
rect 45981 41340 46093 41386
rect 46139 41340 46251 41386
rect 46297 41340 46409 41386
rect 46455 41340 46568 41386
rect 46614 41340 46726 41386
rect 46772 41340 46884 41386
rect 46930 41340 47042 41386
rect 47088 41340 47200 41386
rect 47246 41340 47358 41386
rect 47404 41340 47516 41386
rect 47562 41340 47675 41386
rect 47721 41340 47833 41386
rect 47879 41340 47991 41386
rect 48037 41340 48149 41386
rect 48195 41340 48307 41386
rect 48353 41340 48465 41386
rect 48511 41340 48566 41386
rect 54168 41466 54540 41588
rect 54168 41426 54440 41466
rect 54168 41380 54223 41426
rect 54269 41420 54440 41426
rect 54486 41420 54540 41466
rect 54269 41380 54540 41420
rect 45564 41283 48566 41340
rect 30583 40813 30956 40890
rect 30583 40767 30637 40813
rect 30683 40773 30956 40813
rect 30683 40767 30855 40773
rect 30583 40727 30855 40767
rect 30901 40727 30956 40773
rect 54168 41303 54540 41380
rect 54168 41262 54440 41303
rect 54168 41216 54223 41262
rect 54269 41257 54440 41262
rect 54486 41257 54540 41303
rect 54269 41216 54540 41257
rect 54168 41140 54540 41216
rect 54168 41094 54440 41140
rect 54486 41094 54540 41140
rect 54168 40977 54540 41094
rect 54168 40931 54440 40977
rect 54486 40931 54540 40977
rect 54168 40813 54540 40931
rect 54168 40773 54440 40813
rect 30583 40650 30956 40727
rect 54168 40727 54223 40773
rect 54269 40767 54440 40773
rect 54486 40767 54540 40813
rect 54269 40727 54540 40767
rect 30583 40604 30637 40650
rect 30683 40604 30956 40650
rect 30583 40527 30956 40604
rect 54168 40650 54540 40727
rect 54168 40604 54440 40650
rect 54486 40604 54540 40650
rect 30583 40487 30855 40527
rect 30583 40441 30637 40487
rect 30683 40481 30855 40487
rect 30901 40481 30956 40527
rect 54168 40527 54540 40604
rect 30683 40441 30956 40481
rect 30583 40364 30956 40441
rect 30583 40323 30855 40364
rect 30583 40277 30637 40323
rect 30683 40318 30855 40323
rect 30901 40318 30956 40364
rect 30683 40277 30956 40318
rect 30583 40201 30956 40277
rect 30583 40160 30855 40201
rect 30583 40114 30637 40160
rect 30683 40155 30855 40160
rect 30901 40155 30956 40201
rect 30683 40114 30956 40155
rect 30583 40038 30956 40114
rect 30583 39997 30855 40038
rect 30583 39951 30637 39997
rect 30683 39992 30855 39997
rect 30901 39992 30956 40038
rect 30683 39951 30956 39992
rect 30583 39874 30956 39951
rect 30583 39834 30855 39874
rect 30583 39788 30637 39834
rect 30683 39828 30855 39834
rect 30901 39828 30956 39874
rect 30683 39788 30956 39828
rect 30583 39666 30956 39788
rect 54168 40481 54223 40527
rect 54269 40487 54540 40527
rect 54269 40481 54440 40487
rect 54168 40441 54440 40481
rect 54486 40441 54540 40487
rect 36348 39750 36861 39796
rect 36348 39704 36489 39750
rect 36723 39704 36861 39750
rect 30583 39620 30637 39666
rect 30683 39626 30956 39666
rect 30683 39620 30855 39626
rect 30583 39580 30855 39620
rect 30901 39580 30956 39626
rect 30583 39503 30956 39580
rect 30583 39457 30637 39503
rect 30683 39462 30956 39503
rect 30683 39457 30855 39462
rect 30583 39416 30855 39457
rect 30901 39416 30956 39462
rect 30583 39340 30956 39416
rect 30583 39294 30637 39340
rect 30683 39299 30956 39340
rect 30683 39294 30855 39299
rect 30583 39253 30855 39294
rect 30901 39253 30956 39299
rect 30583 39177 30956 39253
rect 30583 39131 30637 39177
rect 30683 39136 30956 39177
rect 30683 39131 30855 39136
rect 30583 39090 30855 39131
rect 30901 39090 30956 39136
rect 36348 39658 36861 39704
rect 39007 39750 39321 39807
rect 39007 39704 39062 39750
rect 39108 39704 39220 39750
rect 39266 39704 39321 39750
rect 39007 39647 39321 39704
rect 45564 39914 48566 39971
rect 45564 39868 45619 39914
rect 45665 39868 45777 39914
rect 45823 39868 45935 39914
rect 45981 39868 46093 39914
rect 46139 39868 46251 39914
rect 46297 39868 46409 39914
rect 46455 39868 46568 39914
rect 46614 39868 46726 39914
rect 46772 39868 46884 39914
rect 46930 39868 47042 39914
rect 47088 39868 47200 39914
rect 47246 39868 47358 39914
rect 47404 39868 47516 39914
rect 47562 39868 47675 39914
rect 47721 39868 47833 39914
rect 47879 39868 47991 39914
rect 48037 39868 48149 39914
rect 48195 39868 48307 39914
rect 48353 39868 48465 39914
rect 48511 39868 48566 39914
rect 54168 40323 54540 40441
rect 54168 40277 54440 40323
rect 54486 40277 54540 40323
rect 54168 40160 54540 40277
rect 54168 40114 54440 40160
rect 54486 40114 54540 40160
rect 54168 40038 54540 40114
rect 54168 39992 54223 40038
rect 54269 39997 54540 40038
rect 54269 39992 54440 39997
rect 54168 39951 54440 39992
rect 54486 39951 54540 39997
rect 45564 39796 48566 39868
rect 45564 39750 48766 39796
rect 54168 39874 54540 39951
rect 54168 39828 54223 39874
rect 54269 39834 54540 39874
rect 54269 39828 54440 39834
rect 54168 39788 54440 39828
rect 54486 39788 54540 39834
rect 45564 39704 45619 39750
rect 45665 39704 45777 39750
rect 45823 39704 45935 39750
rect 45981 39704 46093 39750
rect 46139 39704 46251 39750
rect 46297 39704 46409 39750
rect 46455 39704 46568 39750
rect 46614 39704 46726 39750
rect 46772 39704 46884 39750
rect 46930 39704 47042 39750
rect 47088 39704 47200 39750
rect 47246 39704 47358 39750
rect 47404 39704 47516 39750
rect 47562 39704 47675 39750
rect 47721 39704 47833 39750
rect 47879 39704 47991 39750
rect 48037 39704 48149 39750
rect 48195 39704 48307 39750
rect 48353 39704 48465 39750
rect 48511 39704 48766 39750
rect 45564 39658 48766 39704
rect 45564 39586 48566 39658
rect 45564 39540 45619 39586
rect 45665 39540 45777 39586
rect 45823 39540 45935 39586
rect 45981 39540 46093 39586
rect 46139 39540 46251 39586
rect 46297 39540 46409 39586
rect 46455 39540 46568 39586
rect 46614 39540 46726 39586
rect 46772 39540 46884 39586
rect 46930 39540 47042 39586
rect 47088 39540 47200 39586
rect 47246 39540 47358 39586
rect 47404 39540 47516 39586
rect 47562 39540 47675 39586
rect 47721 39540 47833 39586
rect 47879 39540 47991 39586
rect 48037 39540 48149 39586
rect 48195 39540 48307 39586
rect 48353 39540 48465 39586
rect 48511 39540 48566 39586
rect 54168 39666 54540 39788
rect 54168 39626 54440 39666
rect 54168 39580 54223 39626
rect 54269 39620 54440 39626
rect 54486 39620 54540 39666
rect 54269 39580 54540 39620
rect 45564 39483 48566 39540
rect 30583 39013 30956 39090
rect 30583 38967 30637 39013
rect 30683 38973 30956 39013
rect 30683 38967 30855 38973
rect 30583 38927 30855 38967
rect 30901 38927 30956 38973
rect 54168 39503 54540 39580
rect 54168 39462 54440 39503
rect 54168 39416 54223 39462
rect 54269 39457 54440 39462
rect 54486 39457 54540 39503
rect 54269 39416 54540 39457
rect 54168 39340 54540 39416
rect 54168 39294 54440 39340
rect 54486 39294 54540 39340
rect 54168 39177 54540 39294
rect 54168 39131 54440 39177
rect 54486 39131 54540 39177
rect 54168 39013 54540 39131
rect 54168 38973 54440 39013
rect 30583 38850 30956 38927
rect 54168 38927 54223 38973
rect 54269 38967 54440 38973
rect 54486 38967 54540 39013
rect 54269 38927 54540 38967
rect 30583 38804 30637 38850
rect 30683 38804 30956 38850
rect 30583 38727 30956 38804
rect 54168 38850 54540 38927
rect 54168 38804 54440 38850
rect 54486 38804 54540 38850
rect 30583 38687 30855 38727
rect 30583 38641 30637 38687
rect 30683 38681 30855 38687
rect 30901 38681 30956 38727
rect 54168 38727 54540 38804
rect 30683 38641 30956 38681
rect 30583 38564 30956 38641
rect 30583 38523 30855 38564
rect 30583 38477 30637 38523
rect 30683 38518 30855 38523
rect 30901 38518 30956 38564
rect 30683 38477 30956 38518
rect 30583 38401 30956 38477
rect 30583 38360 30855 38401
rect 30583 38314 30637 38360
rect 30683 38355 30855 38360
rect 30901 38355 30956 38401
rect 30683 38314 30956 38355
rect 30583 38238 30956 38314
rect 30583 38197 30855 38238
rect 30583 38151 30637 38197
rect 30683 38192 30855 38197
rect 30901 38192 30956 38238
rect 30683 38151 30956 38192
rect 30583 38074 30956 38151
rect 30583 38034 30855 38074
rect 30583 37988 30637 38034
rect 30683 38028 30855 38034
rect 30901 38028 30956 38074
rect 30683 37988 30956 38028
rect 30583 37866 30956 37988
rect 54168 38681 54223 38727
rect 54269 38687 54540 38727
rect 54269 38681 54440 38687
rect 54168 38641 54440 38681
rect 54486 38641 54540 38687
rect 36348 37950 36861 37996
rect 36348 37904 36489 37950
rect 36723 37904 36861 37950
rect 30583 37820 30637 37866
rect 30683 37826 30956 37866
rect 30683 37820 30855 37826
rect 30583 37780 30855 37820
rect 30901 37780 30956 37826
rect 30583 37703 30956 37780
rect 30583 37657 30637 37703
rect 30683 37662 30956 37703
rect 30683 37657 30855 37662
rect 30583 37616 30855 37657
rect 30901 37616 30956 37662
rect 30583 37540 30956 37616
rect 30583 37494 30637 37540
rect 30683 37499 30956 37540
rect 30683 37494 30855 37499
rect 30583 37453 30855 37494
rect 30901 37453 30956 37499
rect 30583 37377 30956 37453
rect 30583 37331 30637 37377
rect 30683 37336 30956 37377
rect 30683 37331 30855 37336
rect 30583 37290 30855 37331
rect 30901 37290 30956 37336
rect 36348 37858 36861 37904
rect 39007 37950 39321 38007
rect 39007 37904 39062 37950
rect 39108 37904 39220 37950
rect 39266 37904 39321 37950
rect 39007 37847 39321 37904
rect 45564 38114 48566 38171
rect 45564 38068 45619 38114
rect 45665 38068 45777 38114
rect 45823 38068 45935 38114
rect 45981 38068 46093 38114
rect 46139 38068 46251 38114
rect 46297 38068 46409 38114
rect 46455 38068 46568 38114
rect 46614 38068 46726 38114
rect 46772 38068 46884 38114
rect 46930 38068 47042 38114
rect 47088 38068 47200 38114
rect 47246 38068 47358 38114
rect 47404 38068 47516 38114
rect 47562 38068 47675 38114
rect 47721 38068 47833 38114
rect 47879 38068 47991 38114
rect 48037 38068 48149 38114
rect 48195 38068 48307 38114
rect 48353 38068 48465 38114
rect 48511 38068 48566 38114
rect 54168 38523 54540 38641
rect 54168 38477 54440 38523
rect 54486 38477 54540 38523
rect 54168 38360 54540 38477
rect 54168 38314 54440 38360
rect 54486 38314 54540 38360
rect 54168 38238 54540 38314
rect 54168 38192 54223 38238
rect 54269 38197 54540 38238
rect 54269 38192 54440 38197
rect 54168 38151 54440 38192
rect 54486 38151 54540 38197
rect 45564 37996 48566 38068
rect 45564 37950 48766 37996
rect 54168 38074 54540 38151
rect 54168 38028 54223 38074
rect 54269 38034 54540 38074
rect 54269 38028 54440 38034
rect 54168 37988 54440 38028
rect 54486 37988 54540 38034
rect 45564 37904 45619 37950
rect 45665 37904 45777 37950
rect 45823 37904 45935 37950
rect 45981 37904 46093 37950
rect 46139 37904 46251 37950
rect 46297 37904 46409 37950
rect 46455 37904 46568 37950
rect 46614 37904 46726 37950
rect 46772 37904 46884 37950
rect 46930 37904 47042 37950
rect 47088 37904 47200 37950
rect 47246 37904 47358 37950
rect 47404 37904 47516 37950
rect 47562 37904 47675 37950
rect 47721 37904 47833 37950
rect 47879 37904 47991 37950
rect 48037 37904 48149 37950
rect 48195 37904 48307 37950
rect 48353 37904 48465 37950
rect 48511 37904 48766 37950
rect 45564 37858 48766 37904
rect 45564 37786 48566 37858
rect 45564 37740 45619 37786
rect 45665 37740 45777 37786
rect 45823 37740 45935 37786
rect 45981 37740 46093 37786
rect 46139 37740 46251 37786
rect 46297 37740 46409 37786
rect 46455 37740 46568 37786
rect 46614 37740 46726 37786
rect 46772 37740 46884 37786
rect 46930 37740 47042 37786
rect 47088 37740 47200 37786
rect 47246 37740 47358 37786
rect 47404 37740 47516 37786
rect 47562 37740 47675 37786
rect 47721 37740 47833 37786
rect 47879 37740 47991 37786
rect 48037 37740 48149 37786
rect 48195 37740 48307 37786
rect 48353 37740 48465 37786
rect 48511 37740 48566 37786
rect 54168 37866 54540 37988
rect 54168 37826 54440 37866
rect 54168 37780 54223 37826
rect 54269 37820 54440 37826
rect 54486 37820 54540 37866
rect 54269 37780 54540 37820
rect 45564 37683 48566 37740
rect 30583 37213 30956 37290
rect 30583 37167 30637 37213
rect 30683 37173 30956 37213
rect 30683 37167 30855 37173
rect 30583 37127 30855 37167
rect 30901 37127 30956 37173
rect 54168 37703 54540 37780
rect 54168 37662 54440 37703
rect 54168 37616 54223 37662
rect 54269 37657 54440 37662
rect 54486 37657 54540 37703
rect 54269 37616 54540 37657
rect 54168 37540 54540 37616
rect 54168 37494 54440 37540
rect 54486 37494 54540 37540
rect 54168 37377 54540 37494
rect 54168 37331 54440 37377
rect 54486 37331 54540 37377
rect 54168 37213 54540 37331
rect 54168 37173 54440 37213
rect 30583 37050 30956 37127
rect 54168 37127 54223 37173
rect 54269 37167 54440 37173
rect 54486 37167 54540 37213
rect 54269 37127 54540 37167
rect 30583 37004 30637 37050
rect 30683 37004 30956 37050
rect 30583 36927 30956 37004
rect 54168 37050 54540 37127
rect 54168 37004 54440 37050
rect 54486 37004 54540 37050
rect 30583 36887 30855 36927
rect 30583 36841 30637 36887
rect 30683 36881 30855 36887
rect 30901 36881 30956 36927
rect 54168 36927 54540 37004
rect 30683 36841 30956 36881
rect 30583 36764 30956 36841
rect 30583 36723 30855 36764
rect 30583 36677 30637 36723
rect 30683 36718 30855 36723
rect 30901 36718 30956 36764
rect 30683 36677 30956 36718
rect 30583 36601 30956 36677
rect 30583 36560 30855 36601
rect 30583 36514 30637 36560
rect 30683 36555 30855 36560
rect 30901 36555 30956 36601
rect 30683 36514 30956 36555
rect 30583 36438 30956 36514
rect 30583 36397 30855 36438
rect 30583 36351 30637 36397
rect 30683 36392 30855 36397
rect 30901 36392 30956 36438
rect 30683 36351 30956 36392
rect 30583 36274 30956 36351
rect 30583 36234 30855 36274
rect 30583 36188 30637 36234
rect 30683 36228 30855 36234
rect 30901 36228 30956 36274
rect 30683 36188 30956 36228
rect 30583 36065 30956 36188
rect 54168 36881 54223 36927
rect 54269 36887 54540 36927
rect 54269 36881 54440 36887
rect 54168 36841 54440 36881
rect 54486 36841 54540 36887
rect 36348 36150 36861 36196
rect 36348 36104 36489 36150
rect 36723 36104 36861 36150
rect 30583 36061 30802 36065
rect 36348 36058 36861 36104
rect 39007 36150 39321 36207
rect 39007 36104 39062 36150
rect 39108 36104 39220 36150
rect 39266 36104 39321 36150
rect 39007 36047 39321 36104
rect 45564 36314 48566 36371
rect 45564 36268 45619 36314
rect 45665 36268 45777 36314
rect 45823 36268 45935 36314
rect 45981 36268 46093 36314
rect 46139 36268 46251 36314
rect 46297 36268 46409 36314
rect 46455 36268 46568 36314
rect 46614 36268 46726 36314
rect 46772 36268 46884 36314
rect 46930 36268 47042 36314
rect 47088 36268 47200 36314
rect 47246 36268 47358 36314
rect 47404 36268 47516 36314
rect 47562 36268 47675 36314
rect 47721 36268 47833 36314
rect 47879 36268 47991 36314
rect 48037 36268 48149 36314
rect 48195 36268 48307 36314
rect 48353 36268 48465 36314
rect 48511 36268 48566 36314
rect 54168 36723 54540 36841
rect 54168 36677 54440 36723
rect 54486 36677 54540 36723
rect 54168 36560 54540 36677
rect 54168 36514 54440 36560
rect 54486 36514 54540 36560
rect 54168 36438 54540 36514
rect 54168 36392 54223 36438
rect 54269 36397 54540 36438
rect 54269 36392 54440 36397
rect 54168 36351 54440 36392
rect 54486 36351 54540 36397
rect 45564 36196 48566 36268
rect 45564 36150 48766 36196
rect 54168 36274 54540 36351
rect 54168 36228 54223 36274
rect 54269 36234 54540 36274
rect 54269 36228 54440 36234
rect 54168 36188 54440 36228
rect 54486 36188 54540 36234
rect 45564 36104 45619 36150
rect 45665 36104 45777 36150
rect 45823 36104 45935 36150
rect 45981 36104 46093 36150
rect 46139 36104 46251 36150
rect 46297 36104 46409 36150
rect 46455 36104 46568 36150
rect 46614 36104 46726 36150
rect 46772 36104 46884 36150
rect 46930 36104 47042 36150
rect 47088 36104 47200 36150
rect 47246 36104 47358 36150
rect 47404 36104 47516 36150
rect 47562 36104 47675 36150
rect 47721 36104 47833 36150
rect 47879 36104 47991 36150
rect 48037 36104 48149 36150
rect 48195 36104 48307 36150
rect 48353 36104 48465 36150
rect 48511 36104 48766 36150
rect 45564 36058 48766 36104
rect 54168 36065 54540 36188
rect 54321 36061 54540 36065
rect 45564 36047 48566 36058
<< mvpsubdiffcont >>
rect 33044 65863 33090 65909
rect 33202 65863 33248 65909
rect 33360 65863 33406 65909
rect 33518 65863 33564 65909
rect 33677 65863 33723 65909
rect 33835 65863 33881 65909
rect 33993 65863 34039 65909
rect 34151 65863 34197 65909
rect 34309 65863 34355 65909
rect 34467 65863 34513 65909
rect 34625 65863 34671 65909
rect 34783 65863 34829 65909
rect 40117 65863 40163 65909
rect 40275 65863 40321 65909
rect 40433 65863 40479 65909
rect 40591 65863 40637 65909
rect 40750 65863 40796 65909
rect 40908 65863 40954 65909
rect 41066 65863 41112 65909
rect 41224 65863 41270 65909
rect 41382 65863 41428 65909
rect 41540 65863 41586 65909
rect 41698 65863 41744 65909
rect 41856 65863 41902 65909
rect 28810 65676 28856 65722
rect 28810 65512 28856 65558
rect 28810 65349 28856 65395
rect 28810 65186 28856 65232
rect 28810 65022 28856 65068
rect 44514 65863 44560 65909
rect 44672 65863 44718 65909
rect 44830 65863 44876 65909
rect 50129 65863 50175 65909
rect 50287 65863 50333 65909
rect 50445 65863 50491 65909
rect 50603 65863 50649 65909
rect 50762 65863 50808 65909
rect 50920 65863 50966 65909
rect 51078 65863 51124 65909
rect 51236 65863 51282 65909
rect 51394 65863 51440 65909
rect 51552 65863 51598 65909
rect 51710 65863 51756 65909
rect 51868 65863 51914 65909
rect 28810 64820 28856 64866
rect 28810 64657 28856 64703
rect 28810 64494 28856 64540
rect 28810 64331 28856 64377
rect 28810 64167 28856 64213
rect 37957 64904 38473 64950
rect 40836 64904 40882 64950
rect 40994 64904 41040 64950
rect 41152 64904 41198 64950
rect 41310 64904 41356 64950
rect 41469 64904 41515 64950
rect 41627 64904 41673 64950
rect 41785 64904 41831 64950
rect 41943 64904 41989 64950
rect 42101 64904 42147 64950
rect 42259 64904 42305 64950
rect 42418 64904 42464 64950
rect 42576 64904 42622 64950
rect 42734 64904 42780 64950
rect 42892 64904 42938 64950
rect 56267 65676 56313 65722
rect 56267 65512 56313 65558
rect 56267 65349 56313 65395
rect 56267 65186 56313 65232
rect 56267 65022 56313 65068
rect 28810 64004 28856 64050
rect 28810 63841 28856 63887
rect 28810 63677 28856 63723
rect 28810 63514 28856 63560
rect 28810 63351 28856 63397
rect 28810 63188 28856 63234
rect 34916 64004 34962 64050
rect 50160 64004 50206 64050
rect 56267 64820 56313 64866
rect 56267 64657 56313 64703
rect 56267 64494 56313 64540
rect 56267 64331 56313 64377
rect 56267 64167 56313 64213
rect 56267 64004 56313 64050
rect 28810 63020 28856 63066
rect 28810 62857 28856 62903
rect 28810 62694 28856 62740
rect 28810 62531 28856 62577
rect 28810 62367 28856 62413
rect 37957 63104 38473 63150
rect 40836 63104 40882 63150
rect 40994 63104 41040 63150
rect 41152 63104 41198 63150
rect 41310 63104 41356 63150
rect 41469 63104 41515 63150
rect 41627 63104 41673 63150
rect 41785 63104 41831 63150
rect 41943 63104 41989 63150
rect 42101 63104 42147 63150
rect 42259 63104 42305 63150
rect 42418 63104 42464 63150
rect 42576 63104 42622 63150
rect 42734 63104 42780 63150
rect 42892 63104 42938 63150
rect 56267 63841 56313 63887
rect 56267 63677 56313 63723
rect 56267 63514 56313 63560
rect 56267 63351 56313 63397
rect 56267 63188 56313 63234
rect 28810 62204 28856 62250
rect 28810 62041 28856 62087
rect 28810 61877 28856 61923
rect 28810 61714 28856 61760
rect 28810 61551 28856 61597
rect 28810 61388 28856 61434
rect 34916 62204 34962 62250
rect 50160 62204 50206 62250
rect 56267 63020 56313 63066
rect 56267 62857 56313 62903
rect 56267 62694 56313 62740
rect 56267 62531 56313 62577
rect 56267 62367 56313 62413
rect 56267 62204 56313 62250
rect 28810 61220 28856 61266
rect 28810 61057 28856 61103
rect 28810 60894 28856 60940
rect 28810 60731 28856 60777
rect 28810 60567 28856 60613
rect 37957 61304 38473 61350
rect 40836 61304 40882 61350
rect 40994 61304 41040 61350
rect 41152 61304 41198 61350
rect 41310 61304 41356 61350
rect 41469 61304 41515 61350
rect 41627 61304 41673 61350
rect 41785 61304 41831 61350
rect 41943 61304 41989 61350
rect 42101 61304 42147 61350
rect 42259 61304 42305 61350
rect 42418 61304 42464 61350
rect 42576 61304 42622 61350
rect 42734 61304 42780 61350
rect 42892 61304 42938 61350
rect 56267 62041 56313 62087
rect 56267 61877 56313 61923
rect 56267 61714 56313 61760
rect 56267 61551 56313 61597
rect 56267 61388 56313 61434
rect 28810 60404 28856 60450
rect 28810 60241 28856 60287
rect 28810 60077 28856 60123
rect 28810 59914 28856 59960
rect 28810 59751 28856 59797
rect 28810 59588 28856 59634
rect 34916 60404 34962 60450
rect 50160 60404 50206 60450
rect 56267 61220 56313 61266
rect 56267 61057 56313 61103
rect 56267 60894 56313 60940
rect 56267 60731 56313 60777
rect 56267 60567 56313 60613
rect 56267 60404 56313 60450
rect 28810 59420 28856 59466
rect 28810 59257 28856 59303
rect 28810 59094 28856 59140
rect 28810 58931 28856 58977
rect 28810 58767 28856 58813
rect 37957 59504 38473 59550
rect 40836 59504 40882 59550
rect 40994 59504 41040 59550
rect 41152 59504 41198 59550
rect 41310 59504 41356 59550
rect 41469 59504 41515 59550
rect 41627 59504 41673 59550
rect 41785 59504 41831 59550
rect 41943 59504 41989 59550
rect 42101 59504 42147 59550
rect 42259 59504 42305 59550
rect 42418 59504 42464 59550
rect 42576 59504 42622 59550
rect 42734 59504 42780 59550
rect 42892 59504 42938 59550
rect 56267 60241 56313 60287
rect 56267 60077 56313 60123
rect 56267 59914 56313 59960
rect 56267 59751 56313 59797
rect 56267 59588 56313 59634
rect 28810 58604 28856 58650
rect 28810 58441 28856 58487
rect 28810 58277 28856 58323
rect 28810 58114 28856 58160
rect 28810 57951 28856 57997
rect 28810 57788 28856 57834
rect 34916 58604 34962 58650
rect 50160 58604 50206 58650
rect 56267 59420 56313 59466
rect 56267 59257 56313 59303
rect 56267 59094 56313 59140
rect 56267 58931 56313 58977
rect 56267 58767 56313 58813
rect 56267 58604 56313 58650
rect 28810 57620 28856 57666
rect 28810 57457 28856 57503
rect 28810 57294 28856 57340
rect 28810 57131 28856 57177
rect 28810 56967 28856 57013
rect 37957 57704 38473 57750
rect 40836 57704 40882 57750
rect 40994 57704 41040 57750
rect 41152 57704 41198 57750
rect 41310 57704 41356 57750
rect 41469 57704 41515 57750
rect 41627 57704 41673 57750
rect 41785 57704 41831 57750
rect 41943 57704 41989 57750
rect 42101 57704 42147 57750
rect 42259 57704 42305 57750
rect 42418 57704 42464 57750
rect 42576 57704 42622 57750
rect 42734 57704 42780 57750
rect 42892 57704 42938 57750
rect 56267 58441 56313 58487
rect 56267 58277 56313 58323
rect 56267 58114 56313 58160
rect 56267 57951 56313 57997
rect 56267 57788 56313 57834
rect 28810 56804 28856 56850
rect 28810 56641 28856 56687
rect 28810 56477 28856 56523
rect 28810 56314 28856 56360
rect 28810 56151 28856 56197
rect 28810 55988 28856 56034
rect 34916 56804 34962 56850
rect 50160 56804 50206 56850
rect 56267 57620 56313 57666
rect 56267 57457 56313 57503
rect 56267 57294 56313 57340
rect 56267 57131 56313 57177
rect 56267 56967 56313 57013
rect 56267 56804 56313 56850
rect 28810 55820 28856 55866
rect 28810 55657 28856 55703
rect 28810 55494 28856 55540
rect 28810 55331 28856 55377
rect 28810 55167 28856 55213
rect 37957 55904 38473 55950
rect 40836 55904 40882 55950
rect 40994 55904 41040 55950
rect 41152 55904 41198 55950
rect 41310 55904 41356 55950
rect 41469 55904 41515 55950
rect 41627 55904 41673 55950
rect 41785 55904 41831 55950
rect 41943 55904 41989 55950
rect 42101 55904 42147 55950
rect 42259 55904 42305 55950
rect 42418 55904 42464 55950
rect 42576 55904 42622 55950
rect 42734 55904 42780 55950
rect 42892 55904 42938 55950
rect 56267 56641 56313 56687
rect 56267 56477 56313 56523
rect 56267 56314 56313 56360
rect 56267 56151 56313 56197
rect 56267 55988 56313 56034
rect 28810 55004 28856 55050
rect 28810 54841 28856 54887
rect 28810 54677 28856 54723
rect 28810 54514 28856 54560
rect 28810 54351 28856 54397
rect 28810 54188 28856 54234
rect 34916 55004 34962 55050
rect 50160 55004 50206 55050
rect 56267 55820 56313 55866
rect 56267 55657 56313 55703
rect 56267 55494 56313 55540
rect 56267 55331 56313 55377
rect 56267 55167 56313 55213
rect 56267 55004 56313 55050
rect 28810 54020 28856 54066
rect 28810 53857 28856 53903
rect 28810 53694 28856 53740
rect 28810 53531 28856 53577
rect 28810 53367 28856 53413
rect 37957 54104 38473 54150
rect 40836 54104 40882 54150
rect 40994 54104 41040 54150
rect 41152 54104 41198 54150
rect 41310 54104 41356 54150
rect 41469 54104 41515 54150
rect 41627 54104 41673 54150
rect 41785 54104 41831 54150
rect 41943 54104 41989 54150
rect 42101 54104 42147 54150
rect 42259 54104 42305 54150
rect 42418 54104 42464 54150
rect 42576 54104 42622 54150
rect 42734 54104 42780 54150
rect 42892 54104 42938 54150
rect 56267 54841 56313 54887
rect 56267 54677 56313 54723
rect 56267 54514 56313 54560
rect 56267 54351 56313 54397
rect 56267 54188 56313 54234
rect 28810 53204 28856 53250
rect 28810 53041 28856 53087
rect 28810 52877 28856 52923
rect 28810 52714 28856 52760
rect 28810 52551 28856 52597
rect 28810 52388 28856 52434
rect 34916 53204 34962 53250
rect 50160 53204 50206 53250
rect 56267 54020 56313 54066
rect 56267 53857 56313 53903
rect 56267 53694 56313 53740
rect 56267 53531 56313 53577
rect 56267 53367 56313 53413
rect 56267 53204 56313 53250
rect 28810 52220 28856 52266
rect 28810 52057 28856 52103
rect 28810 51894 28856 51940
rect 28810 51731 28856 51777
rect 28810 51567 28856 51613
rect 37957 52304 38473 52350
rect 40836 52304 40882 52350
rect 40994 52304 41040 52350
rect 41152 52304 41198 52350
rect 41310 52304 41356 52350
rect 41469 52304 41515 52350
rect 41627 52304 41673 52350
rect 41785 52304 41831 52350
rect 41943 52304 41989 52350
rect 42101 52304 42147 52350
rect 42259 52304 42305 52350
rect 42418 52304 42464 52350
rect 42576 52304 42622 52350
rect 42734 52304 42780 52350
rect 42892 52304 42938 52350
rect 56267 53041 56313 53087
rect 56267 52877 56313 52923
rect 56267 52714 56313 52760
rect 56267 52551 56313 52597
rect 56267 52388 56313 52434
rect 28810 51404 28856 51450
rect 28810 51241 28856 51287
rect 28810 51077 28856 51123
rect 28810 50914 28856 50960
rect 28810 50751 28856 50797
rect 28810 50588 28856 50634
rect 34916 51404 34962 51450
rect 50160 51404 50206 51450
rect 56267 52220 56313 52266
rect 56267 52057 56313 52103
rect 56267 51894 56313 51940
rect 56267 51731 56313 51777
rect 56267 51567 56313 51613
rect 56267 51404 56313 51450
rect 28810 50420 28856 50466
rect 28810 50257 28856 50303
rect 28810 50094 28856 50140
rect 28810 49931 28856 49977
rect 28810 49767 28856 49813
rect 37957 50504 38473 50550
rect 40836 50504 40882 50550
rect 40994 50504 41040 50550
rect 41152 50504 41198 50550
rect 41310 50504 41356 50550
rect 41469 50504 41515 50550
rect 41627 50504 41673 50550
rect 41785 50504 41831 50550
rect 41943 50504 41989 50550
rect 42101 50504 42147 50550
rect 42259 50504 42305 50550
rect 42418 50504 42464 50550
rect 42576 50504 42622 50550
rect 42734 50504 42780 50550
rect 42892 50504 42938 50550
rect 56267 51241 56313 51287
rect 56267 51077 56313 51123
rect 56267 50914 56313 50960
rect 56267 50751 56313 50797
rect 56267 50588 56313 50634
rect 28810 49604 28856 49650
rect 28810 49441 28856 49487
rect 28810 49277 28856 49323
rect 28810 49114 28856 49160
rect 28810 48951 28856 48997
rect 28810 48788 28856 48834
rect 34916 49604 34962 49650
rect 50160 49604 50206 49650
rect 56267 50420 56313 50466
rect 56267 50257 56313 50303
rect 56267 50094 56313 50140
rect 56267 49931 56313 49977
rect 56267 49767 56313 49813
rect 56267 49604 56313 49650
rect 28810 48620 28856 48666
rect 28810 48457 28856 48503
rect 28810 48294 28856 48340
rect 28810 48131 28856 48177
rect 28810 47967 28856 48013
rect 37957 48704 38473 48750
rect 40836 48704 40882 48750
rect 40994 48704 41040 48750
rect 41152 48704 41198 48750
rect 41310 48704 41356 48750
rect 41469 48704 41515 48750
rect 41627 48704 41673 48750
rect 41785 48704 41831 48750
rect 41943 48704 41989 48750
rect 42101 48704 42147 48750
rect 42259 48704 42305 48750
rect 42418 48704 42464 48750
rect 42576 48704 42622 48750
rect 42734 48704 42780 48750
rect 42892 48704 42938 48750
rect 56267 49441 56313 49487
rect 56267 49277 56313 49323
rect 56267 49114 56313 49160
rect 56267 48951 56313 48997
rect 56267 48788 56313 48834
rect 28810 47804 28856 47850
rect 28810 47641 28856 47687
rect 28810 47477 28856 47523
rect 28810 47314 28856 47360
rect 28810 47151 28856 47197
rect 28810 46988 28856 47034
rect 34916 47804 34962 47850
rect 50160 47804 50206 47850
rect 56267 48620 56313 48666
rect 56267 48457 56313 48503
rect 56267 48294 56313 48340
rect 56267 48131 56313 48177
rect 56267 47967 56313 48013
rect 56267 47804 56313 47850
rect 28810 46820 28856 46866
rect 28810 46657 28856 46703
rect 28810 46494 28856 46540
rect 28810 46331 28856 46377
rect 28810 46167 28856 46213
rect 37957 46904 38473 46950
rect 40836 46904 40882 46950
rect 40994 46904 41040 46950
rect 41152 46904 41198 46950
rect 41310 46904 41356 46950
rect 41469 46904 41515 46950
rect 41627 46904 41673 46950
rect 41785 46904 41831 46950
rect 41943 46904 41989 46950
rect 42101 46904 42147 46950
rect 42259 46904 42305 46950
rect 42418 46904 42464 46950
rect 42576 46904 42622 46950
rect 42734 46904 42780 46950
rect 42892 46904 42938 46950
rect 56267 47641 56313 47687
rect 56267 47477 56313 47523
rect 56267 47314 56313 47360
rect 56267 47151 56313 47197
rect 56267 46988 56313 47034
rect 28810 46004 28856 46050
rect 28810 45841 28856 45887
rect 28810 45677 28856 45723
rect 28810 45514 28856 45560
rect 28810 45351 28856 45397
rect 28810 45188 28856 45234
rect 34916 46004 34962 46050
rect 50160 46004 50206 46050
rect 56267 46820 56313 46866
rect 56267 46657 56313 46703
rect 56267 46494 56313 46540
rect 56267 46331 56313 46377
rect 56267 46167 56313 46213
rect 56267 46004 56313 46050
rect 28810 45020 28856 45066
rect 28810 44857 28856 44903
rect 28810 44694 28856 44740
rect 28810 44531 28856 44577
rect 28810 44367 28856 44413
rect 37957 45104 38473 45150
rect 40836 45104 40882 45150
rect 40994 45104 41040 45150
rect 41152 45104 41198 45150
rect 41310 45104 41356 45150
rect 41469 45104 41515 45150
rect 41627 45104 41673 45150
rect 41785 45104 41831 45150
rect 41943 45104 41989 45150
rect 42101 45104 42147 45150
rect 42259 45104 42305 45150
rect 42418 45104 42464 45150
rect 42576 45104 42622 45150
rect 42734 45104 42780 45150
rect 42892 45104 42938 45150
rect 56267 45841 56313 45887
rect 56267 45677 56313 45723
rect 56267 45514 56313 45560
rect 56267 45351 56313 45397
rect 56267 45188 56313 45234
rect 28810 44204 28856 44250
rect 28810 44041 28856 44087
rect 28810 43877 28856 43923
rect 28810 43714 28856 43760
rect 28810 43551 28856 43597
rect 28810 43388 28856 43434
rect 34916 44204 34962 44250
rect 50160 44204 50206 44250
rect 56267 45020 56313 45066
rect 56267 44857 56313 44903
rect 56267 44694 56313 44740
rect 56267 44531 56313 44577
rect 56267 44367 56313 44413
rect 56267 44204 56313 44250
rect 28810 43220 28856 43266
rect 28810 43057 28856 43103
rect 28810 42894 28856 42940
rect 28810 42731 28856 42777
rect 28810 42567 28856 42613
rect 37957 43304 38473 43350
rect 40836 43304 40882 43350
rect 40994 43304 41040 43350
rect 41152 43304 41198 43350
rect 41310 43304 41356 43350
rect 41469 43304 41515 43350
rect 41627 43304 41673 43350
rect 41785 43304 41831 43350
rect 41943 43304 41989 43350
rect 42101 43304 42147 43350
rect 42259 43304 42305 43350
rect 42418 43304 42464 43350
rect 42576 43304 42622 43350
rect 42734 43304 42780 43350
rect 42892 43304 42938 43350
rect 56267 44041 56313 44087
rect 56267 43877 56313 43923
rect 56267 43714 56313 43760
rect 56267 43551 56313 43597
rect 56267 43388 56313 43434
rect 28810 42404 28856 42450
rect 28810 42241 28856 42287
rect 28810 42077 28856 42123
rect 28810 41914 28856 41960
rect 28810 41751 28856 41797
rect 28810 41588 28856 41634
rect 34916 42404 34962 42450
rect 50160 42404 50206 42450
rect 56267 43220 56313 43266
rect 56267 43057 56313 43103
rect 56267 42894 56313 42940
rect 56267 42731 56313 42777
rect 56267 42567 56313 42613
rect 56267 42404 56313 42450
rect 28810 41420 28856 41466
rect 28810 41257 28856 41303
rect 28810 41094 28856 41140
rect 28810 40931 28856 40977
rect 28810 40767 28856 40813
rect 37957 41504 38473 41550
rect 40836 41504 40882 41550
rect 40994 41504 41040 41550
rect 41152 41504 41198 41550
rect 41310 41504 41356 41550
rect 41469 41504 41515 41550
rect 41627 41504 41673 41550
rect 41785 41504 41831 41550
rect 41943 41504 41989 41550
rect 42101 41504 42147 41550
rect 42259 41504 42305 41550
rect 42418 41504 42464 41550
rect 42576 41504 42622 41550
rect 42734 41504 42780 41550
rect 42892 41504 42938 41550
rect 56267 42241 56313 42287
rect 56267 42077 56313 42123
rect 56267 41914 56313 41960
rect 56267 41751 56313 41797
rect 56267 41588 56313 41634
rect 28810 40604 28856 40650
rect 28810 40441 28856 40487
rect 28810 40277 28856 40323
rect 28810 40114 28856 40160
rect 28810 39951 28856 39997
rect 28810 39788 28856 39834
rect 34916 40604 34962 40650
rect 50160 40604 50206 40650
rect 56267 41420 56313 41466
rect 56267 41257 56313 41303
rect 56267 41094 56313 41140
rect 56267 40931 56313 40977
rect 56267 40767 56313 40813
rect 56267 40604 56313 40650
rect 28810 39620 28856 39666
rect 28810 39457 28856 39503
rect 28810 39294 28856 39340
rect 28810 39131 28856 39177
rect 28810 38967 28856 39013
rect 37957 39704 38473 39750
rect 40836 39704 40882 39750
rect 40994 39704 41040 39750
rect 41152 39704 41198 39750
rect 41310 39704 41356 39750
rect 41469 39704 41515 39750
rect 41627 39704 41673 39750
rect 41785 39704 41831 39750
rect 41943 39704 41989 39750
rect 42101 39704 42147 39750
rect 42259 39704 42305 39750
rect 42418 39704 42464 39750
rect 42576 39704 42622 39750
rect 42734 39704 42780 39750
rect 42892 39704 42938 39750
rect 56267 40441 56313 40487
rect 56267 40277 56313 40323
rect 56267 40114 56313 40160
rect 56267 39951 56313 39997
rect 56267 39788 56313 39834
rect 28810 38804 28856 38850
rect 28810 38641 28856 38687
rect 28810 38477 28856 38523
rect 28810 38314 28856 38360
rect 28810 38151 28856 38197
rect 28810 37988 28856 38034
rect 34916 38804 34962 38850
rect 50160 38804 50206 38850
rect 56267 39620 56313 39666
rect 56267 39457 56313 39503
rect 56267 39294 56313 39340
rect 56267 39131 56313 39177
rect 56267 38967 56313 39013
rect 56267 38804 56313 38850
rect 28810 37820 28856 37866
rect 28810 37657 28856 37703
rect 28810 37494 28856 37540
rect 28810 37331 28856 37377
rect 28810 37167 28856 37213
rect 37957 37904 38473 37950
rect 40836 37904 40882 37950
rect 40994 37904 41040 37950
rect 41152 37904 41198 37950
rect 41310 37904 41356 37950
rect 41469 37904 41515 37950
rect 41627 37904 41673 37950
rect 41785 37904 41831 37950
rect 41943 37904 41989 37950
rect 42101 37904 42147 37950
rect 42259 37904 42305 37950
rect 42418 37904 42464 37950
rect 42576 37904 42622 37950
rect 42734 37904 42780 37950
rect 42892 37904 42938 37950
rect 56267 38641 56313 38687
rect 56267 38477 56313 38523
rect 56267 38314 56313 38360
rect 56267 38151 56313 38197
rect 56267 37988 56313 38034
rect 28810 37004 28856 37050
rect 28810 36841 28856 36887
rect 28810 36677 28856 36723
rect 28810 36514 28856 36560
rect 28810 36351 28856 36397
rect 28810 36188 28856 36234
rect 34916 37004 34962 37050
rect 50160 37004 50206 37050
rect 56267 37820 56313 37866
rect 56267 37657 56313 37703
rect 56267 37494 56313 37540
rect 56267 37331 56313 37377
rect 56267 37167 56313 37213
rect 56267 37004 56313 37050
rect 37957 36104 38473 36150
rect 40836 36104 40882 36150
rect 40994 36104 41040 36150
rect 41152 36104 41198 36150
rect 41310 36104 41356 36150
rect 41469 36104 41515 36150
rect 41627 36104 41673 36150
rect 41785 36104 41831 36150
rect 41943 36104 41989 36150
rect 42101 36104 42147 36150
rect 42259 36104 42305 36150
rect 42418 36104 42464 36150
rect 42576 36104 42622 36150
rect 42734 36104 42780 36150
rect 42892 36104 42938 36150
rect 56267 36841 56313 36887
rect 56267 36677 56313 36723
rect 56267 36514 56313 36560
rect 56267 36351 56313 36397
rect 56267 36188 56313 36234
rect 28639 3860 28685 3906
rect 28755 3860 28801 3906
rect 28871 3860 28917 3906
rect 28987 3860 29033 3906
rect 29103 3860 29149 3906
rect 29219 3860 29265 3906
rect 29335 3860 29381 3906
rect 29451 3860 29497 3906
rect 29567 3860 29613 3906
rect 29683 3860 29729 3906
rect 29799 3860 29845 3906
rect 29915 3860 29961 3906
rect 30031 3860 30077 3906
rect 30147 3860 30193 3906
rect 30263 3860 30309 3906
rect 30379 3860 30425 3906
rect 30495 3860 30541 3906
rect 30611 3860 30657 3906
rect 30727 3860 30773 3906
rect 30843 3860 30889 3906
rect 30959 3860 31005 3906
rect 31075 3860 31121 3906
rect 31191 3860 31237 3906
rect 31307 3860 31353 3906
rect 31423 3860 31469 3906
rect 31539 3860 31585 3906
rect 31655 3860 31701 3906
rect 31771 3860 31817 3906
rect 31887 3860 31933 3906
rect 32003 3860 32049 3906
rect 32119 3860 32165 3906
rect 32235 3860 32281 3906
rect 32351 3860 32397 3906
rect 32467 3860 32513 3906
rect 32583 3860 32629 3906
rect 32699 3860 32745 3906
rect 32815 3860 32861 3906
rect 32931 3860 32977 3906
rect 33047 3860 33093 3906
rect 33163 3860 33209 3906
rect 33279 3860 33325 3906
rect 33395 3860 33441 3906
rect 33511 3860 33557 3906
rect 33627 3860 33673 3906
rect 33743 3860 33789 3906
rect 33859 3860 33905 3906
rect 33975 3860 34021 3906
rect 34091 3860 34137 3906
rect 34207 3860 34253 3906
rect 34323 3860 34369 3906
rect 34439 3860 34485 3906
rect 34555 3860 34601 3906
rect 34671 3860 34717 3906
rect 34787 3860 34833 3906
rect 34903 3860 34949 3906
rect 35019 3860 35065 3906
rect 35135 3860 35181 3906
rect 35251 3860 35297 3906
rect 35367 3860 35413 3906
rect 35483 3860 35529 3906
rect 35599 3860 35645 3906
rect 35715 3860 35761 3906
rect 35831 3860 35877 3906
rect 35947 3860 35993 3906
rect 36063 3860 36109 3906
rect 36179 3860 36225 3906
rect 36295 3860 36341 3906
rect 36411 3860 36457 3906
rect 36527 3860 36573 3906
rect 36643 3860 36689 3906
rect 36759 3860 36805 3906
rect 36875 3860 36921 3906
rect 36991 3860 37037 3906
rect 37107 3860 37153 3906
rect 37223 3860 37269 3906
rect 37339 3860 37385 3906
rect 37455 3860 37501 3906
rect 37571 3860 37617 3906
rect 37687 3860 37733 3906
rect 37803 3860 37849 3906
rect 37919 3860 37965 3906
rect 38035 3860 38081 3906
rect 38151 3860 38197 3906
rect 38267 3860 38313 3906
rect 38383 3860 38429 3906
rect 38499 3860 38545 3906
rect 38615 3860 38661 3906
rect 38731 3860 38777 3906
rect 38847 3860 38893 3906
rect 38963 3860 39009 3906
rect 39079 3860 39125 3906
rect 39195 3860 39241 3906
rect 39311 3860 39357 3906
rect 39427 3860 39473 3906
rect 39543 3860 39589 3906
rect 39659 3860 39705 3906
rect 39775 3860 39821 3906
rect 39891 3860 39937 3906
rect 40007 3860 40053 3906
rect 40123 3860 40169 3906
rect 28639 3744 28685 3790
rect 28755 3744 28801 3790
rect 28871 3744 28917 3790
rect 28987 3744 29033 3790
rect 29103 3744 29149 3790
rect 29219 3744 29265 3790
rect 29335 3744 29381 3790
rect 29451 3744 29497 3790
rect 29567 3744 29613 3790
rect 29683 3744 29729 3790
rect 29799 3744 29845 3790
rect 29915 3744 29961 3790
rect 30031 3744 30077 3790
rect 30147 3744 30193 3790
rect 30263 3744 30309 3790
rect 30379 3744 30425 3790
rect 30495 3744 30541 3790
rect 30611 3744 30657 3790
rect 30727 3744 30773 3790
rect 30843 3744 30889 3790
rect 30959 3744 31005 3790
rect 31075 3744 31121 3790
rect 31191 3744 31237 3790
rect 31307 3744 31353 3790
rect 31423 3744 31469 3790
rect 31539 3744 31585 3790
rect 31655 3744 31701 3790
rect 31771 3744 31817 3790
rect 31887 3744 31933 3790
rect 32003 3744 32049 3790
rect 32119 3744 32165 3790
rect 32235 3744 32281 3790
rect 32351 3744 32397 3790
rect 32467 3744 32513 3790
rect 32583 3744 32629 3790
rect 32699 3744 32745 3790
rect 32815 3744 32861 3790
rect 32931 3744 32977 3790
rect 33047 3744 33093 3790
rect 33163 3744 33209 3790
rect 33279 3744 33325 3790
rect 33395 3744 33441 3790
rect 33511 3744 33557 3790
rect 33627 3744 33673 3790
rect 33743 3744 33789 3790
rect 33859 3744 33905 3790
rect 33975 3744 34021 3790
rect 34091 3744 34137 3790
rect 34207 3744 34253 3790
rect 34323 3744 34369 3790
rect 34439 3744 34485 3790
rect 34555 3744 34601 3790
rect 34671 3744 34717 3790
rect 34787 3744 34833 3790
rect 34903 3744 34949 3790
rect 35019 3744 35065 3790
rect 35135 3744 35181 3790
rect 35251 3744 35297 3790
rect 35367 3744 35413 3790
rect 35483 3744 35529 3790
rect 35599 3744 35645 3790
rect 35715 3744 35761 3790
rect 35831 3744 35877 3790
rect 35947 3744 35993 3790
rect 36063 3744 36109 3790
rect 36179 3744 36225 3790
rect 36295 3744 36341 3790
rect 36411 3744 36457 3790
rect 36527 3744 36573 3790
rect 36643 3744 36689 3790
rect 36759 3744 36805 3790
rect 36875 3744 36921 3790
rect 36991 3744 37037 3790
rect 37107 3744 37153 3790
rect 37223 3744 37269 3790
rect 37339 3744 37385 3790
rect 37455 3744 37501 3790
rect 37571 3744 37617 3790
rect 37687 3744 37733 3790
rect 37803 3744 37849 3790
rect 37919 3744 37965 3790
rect 38035 3744 38081 3790
rect 38151 3744 38197 3790
rect 38267 3744 38313 3790
rect 38383 3744 38429 3790
rect 38499 3744 38545 3790
rect 38615 3744 38661 3790
rect 38731 3744 38777 3790
rect 38847 3744 38893 3790
rect 38963 3744 39009 3790
rect 39079 3744 39125 3790
rect 39195 3744 39241 3790
rect 39311 3744 39357 3790
rect 39427 3744 39473 3790
rect 39543 3744 39589 3790
rect 39659 3744 39705 3790
rect 39775 3744 39821 3790
rect 39891 3744 39937 3790
rect 40007 3744 40053 3790
rect 40123 3744 40169 3790
rect 28639 3628 28685 3674
rect 28755 3628 28801 3674
rect 28871 3628 28917 3674
rect 28987 3628 29033 3674
rect 29103 3628 29149 3674
rect 29219 3628 29265 3674
rect 29335 3628 29381 3674
rect 29451 3628 29497 3674
rect 29567 3628 29613 3674
rect 29683 3628 29729 3674
rect 29799 3628 29845 3674
rect 29915 3628 29961 3674
rect 30031 3628 30077 3674
rect 30147 3628 30193 3674
rect 30263 3628 30309 3674
rect 30379 3628 30425 3674
rect 30495 3628 30541 3674
rect 30611 3628 30657 3674
rect 30727 3628 30773 3674
rect 30843 3628 30889 3674
rect 30959 3628 31005 3674
rect 31075 3628 31121 3674
rect 31191 3628 31237 3674
rect 31307 3628 31353 3674
rect 31423 3628 31469 3674
rect 31539 3628 31585 3674
rect 31655 3628 31701 3674
rect 31771 3628 31817 3674
rect 31887 3628 31933 3674
rect 32003 3628 32049 3674
rect 32119 3628 32165 3674
rect 32235 3628 32281 3674
rect 32351 3628 32397 3674
rect 32467 3628 32513 3674
rect 32583 3628 32629 3674
rect 32699 3628 32745 3674
rect 32815 3628 32861 3674
rect 32931 3628 32977 3674
rect 33047 3628 33093 3674
rect 33163 3628 33209 3674
rect 33279 3628 33325 3674
rect 33395 3628 33441 3674
rect 33511 3628 33557 3674
rect 33627 3628 33673 3674
rect 33743 3628 33789 3674
rect 33859 3628 33905 3674
rect 33975 3628 34021 3674
rect 34091 3628 34137 3674
rect 34207 3628 34253 3674
rect 34323 3628 34369 3674
rect 34439 3628 34485 3674
rect 34555 3628 34601 3674
rect 34671 3628 34717 3674
rect 34787 3628 34833 3674
rect 34903 3628 34949 3674
rect 35019 3628 35065 3674
rect 35135 3628 35181 3674
rect 35251 3628 35297 3674
rect 35367 3628 35413 3674
rect 35483 3628 35529 3674
rect 35599 3628 35645 3674
rect 35715 3628 35761 3674
rect 35831 3628 35877 3674
rect 35947 3628 35993 3674
rect 36063 3628 36109 3674
rect 36179 3628 36225 3674
rect 36295 3628 36341 3674
rect 36411 3628 36457 3674
rect 36527 3628 36573 3674
rect 36643 3628 36689 3674
rect 36759 3628 36805 3674
rect 36875 3628 36921 3674
rect 36991 3628 37037 3674
rect 37107 3628 37153 3674
rect 37223 3628 37269 3674
rect 37339 3628 37385 3674
rect 37455 3628 37501 3674
rect 37571 3628 37617 3674
rect 37687 3628 37733 3674
rect 37803 3628 37849 3674
rect 37919 3628 37965 3674
rect 38035 3628 38081 3674
rect 38151 3628 38197 3674
rect 38267 3628 38313 3674
rect 38383 3628 38429 3674
rect 38499 3628 38545 3674
rect 38615 3628 38661 3674
rect 38731 3628 38777 3674
rect 38847 3628 38893 3674
rect 38963 3628 39009 3674
rect 39079 3628 39125 3674
rect 39195 3628 39241 3674
rect 39311 3628 39357 3674
rect 39427 3628 39473 3674
rect 39543 3628 39589 3674
rect 39659 3628 39705 3674
rect 39775 3628 39821 3674
rect 39891 3628 39937 3674
rect 40007 3628 40053 3674
rect 40123 3628 40169 3674
rect 28639 3512 28685 3558
rect 28755 3512 28801 3558
rect 28871 3512 28917 3558
rect 28987 3512 29033 3558
rect 29103 3512 29149 3558
rect 29219 3512 29265 3558
rect 29335 3512 29381 3558
rect 29451 3512 29497 3558
rect 29567 3512 29613 3558
rect 29683 3512 29729 3558
rect 29799 3512 29845 3558
rect 29915 3512 29961 3558
rect 30031 3512 30077 3558
rect 30147 3512 30193 3558
rect 30263 3512 30309 3558
rect 30379 3512 30425 3558
rect 30495 3512 30541 3558
rect 30611 3512 30657 3558
rect 30727 3512 30773 3558
rect 30843 3512 30889 3558
rect 30959 3512 31005 3558
rect 31075 3512 31121 3558
rect 31191 3512 31237 3558
rect 31307 3512 31353 3558
rect 31423 3512 31469 3558
rect 31539 3512 31585 3558
rect 31655 3512 31701 3558
rect 31771 3512 31817 3558
rect 31887 3512 31933 3558
rect 32003 3512 32049 3558
rect 32119 3512 32165 3558
rect 32235 3512 32281 3558
rect 32351 3512 32397 3558
rect 32467 3512 32513 3558
rect 32583 3512 32629 3558
rect 32699 3512 32745 3558
rect 32815 3512 32861 3558
rect 32931 3512 32977 3558
rect 33047 3512 33093 3558
rect 33163 3512 33209 3558
rect 33279 3512 33325 3558
rect 33395 3512 33441 3558
rect 33511 3512 33557 3558
rect 33627 3512 33673 3558
rect 33743 3512 33789 3558
rect 33859 3512 33905 3558
rect 33975 3512 34021 3558
rect 34091 3512 34137 3558
rect 34207 3512 34253 3558
rect 34323 3512 34369 3558
rect 34439 3512 34485 3558
rect 34555 3512 34601 3558
rect 34671 3512 34717 3558
rect 34787 3512 34833 3558
rect 34903 3512 34949 3558
rect 35019 3512 35065 3558
rect 35135 3512 35181 3558
rect 35251 3512 35297 3558
rect 35367 3512 35413 3558
rect 35483 3512 35529 3558
rect 35599 3512 35645 3558
rect 35715 3512 35761 3558
rect 35831 3512 35877 3558
rect 35947 3512 35993 3558
rect 36063 3512 36109 3558
rect 36179 3512 36225 3558
rect 36295 3512 36341 3558
rect 36411 3512 36457 3558
rect 36527 3512 36573 3558
rect 36643 3512 36689 3558
rect 36759 3512 36805 3558
rect 36875 3512 36921 3558
rect 36991 3512 37037 3558
rect 37107 3512 37153 3558
rect 37223 3512 37269 3558
rect 37339 3512 37385 3558
rect 37455 3512 37501 3558
rect 37571 3512 37617 3558
rect 37687 3512 37733 3558
rect 37803 3512 37849 3558
rect 37919 3512 37965 3558
rect 38035 3512 38081 3558
rect 38151 3512 38197 3558
rect 38267 3512 38313 3558
rect 38383 3512 38429 3558
rect 38499 3512 38545 3558
rect 38615 3512 38661 3558
rect 38731 3512 38777 3558
rect 38847 3512 38893 3558
rect 38963 3512 39009 3558
rect 39079 3512 39125 3558
rect 39195 3512 39241 3558
rect 39311 3512 39357 3558
rect 39427 3512 39473 3558
rect 39543 3512 39589 3558
rect 39659 3512 39705 3558
rect 39775 3512 39821 3558
rect 39891 3512 39937 3558
rect 40007 3512 40053 3558
rect 40123 3512 40169 3558
rect 28639 3396 28685 3442
rect 28755 3396 28801 3442
rect 28871 3396 28917 3442
rect 28987 3396 29033 3442
rect 29103 3396 29149 3442
rect 29219 3396 29265 3442
rect 29335 3396 29381 3442
rect 29451 3396 29497 3442
rect 29567 3396 29613 3442
rect 29683 3396 29729 3442
rect 29799 3396 29845 3442
rect 29915 3396 29961 3442
rect 30031 3396 30077 3442
rect 30147 3396 30193 3442
rect 30263 3396 30309 3442
rect 30379 3396 30425 3442
rect 30495 3396 30541 3442
rect 30611 3396 30657 3442
rect 30727 3396 30773 3442
rect 30843 3396 30889 3442
rect 30959 3396 31005 3442
rect 31075 3396 31121 3442
rect 31191 3396 31237 3442
rect 31307 3396 31353 3442
rect 31423 3396 31469 3442
rect 31539 3396 31585 3442
rect 31655 3396 31701 3442
rect 31771 3396 31817 3442
rect 31887 3396 31933 3442
rect 32003 3396 32049 3442
rect 32119 3396 32165 3442
rect 32235 3396 32281 3442
rect 32351 3396 32397 3442
rect 32467 3396 32513 3442
rect 32583 3396 32629 3442
rect 32699 3396 32745 3442
rect 32815 3396 32861 3442
rect 32931 3396 32977 3442
rect 33047 3396 33093 3442
rect 33163 3396 33209 3442
rect 33279 3396 33325 3442
rect 33395 3396 33441 3442
rect 33511 3396 33557 3442
rect 33627 3396 33673 3442
rect 33743 3396 33789 3442
rect 33859 3396 33905 3442
rect 33975 3396 34021 3442
rect 34091 3396 34137 3442
rect 34207 3396 34253 3442
rect 34323 3396 34369 3442
rect 34439 3396 34485 3442
rect 34555 3396 34601 3442
rect 34671 3396 34717 3442
rect 34787 3396 34833 3442
rect 34903 3396 34949 3442
rect 35019 3396 35065 3442
rect 35135 3396 35181 3442
rect 35251 3396 35297 3442
rect 35367 3396 35413 3442
rect 35483 3396 35529 3442
rect 35599 3396 35645 3442
rect 35715 3396 35761 3442
rect 35831 3396 35877 3442
rect 35947 3396 35993 3442
rect 36063 3396 36109 3442
rect 36179 3396 36225 3442
rect 36295 3396 36341 3442
rect 36411 3396 36457 3442
rect 36527 3396 36573 3442
rect 36643 3396 36689 3442
rect 36759 3396 36805 3442
rect 36875 3396 36921 3442
rect 36991 3396 37037 3442
rect 37107 3396 37153 3442
rect 37223 3396 37269 3442
rect 37339 3396 37385 3442
rect 37455 3396 37501 3442
rect 37571 3396 37617 3442
rect 37687 3396 37733 3442
rect 37803 3396 37849 3442
rect 37919 3396 37965 3442
rect 38035 3396 38081 3442
rect 38151 3396 38197 3442
rect 38267 3396 38313 3442
rect 38383 3396 38429 3442
rect 38499 3396 38545 3442
rect 38615 3396 38661 3442
rect 38731 3396 38777 3442
rect 38847 3396 38893 3442
rect 38963 3396 39009 3442
rect 39079 3396 39125 3442
rect 39195 3396 39241 3442
rect 39311 3396 39357 3442
rect 39427 3396 39473 3442
rect 39543 3396 39589 3442
rect 39659 3396 39705 3442
rect 39775 3396 39821 3442
rect 39891 3396 39937 3442
rect 40007 3396 40053 3442
rect 40123 3396 40169 3442
rect 28639 3280 28685 3326
rect 28755 3280 28801 3326
rect 28871 3280 28917 3326
rect 28987 3280 29033 3326
rect 29103 3280 29149 3326
rect 29219 3280 29265 3326
rect 29335 3280 29381 3326
rect 29451 3280 29497 3326
rect 29567 3280 29613 3326
rect 29683 3280 29729 3326
rect 29799 3280 29845 3326
rect 29915 3280 29961 3326
rect 30031 3280 30077 3326
rect 30147 3280 30193 3326
rect 30263 3280 30309 3326
rect 30379 3280 30425 3326
rect 30495 3280 30541 3326
rect 30611 3280 30657 3326
rect 30727 3280 30773 3326
rect 30843 3280 30889 3326
rect 30959 3280 31005 3326
rect 31075 3280 31121 3326
rect 31191 3280 31237 3326
rect 31307 3280 31353 3326
rect 31423 3280 31469 3326
rect 31539 3280 31585 3326
rect 31655 3280 31701 3326
rect 31771 3280 31817 3326
rect 31887 3280 31933 3326
rect 32003 3280 32049 3326
rect 32119 3280 32165 3326
rect 32235 3280 32281 3326
rect 32351 3280 32397 3326
rect 32467 3280 32513 3326
rect 32583 3280 32629 3326
rect 32699 3280 32745 3326
rect 32815 3280 32861 3326
rect 32931 3280 32977 3326
rect 33047 3280 33093 3326
rect 33163 3280 33209 3326
rect 33279 3280 33325 3326
rect 33395 3280 33441 3326
rect 33511 3280 33557 3326
rect 33627 3280 33673 3326
rect 33743 3280 33789 3326
rect 33859 3280 33905 3326
rect 33975 3280 34021 3326
rect 34091 3280 34137 3326
rect 34207 3280 34253 3326
rect 34323 3280 34369 3326
rect 34439 3280 34485 3326
rect 34555 3280 34601 3326
rect 34671 3280 34717 3326
rect 34787 3280 34833 3326
rect 34903 3280 34949 3326
rect 35019 3280 35065 3326
rect 35135 3280 35181 3326
rect 35251 3280 35297 3326
rect 35367 3280 35413 3326
rect 35483 3280 35529 3326
rect 35599 3280 35645 3326
rect 35715 3280 35761 3326
rect 35831 3280 35877 3326
rect 35947 3280 35993 3326
rect 36063 3280 36109 3326
rect 36179 3280 36225 3326
rect 36295 3280 36341 3326
rect 36411 3280 36457 3326
rect 36527 3280 36573 3326
rect 36643 3280 36689 3326
rect 36759 3280 36805 3326
rect 36875 3280 36921 3326
rect 36991 3280 37037 3326
rect 37107 3280 37153 3326
rect 37223 3280 37269 3326
rect 37339 3280 37385 3326
rect 37455 3280 37501 3326
rect 37571 3280 37617 3326
rect 37687 3280 37733 3326
rect 37803 3280 37849 3326
rect 37919 3280 37965 3326
rect 38035 3280 38081 3326
rect 38151 3280 38197 3326
rect 38267 3280 38313 3326
rect 38383 3280 38429 3326
rect 38499 3280 38545 3326
rect 38615 3280 38661 3326
rect 38731 3280 38777 3326
rect 38847 3280 38893 3326
rect 38963 3280 39009 3326
rect 39079 3280 39125 3326
rect 39195 3280 39241 3326
rect 39311 3280 39357 3326
rect 39427 3280 39473 3326
rect 39543 3280 39589 3326
rect 39659 3280 39705 3326
rect 39775 3280 39821 3326
rect 39891 3280 39937 3326
rect 40007 3280 40053 3326
rect 40123 3280 40169 3326
rect 28639 3164 28685 3210
rect 28755 3164 28801 3210
rect 28871 3164 28917 3210
rect 28987 3164 29033 3210
rect 29103 3164 29149 3210
rect 29219 3164 29265 3210
rect 29335 3164 29381 3210
rect 29451 3164 29497 3210
rect 29567 3164 29613 3210
rect 29683 3164 29729 3210
rect 29799 3164 29845 3210
rect 29915 3164 29961 3210
rect 30031 3164 30077 3210
rect 30147 3164 30193 3210
rect 30263 3164 30309 3210
rect 30379 3164 30425 3210
rect 30495 3164 30541 3210
rect 30611 3164 30657 3210
rect 30727 3164 30773 3210
rect 30843 3164 30889 3210
rect 30959 3164 31005 3210
rect 31075 3164 31121 3210
rect 31191 3164 31237 3210
rect 31307 3164 31353 3210
rect 31423 3164 31469 3210
rect 31539 3164 31585 3210
rect 31655 3164 31701 3210
rect 31771 3164 31817 3210
rect 31887 3164 31933 3210
rect 32003 3164 32049 3210
rect 32119 3164 32165 3210
rect 32235 3164 32281 3210
rect 32351 3164 32397 3210
rect 32467 3164 32513 3210
rect 32583 3164 32629 3210
rect 32699 3164 32745 3210
rect 32815 3164 32861 3210
rect 32931 3164 32977 3210
rect 33047 3164 33093 3210
rect 33163 3164 33209 3210
rect 33279 3164 33325 3210
rect 33395 3164 33441 3210
rect 33511 3164 33557 3210
rect 33627 3164 33673 3210
rect 33743 3164 33789 3210
rect 33859 3164 33905 3210
rect 33975 3164 34021 3210
rect 34091 3164 34137 3210
rect 34207 3164 34253 3210
rect 34323 3164 34369 3210
rect 34439 3164 34485 3210
rect 34555 3164 34601 3210
rect 34671 3164 34717 3210
rect 34787 3164 34833 3210
rect 34903 3164 34949 3210
rect 35019 3164 35065 3210
rect 35135 3164 35181 3210
rect 35251 3164 35297 3210
rect 35367 3164 35413 3210
rect 35483 3164 35529 3210
rect 35599 3164 35645 3210
rect 35715 3164 35761 3210
rect 35831 3164 35877 3210
rect 35947 3164 35993 3210
rect 36063 3164 36109 3210
rect 36179 3164 36225 3210
rect 36295 3164 36341 3210
rect 36411 3164 36457 3210
rect 36527 3164 36573 3210
rect 36643 3164 36689 3210
rect 36759 3164 36805 3210
rect 36875 3164 36921 3210
rect 36991 3164 37037 3210
rect 37107 3164 37153 3210
rect 37223 3164 37269 3210
rect 37339 3164 37385 3210
rect 37455 3164 37501 3210
rect 37571 3164 37617 3210
rect 37687 3164 37733 3210
rect 37803 3164 37849 3210
rect 37919 3164 37965 3210
rect 38035 3164 38081 3210
rect 38151 3164 38197 3210
rect 38267 3164 38313 3210
rect 38383 3164 38429 3210
rect 38499 3164 38545 3210
rect 38615 3164 38661 3210
rect 38731 3164 38777 3210
rect 38847 3164 38893 3210
rect 38963 3164 39009 3210
rect 39079 3164 39125 3210
rect 39195 3164 39241 3210
rect 39311 3164 39357 3210
rect 39427 3164 39473 3210
rect 39543 3164 39589 3210
rect 39659 3164 39705 3210
rect 39775 3164 39821 3210
rect 39891 3164 39937 3210
rect 40007 3164 40053 3210
rect 40123 3164 40169 3210
rect 28639 3048 28685 3094
rect 28755 3048 28801 3094
rect 28871 3048 28917 3094
rect 28987 3048 29033 3094
rect 29103 3048 29149 3094
rect 29219 3048 29265 3094
rect 29335 3048 29381 3094
rect 29451 3048 29497 3094
rect 29567 3048 29613 3094
rect 29683 3048 29729 3094
rect 29799 3048 29845 3094
rect 29915 3048 29961 3094
rect 30031 3048 30077 3094
rect 30147 3048 30193 3094
rect 30263 3048 30309 3094
rect 30379 3048 30425 3094
rect 30495 3048 30541 3094
rect 30611 3048 30657 3094
rect 30727 3048 30773 3094
rect 30843 3048 30889 3094
rect 30959 3048 31005 3094
rect 31075 3048 31121 3094
rect 31191 3048 31237 3094
rect 31307 3048 31353 3094
rect 31423 3048 31469 3094
rect 31539 3048 31585 3094
rect 31655 3048 31701 3094
rect 31771 3048 31817 3094
rect 31887 3048 31933 3094
rect 32003 3048 32049 3094
rect 32119 3048 32165 3094
rect 32235 3048 32281 3094
rect 32351 3048 32397 3094
rect 32467 3048 32513 3094
rect 32583 3048 32629 3094
rect 32699 3048 32745 3094
rect 32815 3048 32861 3094
rect 32931 3048 32977 3094
rect 33047 3048 33093 3094
rect 33163 3048 33209 3094
rect 33279 3048 33325 3094
rect 33395 3048 33441 3094
rect 33511 3048 33557 3094
rect 33627 3048 33673 3094
rect 33743 3048 33789 3094
rect 33859 3048 33905 3094
rect 33975 3048 34021 3094
rect 34091 3048 34137 3094
rect 34207 3048 34253 3094
rect 34323 3048 34369 3094
rect 34439 3048 34485 3094
rect 34555 3048 34601 3094
rect 34671 3048 34717 3094
rect 34787 3048 34833 3094
rect 34903 3048 34949 3094
rect 35019 3048 35065 3094
rect 35135 3048 35181 3094
rect 35251 3048 35297 3094
rect 35367 3048 35413 3094
rect 35483 3048 35529 3094
rect 35599 3048 35645 3094
rect 35715 3048 35761 3094
rect 35831 3048 35877 3094
rect 35947 3048 35993 3094
rect 36063 3048 36109 3094
rect 36179 3048 36225 3094
rect 36295 3048 36341 3094
rect 36411 3048 36457 3094
rect 36527 3048 36573 3094
rect 36643 3048 36689 3094
rect 36759 3048 36805 3094
rect 36875 3048 36921 3094
rect 36991 3048 37037 3094
rect 37107 3048 37153 3094
rect 37223 3048 37269 3094
rect 37339 3048 37385 3094
rect 37455 3048 37501 3094
rect 37571 3048 37617 3094
rect 37687 3048 37733 3094
rect 37803 3048 37849 3094
rect 37919 3048 37965 3094
rect 38035 3048 38081 3094
rect 38151 3048 38197 3094
rect 38267 3048 38313 3094
rect 38383 3048 38429 3094
rect 38499 3048 38545 3094
rect 38615 3048 38661 3094
rect 38731 3048 38777 3094
rect 38847 3048 38893 3094
rect 38963 3048 39009 3094
rect 39079 3048 39125 3094
rect 39195 3048 39241 3094
rect 39311 3048 39357 3094
rect 39427 3048 39473 3094
rect 39543 3048 39589 3094
rect 39659 3048 39705 3094
rect 39775 3048 39821 3094
rect 39891 3048 39937 3094
rect 40007 3048 40053 3094
rect 40123 3048 40169 3094
rect 28639 2932 28685 2978
rect 28755 2932 28801 2978
rect 28871 2932 28917 2978
rect 28987 2932 29033 2978
rect 29103 2932 29149 2978
rect 29219 2932 29265 2978
rect 29335 2932 29381 2978
rect 29451 2932 29497 2978
rect 29567 2932 29613 2978
rect 29683 2932 29729 2978
rect 29799 2932 29845 2978
rect 29915 2932 29961 2978
rect 30031 2932 30077 2978
rect 30147 2932 30193 2978
rect 30263 2932 30309 2978
rect 30379 2932 30425 2978
rect 30495 2932 30541 2978
rect 30611 2932 30657 2978
rect 30727 2932 30773 2978
rect 30843 2932 30889 2978
rect 30959 2932 31005 2978
rect 31075 2932 31121 2978
rect 31191 2932 31237 2978
rect 31307 2932 31353 2978
rect 31423 2932 31469 2978
rect 31539 2932 31585 2978
rect 31655 2932 31701 2978
rect 31771 2932 31817 2978
rect 31887 2932 31933 2978
rect 32003 2932 32049 2978
rect 32119 2932 32165 2978
rect 32235 2932 32281 2978
rect 32351 2932 32397 2978
rect 32467 2932 32513 2978
rect 32583 2932 32629 2978
rect 32699 2932 32745 2978
rect 32815 2932 32861 2978
rect 32931 2932 32977 2978
rect 33047 2932 33093 2978
rect 33163 2932 33209 2978
rect 33279 2932 33325 2978
rect 33395 2932 33441 2978
rect 33511 2932 33557 2978
rect 33627 2932 33673 2978
rect 33743 2932 33789 2978
rect 33859 2932 33905 2978
rect 33975 2932 34021 2978
rect 34091 2932 34137 2978
rect 34207 2932 34253 2978
rect 34323 2932 34369 2978
rect 34439 2932 34485 2978
rect 34555 2932 34601 2978
rect 34671 2932 34717 2978
rect 34787 2932 34833 2978
rect 34903 2932 34949 2978
rect 35019 2932 35065 2978
rect 35135 2932 35181 2978
rect 35251 2932 35297 2978
rect 35367 2932 35413 2978
rect 35483 2932 35529 2978
rect 35599 2932 35645 2978
rect 35715 2932 35761 2978
rect 35831 2932 35877 2978
rect 35947 2932 35993 2978
rect 36063 2932 36109 2978
rect 36179 2932 36225 2978
rect 36295 2932 36341 2978
rect 36411 2932 36457 2978
rect 36527 2932 36573 2978
rect 36643 2932 36689 2978
rect 36759 2932 36805 2978
rect 36875 2932 36921 2978
rect 36991 2932 37037 2978
rect 37107 2932 37153 2978
rect 37223 2932 37269 2978
rect 37339 2932 37385 2978
rect 37455 2932 37501 2978
rect 37571 2932 37617 2978
rect 37687 2932 37733 2978
rect 37803 2932 37849 2978
rect 37919 2932 37965 2978
rect 38035 2932 38081 2978
rect 38151 2932 38197 2978
rect 38267 2932 38313 2978
rect 38383 2932 38429 2978
rect 38499 2932 38545 2978
rect 38615 2932 38661 2978
rect 38731 2932 38777 2978
rect 38847 2932 38893 2978
rect 38963 2932 39009 2978
rect 39079 2932 39125 2978
rect 39195 2932 39241 2978
rect 39311 2932 39357 2978
rect 39427 2932 39473 2978
rect 39543 2932 39589 2978
rect 39659 2932 39705 2978
rect 39775 2932 39821 2978
rect 39891 2932 39937 2978
rect 40007 2932 40053 2978
rect 40123 2932 40169 2978
rect 28639 2816 28685 2862
rect 28755 2816 28801 2862
rect 28871 2816 28917 2862
rect 28987 2816 29033 2862
rect 29103 2816 29149 2862
rect 29219 2816 29265 2862
rect 29335 2816 29381 2862
rect 29451 2816 29497 2862
rect 29567 2816 29613 2862
rect 29683 2816 29729 2862
rect 29799 2816 29845 2862
rect 29915 2816 29961 2862
rect 30031 2816 30077 2862
rect 30147 2816 30193 2862
rect 30263 2816 30309 2862
rect 30379 2816 30425 2862
rect 30495 2816 30541 2862
rect 30611 2816 30657 2862
rect 30727 2816 30773 2862
rect 30843 2816 30889 2862
rect 30959 2816 31005 2862
rect 31075 2816 31121 2862
rect 31191 2816 31237 2862
rect 31307 2816 31353 2862
rect 31423 2816 31469 2862
rect 31539 2816 31585 2862
rect 31655 2816 31701 2862
rect 31771 2816 31817 2862
rect 31887 2816 31933 2862
rect 32003 2816 32049 2862
rect 32119 2816 32165 2862
rect 32235 2816 32281 2862
rect 32351 2816 32397 2862
rect 32467 2816 32513 2862
rect 32583 2816 32629 2862
rect 32699 2816 32745 2862
rect 32815 2816 32861 2862
rect 32931 2816 32977 2862
rect 33047 2816 33093 2862
rect 33163 2816 33209 2862
rect 33279 2816 33325 2862
rect 33395 2816 33441 2862
rect 33511 2816 33557 2862
rect 33627 2816 33673 2862
rect 33743 2816 33789 2862
rect 33859 2816 33905 2862
rect 33975 2816 34021 2862
rect 34091 2816 34137 2862
rect 34207 2816 34253 2862
rect 34323 2816 34369 2862
rect 34439 2816 34485 2862
rect 34555 2816 34601 2862
rect 34671 2816 34717 2862
rect 34787 2816 34833 2862
rect 34903 2816 34949 2862
rect 35019 2816 35065 2862
rect 35135 2816 35181 2862
rect 35251 2816 35297 2862
rect 35367 2816 35413 2862
rect 35483 2816 35529 2862
rect 35599 2816 35645 2862
rect 35715 2816 35761 2862
rect 35831 2816 35877 2862
rect 35947 2816 35993 2862
rect 36063 2816 36109 2862
rect 36179 2816 36225 2862
rect 36295 2816 36341 2862
rect 36411 2816 36457 2862
rect 36527 2816 36573 2862
rect 36643 2816 36689 2862
rect 36759 2816 36805 2862
rect 36875 2816 36921 2862
rect 36991 2816 37037 2862
rect 37107 2816 37153 2862
rect 37223 2816 37269 2862
rect 37339 2816 37385 2862
rect 37455 2816 37501 2862
rect 37571 2816 37617 2862
rect 37687 2816 37733 2862
rect 37803 2816 37849 2862
rect 37919 2816 37965 2862
rect 38035 2816 38081 2862
rect 38151 2816 38197 2862
rect 38267 2816 38313 2862
rect 38383 2816 38429 2862
rect 38499 2816 38545 2862
rect 38615 2816 38661 2862
rect 38731 2816 38777 2862
rect 38847 2816 38893 2862
rect 38963 2816 39009 2862
rect 39079 2816 39125 2862
rect 39195 2816 39241 2862
rect 39311 2816 39357 2862
rect 39427 2816 39473 2862
rect 39543 2816 39589 2862
rect 39659 2816 39705 2862
rect 39775 2816 39821 2862
rect 39891 2816 39937 2862
rect 40007 2816 40053 2862
rect 40123 2816 40169 2862
rect 28639 2700 28685 2746
rect 28755 2700 28801 2746
rect 28871 2700 28917 2746
rect 28987 2700 29033 2746
rect 29103 2700 29149 2746
rect 29219 2700 29265 2746
rect 29335 2700 29381 2746
rect 29451 2700 29497 2746
rect 29567 2700 29613 2746
rect 29683 2700 29729 2746
rect 29799 2700 29845 2746
rect 29915 2700 29961 2746
rect 30031 2700 30077 2746
rect 30147 2700 30193 2746
rect 30263 2700 30309 2746
rect 30379 2700 30425 2746
rect 30495 2700 30541 2746
rect 30611 2700 30657 2746
rect 30727 2700 30773 2746
rect 30843 2700 30889 2746
rect 30959 2700 31005 2746
rect 31075 2700 31121 2746
rect 31191 2700 31237 2746
rect 31307 2700 31353 2746
rect 31423 2700 31469 2746
rect 31539 2700 31585 2746
rect 31655 2700 31701 2746
rect 31771 2700 31817 2746
rect 31887 2700 31933 2746
rect 32003 2700 32049 2746
rect 32119 2700 32165 2746
rect 32235 2700 32281 2746
rect 32351 2700 32397 2746
rect 32467 2700 32513 2746
rect 32583 2700 32629 2746
rect 32699 2700 32745 2746
rect 32815 2700 32861 2746
rect 32931 2700 32977 2746
rect 33047 2700 33093 2746
rect 33163 2700 33209 2746
rect 33279 2700 33325 2746
rect 33395 2700 33441 2746
rect 33511 2700 33557 2746
rect 33627 2700 33673 2746
rect 33743 2700 33789 2746
rect 33859 2700 33905 2746
rect 33975 2700 34021 2746
rect 34091 2700 34137 2746
rect 34207 2700 34253 2746
rect 34323 2700 34369 2746
rect 34439 2700 34485 2746
rect 34555 2700 34601 2746
rect 34671 2700 34717 2746
rect 34787 2700 34833 2746
rect 34903 2700 34949 2746
rect 35019 2700 35065 2746
rect 35135 2700 35181 2746
rect 35251 2700 35297 2746
rect 35367 2700 35413 2746
rect 35483 2700 35529 2746
rect 35599 2700 35645 2746
rect 35715 2700 35761 2746
rect 35831 2700 35877 2746
rect 35947 2700 35993 2746
rect 36063 2700 36109 2746
rect 36179 2700 36225 2746
rect 36295 2700 36341 2746
rect 36411 2700 36457 2746
rect 36527 2700 36573 2746
rect 36643 2700 36689 2746
rect 36759 2700 36805 2746
rect 36875 2700 36921 2746
rect 36991 2700 37037 2746
rect 37107 2700 37153 2746
rect 37223 2700 37269 2746
rect 37339 2700 37385 2746
rect 37455 2700 37501 2746
rect 37571 2700 37617 2746
rect 37687 2700 37733 2746
rect 37803 2700 37849 2746
rect 37919 2700 37965 2746
rect 38035 2700 38081 2746
rect 38151 2700 38197 2746
rect 38267 2700 38313 2746
rect 38383 2700 38429 2746
rect 38499 2700 38545 2746
rect 38615 2700 38661 2746
rect 38731 2700 38777 2746
rect 38847 2700 38893 2746
rect 38963 2700 39009 2746
rect 39079 2700 39125 2746
rect 39195 2700 39241 2746
rect 39311 2700 39357 2746
rect 39427 2700 39473 2746
rect 39543 2700 39589 2746
rect 39659 2700 39705 2746
rect 39775 2700 39821 2746
rect 39891 2700 39937 2746
rect 40007 2700 40053 2746
rect 40123 2700 40169 2746
rect 28639 2584 28685 2630
rect 28755 2584 28801 2630
rect 28871 2584 28917 2630
rect 28987 2584 29033 2630
rect 29103 2584 29149 2630
rect 29219 2584 29265 2630
rect 29335 2584 29381 2630
rect 29451 2584 29497 2630
rect 29567 2584 29613 2630
rect 29683 2584 29729 2630
rect 29799 2584 29845 2630
rect 29915 2584 29961 2630
rect 30031 2584 30077 2630
rect 30147 2584 30193 2630
rect 30263 2584 30309 2630
rect 30379 2584 30425 2630
rect 30495 2584 30541 2630
rect 30611 2584 30657 2630
rect 30727 2584 30773 2630
rect 30843 2584 30889 2630
rect 30959 2584 31005 2630
rect 31075 2584 31121 2630
rect 31191 2584 31237 2630
rect 31307 2584 31353 2630
rect 31423 2584 31469 2630
rect 31539 2584 31585 2630
rect 31655 2584 31701 2630
rect 31771 2584 31817 2630
rect 31887 2584 31933 2630
rect 32003 2584 32049 2630
rect 32119 2584 32165 2630
rect 32235 2584 32281 2630
rect 32351 2584 32397 2630
rect 32467 2584 32513 2630
rect 32583 2584 32629 2630
rect 32699 2584 32745 2630
rect 32815 2584 32861 2630
rect 32931 2584 32977 2630
rect 33047 2584 33093 2630
rect 33163 2584 33209 2630
rect 33279 2584 33325 2630
rect 33395 2584 33441 2630
rect 33511 2584 33557 2630
rect 33627 2584 33673 2630
rect 33743 2584 33789 2630
rect 33859 2584 33905 2630
rect 33975 2584 34021 2630
rect 34091 2584 34137 2630
rect 34207 2584 34253 2630
rect 34323 2584 34369 2630
rect 34439 2584 34485 2630
rect 34555 2584 34601 2630
rect 34671 2584 34717 2630
rect 34787 2584 34833 2630
rect 34903 2584 34949 2630
rect 35019 2584 35065 2630
rect 35135 2584 35181 2630
rect 35251 2584 35297 2630
rect 35367 2584 35413 2630
rect 35483 2584 35529 2630
rect 35599 2584 35645 2630
rect 35715 2584 35761 2630
rect 35831 2584 35877 2630
rect 35947 2584 35993 2630
rect 36063 2584 36109 2630
rect 36179 2584 36225 2630
rect 36295 2584 36341 2630
rect 36411 2584 36457 2630
rect 36527 2584 36573 2630
rect 36643 2584 36689 2630
rect 36759 2584 36805 2630
rect 36875 2584 36921 2630
rect 36991 2584 37037 2630
rect 37107 2584 37153 2630
rect 37223 2584 37269 2630
rect 37339 2584 37385 2630
rect 37455 2584 37501 2630
rect 37571 2584 37617 2630
rect 37687 2584 37733 2630
rect 37803 2584 37849 2630
rect 37919 2584 37965 2630
rect 38035 2584 38081 2630
rect 38151 2584 38197 2630
rect 38267 2584 38313 2630
rect 38383 2584 38429 2630
rect 38499 2584 38545 2630
rect 38615 2584 38661 2630
rect 38731 2584 38777 2630
rect 38847 2584 38893 2630
rect 38963 2584 39009 2630
rect 39079 2584 39125 2630
rect 39195 2584 39241 2630
rect 39311 2584 39357 2630
rect 39427 2584 39473 2630
rect 39543 2584 39589 2630
rect 39659 2584 39705 2630
rect 39775 2584 39821 2630
rect 39891 2584 39937 2630
rect 40007 2584 40053 2630
rect 40123 2584 40169 2630
rect 28639 2468 28685 2514
rect 28755 2468 28801 2514
rect 28871 2468 28917 2514
rect 28987 2468 29033 2514
rect 29103 2468 29149 2514
rect 29219 2468 29265 2514
rect 29335 2468 29381 2514
rect 29451 2468 29497 2514
rect 29567 2468 29613 2514
rect 29683 2468 29729 2514
rect 29799 2468 29845 2514
rect 29915 2468 29961 2514
rect 30031 2468 30077 2514
rect 30147 2468 30193 2514
rect 30263 2468 30309 2514
rect 30379 2468 30425 2514
rect 30495 2468 30541 2514
rect 30611 2468 30657 2514
rect 30727 2468 30773 2514
rect 30843 2468 30889 2514
rect 30959 2468 31005 2514
rect 31075 2468 31121 2514
rect 31191 2468 31237 2514
rect 31307 2468 31353 2514
rect 31423 2468 31469 2514
rect 31539 2468 31585 2514
rect 31655 2468 31701 2514
rect 31771 2468 31817 2514
rect 31887 2468 31933 2514
rect 32003 2468 32049 2514
rect 32119 2468 32165 2514
rect 32235 2468 32281 2514
rect 32351 2468 32397 2514
rect 32467 2468 32513 2514
rect 32583 2468 32629 2514
rect 32699 2468 32745 2514
rect 32815 2468 32861 2514
rect 32931 2468 32977 2514
rect 33047 2468 33093 2514
rect 33163 2468 33209 2514
rect 33279 2468 33325 2514
rect 33395 2468 33441 2514
rect 33511 2468 33557 2514
rect 33627 2468 33673 2514
rect 33743 2468 33789 2514
rect 33859 2468 33905 2514
rect 33975 2468 34021 2514
rect 34091 2468 34137 2514
rect 34207 2468 34253 2514
rect 34323 2468 34369 2514
rect 34439 2468 34485 2514
rect 34555 2468 34601 2514
rect 34671 2468 34717 2514
rect 34787 2468 34833 2514
rect 34903 2468 34949 2514
rect 35019 2468 35065 2514
rect 35135 2468 35181 2514
rect 35251 2468 35297 2514
rect 35367 2468 35413 2514
rect 35483 2468 35529 2514
rect 35599 2468 35645 2514
rect 35715 2468 35761 2514
rect 35831 2468 35877 2514
rect 35947 2468 35993 2514
rect 36063 2468 36109 2514
rect 36179 2468 36225 2514
rect 36295 2468 36341 2514
rect 36411 2468 36457 2514
rect 36527 2468 36573 2514
rect 36643 2468 36689 2514
rect 36759 2468 36805 2514
rect 36875 2468 36921 2514
rect 36991 2468 37037 2514
rect 37107 2468 37153 2514
rect 37223 2468 37269 2514
rect 37339 2468 37385 2514
rect 37455 2468 37501 2514
rect 37571 2468 37617 2514
rect 37687 2468 37733 2514
rect 37803 2468 37849 2514
rect 37919 2468 37965 2514
rect 38035 2468 38081 2514
rect 38151 2468 38197 2514
rect 38267 2468 38313 2514
rect 38383 2468 38429 2514
rect 38499 2468 38545 2514
rect 38615 2468 38661 2514
rect 38731 2468 38777 2514
rect 38847 2468 38893 2514
rect 38963 2468 39009 2514
rect 39079 2468 39125 2514
rect 39195 2468 39241 2514
rect 39311 2468 39357 2514
rect 39427 2468 39473 2514
rect 39543 2468 39589 2514
rect 39659 2468 39705 2514
rect 39775 2468 39821 2514
rect 39891 2468 39937 2514
rect 40007 2468 40053 2514
rect 40123 2468 40169 2514
rect 28639 2352 28685 2398
rect 28755 2352 28801 2398
rect 28871 2352 28917 2398
rect 28987 2352 29033 2398
rect 29103 2352 29149 2398
rect 29219 2352 29265 2398
rect 29335 2352 29381 2398
rect 29451 2352 29497 2398
rect 29567 2352 29613 2398
rect 29683 2352 29729 2398
rect 29799 2352 29845 2398
rect 29915 2352 29961 2398
rect 30031 2352 30077 2398
rect 30147 2352 30193 2398
rect 30263 2352 30309 2398
rect 30379 2352 30425 2398
rect 30495 2352 30541 2398
rect 30611 2352 30657 2398
rect 30727 2352 30773 2398
rect 30843 2352 30889 2398
rect 30959 2352 31005 2398
rect 31075 2352 31121 2398
rect 31191 2352 31237 2398
rect 31307 2352 31353 2398
rect 31423 2352 31469 2398
rect 31539 2352 31585 2398
rect 31655 2352 31701 2398
rect 31771 2352 31817 2398
rect 31887 2352 31933 2398
rect 32003 2352 32049 2398
rect 32119 2352 32165 2398
rect 32235 2352 32281 2398
rect 32351 2352 32397 2398
rect 32467 2352 32513 2398
rect 32583 2352 32629 2398
rect 32699 2352 32745 2398
rect 32815 2352 32861 2398
rect 32931 2352 32977 2398
rect 33047 2352 33093 2398
rect 33163 2352 33209 2398
rect 33279 2352 33325 2398
rect 33395 2352 33441 2398
rect 33511 2352 33557 2398
rect 33627 2352 33673 2398
rect 33743 2352 33789 2398
rect 33859 2352 33905 2398
rect 33975 2352 34021 2398
rect 34091 2352 34137 2398
rect 34207 2352 34253 2398
rect 34323 2352 34369 2398
rect 34439 2352 34485 2398
rect 34555 2352 34601 2398
rect 34671 2352 34717 2398
rect 34787 2352 34833 2398
rect 34903 2352 34949 2398
rect 35019 2352 35065 2398
rect 35135 2352 35181 2398
rect 35251 2352 35297 2398
rect 35367 2352 35413 2398
rect 35483 2352 35529 2398
rect 35599 2352 35645 2398
rect 35715 2352 35761 2398
rect 35831 2352 35877 2398
rect 35947 2352 35993 2398
rect 36063 2352 36109 2398
rect 36179 2352 36225 2398
rect 36295 2352 36341 2398
rect 36411 2352 36457 2398
rect 36527 2352 36573 2398
rect 36643 2352 36689 2398
rect 36759 2352 36805 2398
rect 36875 2352 36921 2398
rect 36991 2352 37037 2398
rect 37107 2352 37153 2398
rect 37223 2352 37269 2398
rect 37339 2352 37385 2398
rect 37455 2352 37501 2398
rect 37571 2352 37617 2398
rect 37687 2352 37733 2398
rect 37803 2352 37849 2398
rect 37919 2352 37965 2398
rect 38035 2352 38081 2398
rect 38151 2352 38197 2398
rect 38267 2352 38313 2398
rect 38383 2352 38429 2398
rect 38499 2352 38545 2398
rect 38615 2352 38661 2398
rect 38731 2352 38777 2398
rect 38847 2352 38893 2398
rect 38963 2352 39009 2398
rect 39079 2352 39125 2398
rect 39195 2352 39241 2398
rect 39311 2352 39357 2398
rect 39427 2352 39473 2398
rect 39543 2352 39589 2398
rect 39659 2352 39705 2398
rect 39775 2352 39821 2398
rect 39891 2352 39937 2398
rect 40007 2352 40053 2398
rect 40123 2352 40169 2398
rect 28639 2236 28685 2282
rect 28755 2236 28801 2282
rect 28871 2236 28917 2282
rect 28987 2236 29033 2282
rect 29103 2236 29149 2282
rect 29219 2236 29265 2282
rect 29335 2236 29381 2282
rect 29451 2236 29497 2282
rect 29567 2236 29613 2282
rect 29683 2236 29729 2282
rect 29799 2236 29845 2282
rect 29915 2236 29961 2282
rect 30031 2236 30077 2282
rect 30147 2236 30193 2282
rect 30263 2236 30309 2282
rect 30379 2236 30425 2282
rect 30495 2236 30541 2282
rect 30611 2236 30657 2282
rect 30727 2236 30773 2282
rect 30843 2236 30889 2282
rect 30959 2236 31005 2282
rect 31075 2236 31121 2282
rect 31191 2236 31237 2282
rect 31307 2236 31353 2282
rect 31423 2236 31469 2282
rect 31539 2236 31585 2282
rect 31655 2236 31701 2282
rect 31771 2236 31817 2282
rect 31887 2236 31933 2282
rect 32003 2236 32049 2282
rect 32119 2236 32165 2282
rect 32235 2236 32281 2282
rect 32351 2236 32397 2282
rect 32467 2236 32513 2282
rect 32583 2236 32629 2282
rect 32699 2236 32745 2282
rect 32815 2236 32861 2282
rect 32931 2236 32977 2282
rect 33047 2236 33093 2282
rect 33163 2236 33209 2282
rect 33279 2236 33325 2282
rect 33395 2236 33441 2282
rect 33511 2236 33557 2282
rect 33627 2236 33673 2282
rect 33743 2236 33789 2282
rect 33859 2236 33905 2282
rect 33975 2236 34021 2282
rect 34091 2236 34137 2282
rect 34207 2236 34253 2282
rect 34323 2236 34369 2282
rect 34439 2236 34485 2282
rect 34555 2236 34601 2282
rect 34671 2236 34717 2282
rect 34787 2236 34833 2282
rect 34903 2236 34949 2282
rect 35019 2236 35065 2282
rect 35135 2236 35181 2282
rect 35251 2236 35297 2282
rect 35367 2236 35413 2282
rect 35483 2236 35529 2282
rect 35599 2236 35645 2282
rect 35715 2236 35761 2282
rect 35831 2236 35877 2282
rect 35947 2236 35993 2282
rect 36063 2236 36109 2282
rect 36179 2236 36225 2282
rect 36295 2236 36341 2282
rect 36411 2236 36457 2282
rect 36527 2236 36573 2282
rect 36643 2236 36689 2282
rect 36759 2236 36805 2282
rect 36875 2236 36921 2282
rect 36991 2236 37037 2282
rect 37107 2236 37153 2282
rect 37223 2236 37269 2282
rect 37339 2236 37385 2282
rect 37455 2236 37501 2282
rect 37571 2236 37617 2282
rect 37687 2236 37733 2282
rect 37803 2236 37849 2282
rect 37919 2236 37965 2282
rect 38035 2236 38081 2282
rect 38151 2236 38197 2282
rect 38267 2236 38313 2282
rect 38383 2236 38429 2282
rect 38499 2236 38545 2282
rect 38615 2236 38661 2282
rect 38731 2236 38777 2282
rect 38847 2236 38893 2282
rect 38963 2236 39009 2282
rect 39079 2236 39125 2282
rect 39195 2236 39241 2282
rect 39311 2236 39357 2282
rect 39427 2236 39473 2282
rect 39543 2236 39589 2282
rect 39659 2236 39705 2282
rect 39775 2236 39821 2282
rect 39891 2236 39937 2282
rect 40007 2236 40053 2282
rect 40123 2236 40169 2282
rect 28639 2120 28685 2166
rect 28755 2120 28801 2166
rect 28871 2120 28917 2166
rect 28987 2120 29033 2166
rect 29103 2120 29149 2166
rect 29219 2120 29265 2166
rect 29335 2120 29381 2166
rect 29451 2120 29497 2166
rect 29567 2120 29613 2166
rect 29683 2120 29729 2166
rect 29799 2120 29845 2166
rect 29915 2120 29961 2166
rect 30031 2120 30077 2166
rect 30147 2120 30193 2166
rect 30263 2120 30309 2166
rect 30379 2120 30425 2166
rect 30495 2120 30541 2166
rect 30611 2120 30657 2166
rect 30727 2120 30773 2166
rect 30843 2120 30889 2166
rect 30959 2120 31005 2166
rect 31075 2120 31121 2166
rect 31191 2120 31237 2166
rect 31307 2120 31353 2166
rect 31423 2120 31469 2166
rect 31539 2120 31585 2166
rect 31655 2120 31701 2166
rect 31771 2120 31817 2166
rect 31887 2120 31933 2166
rect 32003 2120 32049 2166
rect 32119 2120 32165 2166
rect 32235 2120 32281 2166
rect 32351 2120 32397 2166
rect 32467 2120 32513 2166
rect 32583 2120 32629 2166
rect 32699 2120 32745 2166
rect 32815 2120 32861 2166
rect 32931 2120 32977 2166
rect 33047 2120 33093 2166
rect 33163 2120 33209 2166
rect 33279 2120 33325 2166
rect 33395 2120 33441 2166
rect 33511 2120 33557 2166
rect 33627 2120 33673 2166
rect 33743 2120 33789 2166
rect 33859 2120 33905 2166
rect 33975 2120 34021 2166
rect 34091 2120 34137 2166
rect 34207 2120 34253 2166
rect 34323 2120 34369 2166
rect 34439 2120 34485 2166
rect 34555 2120 34601 2166
rect 34671 2120 34717 2166
rect 34787 2120 34833 2166
rect 34903 2120 34949 2166
rect 35019 2120 35065 2166
rect 35135 2120 35181 2166
rect 35251 2120 35297 2166
rect 35367 2120 35413 2166
rect 35483 2120 35529 2166
rect 35599 2120 35645 2166
rect 35715 2120 35761 2166
rect 35831 2120 35877 2166
rect 35947 2120 35993 2166
rect 36063 2120 36109 2166
rect 36179 2120 36225 2166
rect 36295 2120 36341 2166
rect 36411 2120 36457 2166
rect 36527 2120 36573 2166
rect 36643 2120 36689 2166
rect 36759 2120 36805 2166
rect 36875 2120 36921 2166
rect 36991 2120 37037 2166
rect 37107 2120 37153 2166
rect 37223 2120 37269 2166
rect 37339 2120 37385 2166
rect 37455 2120 37501 2166
rect 37571 2120 37617 2166
rect 37687 2120 37733 2166
rect 37803 2120 37849 2166
rect 37919 2120 37965 2166
rect 38035 2120 38081 2166
rect 38151 2120 38197 2166
rect 38267 2120 38313 2166
rect 38383 2120 38429 2166
rect 38499 2120 38545 2166
rect 38615 2120 38661 2166
rect 38731 2120 38777 2166
rect 38847 2120 38893 2166
rect 38963 2120 39009 2166
rect 39079 2120 39125 2166
rect 39195 2120 39241 2166
rect 39311 2120 39357 2166
rect 39427 2120 39473 2166
rect 39543 2120 39589 2166
rect 39659 2120 39705 2166
rect 39775 2120 39821 2166
rect 39891 2120 39937 2166
rect 40007 2120 40053 2166
rect 40123 2120 40169 2166
rect 28639 2004 28685 2050
rect 28755 2004 28801 2050
rect 28871 2004 28917 2050
rect 28987 2004 29033 2050
rect 29103 2004 29149 2050
rect 29219 2004 29265 2050
rect 29335 2004 29381 2050
rect 29451 2004 29497 2050
rect 29567 2004 29613 2050
rect 29683 2004 29729 2050
rect 29799 2004 29845 2050
rect 29915 2004 29961 2050
rect 30031 2004 30077 2050
rect 30147 2004 30193 2050
rect 30263 2004 30309 2050
rect 30379 2004 30425 2050
rect 30495 2004 30541 2050
rect 30611 2004 30657 2050
rect 30727 2004 30773 2050
rect 30843 2004 30889 2050
rect 30959 2004 31005 2050
rect 31075 2004 31121 2050
rect 31191 2004 31237 2050
rect 31307 2004 31353 2050
rect 31423 2004 31469 2050
rect 31539 2004 31585 2050
rect 31655 2004 31701 2050
rect 31771 2004 31817 2050
rect 31887 2004 31933 2050
rect 32003 2004 32049 2050
rect 32119 2004 32165 2050
rect 32235 2004 32281 2050
rect 32351 2004 32397 2050
rect 32467 2004 32513 2050
rect 32583 2004 32629 2050
rect 32699 2004 32745 2050
rect 32815 2004 32861 2050
rect 32931 2004 32977 2050
rect 33047 2004 33093 2050
rect 33163 2004 33209 2050
rect 33279 2004 33325 2050
rect 33395 2004 33441 2050
rect 33511 2004 33557 2050
rect 33627 2004 33673 2050
rect 33743 2004 33789 2050
rect 33859 2004 33905 2050
rect 33975 2004 34021 2050
rect 34091 2004 34137 2050
rect 34207 2004 34253 2050
rect 34323 2004 34369 2050
rect 34439 2004 34485 2050
rect 34555 2004 34601 2050
rect 34671 2004 34717 2050
rect 34787 2004 34833 2050
rect 34903 2004 34949 2050
rect 35019 2004 35065 2050
rect 35135 2004 35181 2050
rect 35251 2004 35297 2050
rect 35367 2004 35413 2050
rect 35483 2004 35529 2050
rect 35599 2004 35645 2050
rect 35715 2004 35761 2050
rect 35831 2004 35877 2050
rect 35947 2004 35993 2050
rect 36063 2004 36109 2050
rect 36179 2004 36225 2050
rect 36295 2004 36341 2050
rect 36411 2004 36457 2050
rect 36527 2004 36573 2050
rect 36643 2004 36689 2050
rect 36759 2004 36805 2050
rect 36875 2004 36921 2050
rect 36991 2004 37037 2050
rect 37107 2004 37153 2050
rect 37223 2004 37269 2050
rect 37339 2004 37385 2050
rect 37455 2004 37501 2050
rect 37571 2004 37617 2050
rect 37687 2004 37733 2050
rect 37803 2004 37849 2050
rect 37919 2004 37965 2050
rect 38035 2004 38081 2050
rect 38151 2004 38197 2050
rect 38267 2004 38313 2050
rect 38383 2004 38429 2050
rect 38499 2004 38545 2050
rect 38615 2004 38661 2050
rect 38731 2004 38777 2050
rect 38847 2004 38893 2050
rect 38963 2004 39009 2050
rect 39079 2004 39125 2050
rect 39195 2004 39241 2050
rect 39311 2004 39357 2050
rect 39427 2004 39473 2050
rect 39543 2004 39589 2050
rect 39659 2004 39705 2050
rect 39775 2004 39821 2050
rect 39891 2004 39937 2050
rect 40007 2004 40053 2050
rect 40123 2004 40169 2050
rect 28639 1888 28685 1934
rect 28755 1888 28801 1934
rect 28871 1888 28917 1934
rect 28987 1888 29033 1934
rect 29103 1888 29149 1934
rect 29219 1888 29265 1934
rect 29335 1888 29381 1934
rect 29451 1888 29497 1934
rect 29567 1888 29613 1934
rect 29683 1888 29729 1934
rect 29799 1888 29845 1934
rect 29915 1888 29961 1934
rect 30031 1888 30077 1934
rect 30147 1888 30193 1934
rect 30263 1888 30309 1934
rect 30379 1888 30425 1934
rect 30495 1888 30541 1934
rect 30611 1888 30657 1934
rect 30727 1888 30773 1934
rect 30843 1888 30889 1934
rect 30959 1888 31005 1934
rect 31075 1888 31121 1934
rect 31191 1888 31237 1934
rect 31307 1888 31353 1934
rect 31423 1888 31469 1934
rect 31539 1888 31585 1934
rect 31655 1888 31701 1934
rect 31771 1888 31817 1934
rect 31887 1888 31933 1934
rect 32003 1888 32049 1934
rect 32119 1888 32165 1934
rect 32235 1888 32281 1934
rect 32351 1888 32397 1934
rect 32467 1888 32513 1934
rect 32583 1888 32629 1934
rect 32699 1888 32745 1934
rect 32815 1888 32861 1934
rect 32931 1888 32977 1934
rect 33047 1888 33093 1934
rect 33163 1888 33209 1934
rect 33279 1888 33325 1934
rect 33395 1888 33441 1934
rect 33511 1888 33557 1934
rect 33627 1888 33673 1934
rect 33743 1888 33789 1934
rect 33859 1888 33905 1934
rect 33975 1888 34021 1934
rect 34091 1888 34137 1934
rect 34207 1888 34253 1934
rect 34323 1888 34369 1934
rect 34439 1888 34485 1934
rect 34555 1888 34601 1934
rect 34671 1888 34717 1934
rect 34787 1888 34833 1934
rect 34903 1888 34949 1934
rect 35019 1888 35065 1934
rect 35135 1888 35181 1934
rect 35251 1888 35297 1934
rect 35367 1888 35413 1934
rect 35483 1888 35529 1934
rect 35599 1888 35645 1934
rect 35715 1888 35761 1934
rect 35831 1888 35877 1934
rect 35947 1888 35993 1934
rect 36063 1888 36109 1934
rect 36179 1888 36225 1934
rect 36295 1888 36341 1934
rect 36411 1888 36457 1934
rect 36527 1888 36573 1934
rect 36643 1888 36689 1934
rect 36759 1888 36805 1934
rect 36875 1888 36921 1934
rect 36991 1888 37037 1934
rect 37107 1888 37153 1934
rect 37223 1888 37269 1934
rect 37339 1888 37385 1934
rect 37455 1888 37501 1934
rect 37571 1888 37617 1934
rect 37687 1888 37733 1934
rect 37803 1888 37849 1934
rect 37919 1888 37965 1934
rect 38035 1888 38081 1934
rect 38151 1888 38197 1934
rect 38267 1888 38313 1934
rect 38383 1888 38429 1934
rect 38499 1888 38545 1934
rect 38615 1888 38661 1934
rect 38731 1888 38777 1934
rect 38847 1888 38893 1934
rect 38963 1888 39009 1934
rect 39079 1888 39125 1934
rect 39195 1888 39241 1934
rect 39311 1888 39357 1934
rect 39427 1888 39473 1934
rect 39543 1888 39589 1934
rect 39659 1888 39705 1934
rect 39775 1888 39821 1934
rect 39891 1888 39937 1934
rect 40007 1888 40053 1934
rect 40123 1888 40169 1934
rect 28639 1772 28685 1818
rect 28755 1772 28801 1818
rect 28871 1772 28917 1818
rect 28987 1772 29033 1818
rect 29103 1772 29149 1818
rect 29219 1772 29265 1818
rect 29335 1772 29381 1818
rect 29451 1772 29497 1818
rect 29567 1772 29613 1818
rect 29683 1772 29729 1818
rect 29799 1772 29845 1818
rect 29915 1772 29961 1818
rect 30031 1772 30077 1818
rect 30147 1772 30193 1818
rect 30263 1772 30309 1818
rect 30379 1772 30425 1818
rect 30495 1772 30541 1818
rect 30611 1772 30657 1818
rect 30727 1772 30773 1818
rect 30843 1772 30889 1818
rect 30959 1772 31005 1818
rect 31075 1772 31121 1818
rect 31191 1772 31237 1818
rect 31307 1772 31353 1818
rect 31423 1772 31469 1818
rect 31539 1772 31585 1818
rect 31655 1772 31701 1818
rect 31771 1772 31817 1818
rect 31887 1772 31933 1818
rect 32003 1772 32049 1818
rect 32119 1772 32165 1818
rect 32235 1772 32281 1818
rect 32351 1772 32397 1818
rect 32467 1772 32513 1818
rect 32583 1772 32629 1818
rect 32699 1772 32745 1818
rect 32815 1772 32861 1818
rect 32931 1772 32977 1818
rect 33047 1772 33093 1818
rect 33163 1772 33209 1818
rect 33279 1772 33325 1818
rect 33395 1772 33441 1818
rect 33511 1772 33557 1818
rect 33627 1772 33673 1818
rect 33743 1772 33789 1818
rect 33859 1772 33905 1818
rect 33975 1772 34021 1818
rect 34091 1772 34137 1818
rect 34207 1772 34253 1818
rect 34323 1772 34369 1818
rect 34439 1772 34485 1818
rect 34555 1772 34601 1818
rect 34671 1772 34717 1818
rect 34787 1772 34833 1818
rect 34903 1772 34949 1818
rect 35019 1772 35065 1818
rect 35135 1772 35181 1818
rect 35251 1772 35297 1818
rect 35367 1772 35413 1818
rect 35483 1772 35529 1818
rect 35599 1772 35645 1818
rect 35715 1772 35761 1818
rect 35831 1772 35877 1818
rect 35947 1772 35993 1818
rect 36063 1772 36109 1818
rect 36179 1772 36225 1818
rect 36295 1772 36341 1818
rect 36411 1772 36457 1818
rect 36527 1772 36573 1818
rect 36643 1772 36689 1818
rect 36759 1772 36805 1818
rect 36875 1772 36921 1818
rect 36991 1772 37037 1818
rect 37107 1772 37153 1818
rect 37223 1772 37269 1818
rect 37339 1772 37385 1818
rect 37455 1772 37501 1818
rect 37571 1772 37617 1818
rect 37687 1772 37733 1818
rect 37803 1772 37849 1818
rect 37919 1772 37965 1818
rect 38035 1772 38081 1818
rect 38151 1772 38197 1818
rect 38267 1772 38313 1818
rect 38383 1772 38429 1818
rect 38499 1772 38545 1818
rect 38615 1772 38661 1818
rect 38731 1772 38777 1818
rect 38847 1772 38893 1818
rect 38963 1772 39009 1818
rect 39079 1772 39125 1818
rect 39195 1772 39241 1818
rect 39311 1772 39357 1818
rect 39427 1772 39473 1818
rect 39543 1772 39589 1818
rect 39659 1772 39705 1818
rect 39775 1772 39821 1818
rect 39891 1772 39937 1818
rect 40007 1772 40053 1818
rect 40123 1772 40169 1818
rect 28639 1656 28685 1702
rect 28755 1656 28801 1702
rect 28871 1656 28917 1702
rect 28987 1656 29033 1702
rect 29103 1656 29149 1702
rect 29219 1656 29265 1702
rect 29335 1656 29381 1702
rect 29451 1656 29497 1702
rect 29567 1656 29613 1702
rect 29683 1656 29729 1702
rect 29799 1656 29845 1702
rect 29915 1656 29961 1702
rect 30031 1656 30077 1702
rect 30147 1656 30193 1702
rect 30263 1656 30309 1702
rect 30379 1656 30425 1702
rect 30495 1656 30541 1702
rect 30611 1656 30657 1702
rect 30727 1656 30773 1702
rect 30843 1656 30889 1702
rect 30959 1656 31005 1702
rect 31075 1656 31121 1702
rect 31191 1656 31237 1702
rect 31307 1656 31353 1702
rect 31423 1656 31469 1702
rect 31539 1656 31585 1702
rect 31655 1656 31701 1702
rect 31771 1656 31817 1702
rect 31887 1656 31933 1702
rect 32003 1656 32049 1702
rect 32119 1656 32165 1702
rect 32235 1656 32281 1702
rect 32351 1656 32397 1702
rect 32467 1656 32513 1702
rect 32583 1656 32629 1702
rect 32699 1656 32745 1702
rect 32815 1656 32861 1702
rect 32931 1656 32977 1702
rect 33047 1656 33093 1702
rect 33163 1656 33209 1702
rect 33279 1656 33325 1702
rect 33395 1656 33441 1702
rect 33511 1656 33557 1702
rect 33627 1656 33673 1702
rect 33743 1656 33789 1702
rect 33859 1656 33905 1702
rect 33975 1656 34021 1702
rect 34091 1656 34137 1702
rect 34207 1656 34253 1702
rect 34323 1656 34369 1702
rect 34439 1656 34485 1702
rect 34555 1656 34601 1702
rect 34671 1656 34717 1702
rect 34787 1656 34833 1702
rect 34903 1656 34949 1702
rect 35019 1656 35065 1702
rect 35135 1656 35181 1702
rect 35251 1656 35297 1702
rect 35367 1656 35413 1702
rect 35483 1656 35529 1702
rect 35599 1656 35645 1702
rect 35715 1656 35761 1702
rect 35831 1656 35877 1702
rect 35947 1656 35993 1702
rect 36063 1656 36109 1702
rect 36179 1656 36225 1702
rect 36295 1656 36341 1702
rect 36411 1656 36457 1702
rect 36527 1656 36573 1702
rect 36643 1656 36689 1702
rect 36759 1656 36805 1702
rect 36875 1656 36921 1702
rect 36991 1656 37037 1702
rect 37107 1656 37153 1702
rect 37223 1656 37269 1702
rect 37339 1656 37385 1702
rect 37455 1656 37501 1702
rect 37571 1656 37617 1702
rect 37687 1656 37733 1702
rect 37803 1656 37849 1702
rect 37919 1656 37965 1702
rect 38035 1656 38081 1702
rect 38151 1656 38197 1702
rect 38267 1656 38313 1702
rect 38383 1656 38429 1702
rect 38499 1656 38545 1702
rect 38615 1656 38661 1702
rect 38731 1656 38777 1702
rect 38847 1656 38893 1702
rect 38963 1656 39009 1702
rect 39079 1656 39125 1702
rect 39195 1656 39241 1702
rect 39311 1656 39357 1702
rect 39427 1656 39473 1702
rect 39543 1656 39589 1702
rect 39659 1656 39705 1702
rect 39775 1656 39821 1702
rect 39891 1656 39937 1702
rect 40007 1656 40053 1702
rect 40123 1656 40169 1702
rect 50845 3860 50891 3906
rect 50961 3860 51007 3906
rect 51077 3860 51123 3906
rect 51193 3860 51239 3906
rect 51309 3860 51355 3906
rect 51425 3860 51471 3906
rect 51541 3860 51587 3906
rect 51657 3860 51703 3906
rect 51773 3860 51819 3906
rect 51889 3860 51935 3906
rect 52005 3860 52051 3906
rect 52121 3860 52167 3906
rect 52237 3860 52283 3906
rect 52353 3860 52399 3906
rect 52469 3860 52515 3906
rect 52585 3860 52631 3906
rect 52701 3860 52747 3906
rect 52817 3860 52863 3906
rect 52933 3860 52979 3906
rect 53049 3860 53095 3906
rect 53165 3860 53211 3906
rect 53281 3860 53327 3906
rect 53397 3860 53443 3906
rect 53513 3860 53559 3906
rect 53629 3860 53675 3906
rect 53745 3860 53791 3906
rect 53861 3860 53907 3906
rect 53977 3860 54023 3906
rect 54093 3860 54139 3906
rect 54209 3860 54255 3906
rect 54325 3860 54371 3906
rect 54441 3860 54487 3906
rect 54557 3860 54603 3906
rect 54673 3860 54719 3906
rect 54789 3860 54835 3906
rect 54905 3860 54951 3906
rect 55021 3860 55067 3906
rect 55137 3860 55183 3906
rect 55253 3860 55299 3906
rect 55369 3860 55415 3906
rect 55485 3860 55531 3906
rect 55601 3860 55647 3906
rect 55717 3860 55763 3906
rect 55833 3860 55879 3906
rect 55949 3860 55995 3906
rect 56065 3860 56111 3906
rect 56181 3860 56227 3906
rect 56297 3860 56343 3906
rect 56413 3860 56459 3906
rect 56529 3860 56575 3906
rect 50845 3744 50891 3790
rect 50961 3744 51007 3790
rect 51077 3744 51123 3790
rect 51193 3744 51239 3790
rect 51309 3744 51355 3790
rect 51425 3744 51471 3790
rect 51541 3744 51587 3790
rect 51657 3744 51703 3790
rect 51773 3744 51819 3790
rect 51889 3744 51935 3790
rect 52005 3744 52051 3790
rect 52121 3744 52167 3790
rect 52237 3744 52283 3790
rect 52353 3744 52399 3790
rect 52469 3744 52515 3790
rect 52585 3744 52631 3790
rect 52701 3744 52747 3790
rect 52817 3744 52863 3790
rect 52933 3744 52979 3790
rect 53049 3744 53095 3790
rect 53165 3744 53211 3790
rect 53281 3744 53327 3790
rect 53397 3744 53443 3790
rect 53513 3744 53559 3790
rect 53629 3744 53675 3790
rect 53745 3744 53791 3790
rect 53861 3744 53907 3790
rect 53977 3744 54023 3790
rect 54093 3744 54139 3790
rect 54209 3744 54255 3790
rect 54325 3744 54371 3790
rect 54441 3744 54487 3790
rect 54557 3744 54603 3790
rect 54673 3744 54719 3790
rect 54789 3744 54835 3790
rect 54905 3744 54951 3790
rect 55021 3744 55067 3790
rect 55137 3744 55183 3790
rect 55253 3744 55299 3790
rect 55369 3744 55415 3790
rect 55485 3744 55531 3790
rect 55601 3744 55647 3790
rect 55717 3744 55763 3790
rect 55833 3744 55879 3790
rect 55949 3744 55995 3790
rect 56065 3744 56111 3790
rect 56181 3744 56227 3790
rect 56297 3744 56343 3790
rect 56413 3744 56459 3790
rect 56529 3744 56575 3790
rect 50845 3628 50891 3674
rect 50961 3628 51007 3674
rect 51077 3628 51123 3674
rect 51193 3628 51239 3674
rect 51309 3628 51355 3674
rect 51425 3628 51471 3674
rect 51541 3628 51587 3674
rect 51657 3628 51703 3674
rect 51773 3628 51819 3674
rect 51889 3628 51935 3674
rect 52005 3628 52051 3674
rect 52121 3628 52167 3674
rect 52237 3628 52283 3674
rect 52353 3628 52399 3674
rect 52469 3628 52515 3674
rect 52585 3628 52631 3674
rect 52701 3628 52747 3674
rect 52817 3628 52863 3674
rect 52933 3628 52979 3674
rect 53049 3628 53095 3674
rect 53165 3628 53211 3674
rect 53281 3628 53327 3674
rect 53397 3628 53443 3674
rect 53513 3628 53559 3674
rect 53629 3628 53675 3674
rect 53745 3628 53791 3674
rect 53861 3628 53907 3674
rect 53977 3628 54023 3674
rect 54093 3628 54139 3674
rect 54209 3628 54255 3674
rect 54325 3628 54371 3674
rect 54441 3628 54487 3674
rect 54557 3628 54603 3674
rect 54673 3628 54719 3674
rect 54789 3628 54835 3674
rect 54905 3628 54951 3674
rect 55021 3628 55067 3674
rect 55137 3628 55183 3674
rect 55253 3628 55299 3674
rect 55369 3628 55415 3674
rect 55485 3628 55531 3674
rect 55601 3628 55647 3674
rect 55717 3628 55763 3674
rect 55833 3628 55879 3674
rect 55949 3628 55995 3674
rect 56065 3628 56111 3674
rect 56181 3628 56227 3674
rect 56297 3628 56343 3674
rect 56413 3628 56459 3674
rect 56529 3628 56575 3674
rect 50845 3512 50891 3558
rect 50961 3512 51007 3558
rect 51077 3512 51123 3558
rect 51193 3512 51239 3558
rect 51309 3512 51355 3558
rect 51425 3512 51471 3558
rect 51541 3512 51587 3558
rect 51657 3512 51703 3558
rect 51773 3512 51819 3558
rect 51889 3512 51935 3558
rect 52005 3512 52051 3558
rect 52121 3512 52167 3558
rect 52237 3512 52283 3558
rect 52353 3512 52399 3558
rect 52469 3512 52515 3558
rect 52585 3512 52631 3558
rect 52701 3512 52747 3558
rect 52817 3512 52863 3558
rect 52933 3512 52979 3558
rect 53049 3512 53095 3558
rect 53165 3512 53211 3558
rect 53281 3512 53327 3558
rect 53397 3512 53443 3558
rect 53513 3512 53559 3558
rect 53629 3512 53675 3558
rect 53745 3512 53791 3558
rect 53861 3512 53907 3558
rect 53977 3512 54023 3558
rect 54093 3512 54139 3558
rect 54209 3512 54255 3558
rect 54325 3512 54371 3558
rect 54441 3512 54487 3558
rect 54557 3512 54603 3558
rect 54673 3512 54719 3558
rect 54789 3512 54835 3558
rect 54905 3512 54951 3558
rect 55021 3512 55067 3558
rect 55137 3512 55183 3558
rect 55253 3512 55299 3558
rect 55369 3512 55415 3558
rect 55485 3512 55531 3558
rect 55601 3512 55647 3558
rect 55717 3512 55763 3558
rect 55833 3512 55879 3558
rect 55949 3512 55995 3558
rect 56065 3512 56111 3558
rect 56181 3512 56227 3558
rect 56297 3512 56343 3558
rect 56413 3512 56459 3558
rect 56529 3512 56575 3558
rect 50845 3396 50891 3442
rect 50961 3396 51007 3442
rect 51077 3396 51123 3442
rect 51193 3396 51239 3442
rect 51309 3396 51355 3442
rect 51425 3396 51471 3442
rect 51541 3396 51587 3442
rect 51657 3396 51703 3442
rect 51773 3396 51819 3442
rect 51889 3396 51935 3442
rect 52005 3396 52051 3442
rect 52121 3396 52167 3442
rect 52237 3396 52283 3442
rect 52353 3396 52399 3442
rect 52469 3396 52515 3442
rect 52585 3396 52631 3442
rect 52701 3396 52747 3442
rect 52817 3396 52863 3442
rect 52933 3396 52979 3442
rect 53049 3396 53095 3442
rect 53165 3396 53211 3442
rect 53281 3396 53327 3442
rect 53397 3396 53443 3442
rect 53513 3396 53559 3442
rect 53629 3396 53675 3442
rect 53745 3396 53791 3442
rect 53861 3396 53907 3442
rect 53977 3396 54023 3442
rect 54093 3396 54139 3442
rect 54209 3396 54255 3442
rect 54325 3396 54371 3442
rect 54441 3396 54487 3442
rect 54557 3396 54603 3442
rect 54673 3396 54719 3442
rect 54789 3396 54835 3442
rect 54905 3396 54951 3442
rect 55021 3396 55067 3442
rect 55137 3396 55183 3442
rect 55253 3396 55299 3442
rect 55369 3396 55415 3442
rect 55485 3396 55531 3442
rect 55601 3396 55647 3442
rect 55717 3396 55763 3442
rect 55833 3396 55879 3442
rect 55949 3396 55995 3442
rect 56065 3396 56111 3442
rect 56181 3396 56227 3442
rect 56297 3396 56343 3442
rect 56413 3396 56459 3442
rect 56529 3396 56575 3442
rect 50845 3280 50891 3326
rect 50961 3280 51007 3326
rect 51077 3280 51123 3326
rect 51193 3280 51239 3326
rect 51309 3280 51355 3326
rect 51425 3280 51471 3326
rect 51541 3280 51587 3326
rect 51657 3280 51703 3326
rect 51773 3280 51819 3326
rect 51889 3280 51935 3326
rect 52005 3280 52051 3326
rect 52121 3280 52167 3326
rect 52237 3280 52283 3326
rect 52353 3280 52399 3326
rect 52469 3280 52515 3326
rect 52585 3280 52631 3326
rect 52701 3280 52747 3326
rect 52817 3280 52863 3326
rect 52933 3280 52979 3326
rect 53049 3280 53095 3326
rect 53165 3280 53211 3326
rect 53281 3280 53327 3326
rect 53397 3280 53443 3326
rect 53513 3280 53559 3326
rect 53629 3280 53675 3326
rect 53745 3280 53791 3326
rect 53861 3280 53907 3326
rect 53977 3280 54023 3326
rect 54093 3280 54139 3326
rect 54209 3280 54255 3326
rect 54325 3280 54371 3326
rect 54441 3280 54487 3326
rect 54557 3280 54603 3326
rect 54673 3280 54719 3326
rect 54789 3280 54835 3326
rect 54905 3280 54951 3326
rect 55021 3280 55067 3326
rect 55137 3280 55183 3326
rect 55253 3280 55299 3326
rect 55369 3280 55415 3326
rect 55485 3280 55531 3326
rect 55601 3280 55647 3326
rect 55717 3280 55763 3326
rect 55833 3280 55879 3326
rect 55949 3280 55995 3326
rect 56065 3280 56111 3326
rect 56181 3280 56227 3326
rect 56297 3280 56343 3326
rect 56413 3280 56459 3326
rect 56529 3280 56575 3326
rect 50845 3164 50891 3210
rect 50961 3164 51007 3210
rect 51077 3164 51123 3210
rect 51193 3164 51239 3210
rect 51309 3164 51355 3210
rect 51425 3164 51471 3210
rect 51541 3164 51587 3210
rect 51657 3164 51703 3210
rect 51773 3164 51819 3210
rect 51889 3164 51935 3210
rect 52005 3164 52051 3210
rect 52121 3164 52167 3210
rect 52237 3164 52283 3210
rect 52353 3164 52399 3210
rect 52469 3164 52515 3210
rect 52585 3164 52631 3210
rect 52701 3164 52747 3210
rect 52817 3164 52863 3210
rect 52933 3164 52979 3210
rect 53049 3164 53095 3210
rect 53165 3164 53211 3210
rect 53281 3164 53327 3210
rect 53397 3164 53443 3210
rect 53513 3164 53559 3210
rect 53629 3164 53675 3210
rect 53745 3164 53791 3210
rect 53861 3164 53907 3210
rect 53977 3164 54023 3210
rect 54093 3164 54139 3210
rect 54209 3164 54255 3210
rect 54325 3164 54371 3210
rect 54441 3164 54487 3210
rect 54557 3164 54603 3210
rect 54673 3164 54719 3210
rect 54789 3164 54835 3210
rect 54905 3164 54951 3210
rect 55021 3164 55067 3210
rect 55137 3164 55183 3210
rect 55253 3164 55299 3210
rect 55369 3164 55415 3210
rect 55485 3164 55531 3210
rect 55601 3164 55647 3210
rect 55717 3164 55763 3210
rect 55833 3164 55879 3210
rect 55949 3164 55995 3210
rect 56065 3164 56111 3210
rect 56181 3164 56227 3210
rect 56297 3164 56343 3210
rect 56413 3164 56459 3210
rect 56529 3164 56575 3210
rect 50845 3048 50891 3094
rect 50961 3048 51007 3094
rect 51077 3048 51123 3094
rect 51193 3048 51239 3094
rect 51309 3048 51355 3094
rect 51425 3048 51471 3094
rect 51541 3048 51587 3094
rect 51657 3048 51703 3094
rect 51773 3048 51819 3094
rect 51889 3048 51935 3094
rect 52005 3048 52051 3094
rect 52121 3048 52167 3094
rect 52237 3048 52283 3094
rect 52353 3048 52399 3094
rect 52469 3048 52515 3094
rect 52585 3048 52631 3094
rect 52701 3048 52747 3094
rect 52817 3048 52863 3094
rect 52933 3048 52979 3094
rect 53049 3048 53095 3094
rect 53165 3048 53211 3094
rect 53281 3048 53327 3094
rect 53397 3048 53443 3094
rect 53513 3048 53559 3094
rect 53629 3048 53675 3094
rect 53745 3048 53791 3094
rect 53861 3048 53907 3094
rect 53977 3048 54023 3094
rect 54093 3048 54139 3094
rect 54209 3048 54255 3094
rect 54325 3048 54371 3094
rect 54441 3048 54487 3094
rect 54557 3048 54603 3094
rect 54673 3048 54719 3094
rect 54789 3048 54835 3094
rect 54905 3048 54951 3094
rect 55021 3048 55067 3094
rect 55137 3048 55183 3094
rect 55253 3048 55299 3094
rect 55369 3048 55415 3094
rect 55485 3048 55531 3094
rect 55601 3048 55647 3094
rect 55717 3048 55763 3094
rect 55833 3048 55879 3094
rect 55949 3048 55995 3094
rect 56065 3048 56111 3094
rect 56181 3048 56227 3094
rect 56297 3048 56343 3094
rect 56413 3048 56459 3094
rect 56529 3048 56575 3094
rect 50845 2932 50891 2978
rect 50961 2932 51007 2978
rect 51077 2932 51123 2978
rect 51193 2932 51239 2978
rect 51309 2932 51355 2978
rect 51425 2932 51471 2978
rect 51541 2932 51587 2978
rect 51657 2932 51703 2978
rect 51773 2932 51819 2978
rect 51889 2932 51935 2978
rect 52005 2932 52051 2978
rect 52121 2932 52167 2978
rect 52237 2932 52283 2978
rect 52353 2932 52399 2978
rect 52469 2932 52515 2978
rect 52585 2932 52631 2978
rect 52701 2932 52747 2978
rect 52817 2932 52863 2978
rect 52933 2932 52979 2978
rect 53049 2932 53095 2978
rect 53165 2932 53211 2978
rect 53281 2932 53327 2978
rect 53397 2932 53443 2978
rect 53513 2932 53559 2978
rect 53629 2932 53675 2978
rect 53745 2932 53791 2978
rect 53861 2932 53907 2978
rect 53977 2932 54023 2978
rect 54093 2932 54139 2978
rect 54209 2932 54255 2978
rect 54325 2932 54371 2978
rect 54441 2932 54487 2978
rect 54557 2932 54603 2978
rect 54673 2932 54719 2978
rect 54789 2932 54835 2978
rect 54905 2932 54951 2978
rect 55021 2932 55067 2978
rect 55137 2932 55183 2978
rect 55253 2932 55299 2978
rect 55369 2932 55415 2978
rect 55485 2932 55531 2978
rect 55601 2932 55647 2978
rect 55717 2932 55763 2978
rect 55833 2932 55879 2978
rect 55949 2932 55995 2978
rect 56065 2932 56111 2978
rect 56181 2932 56227 2978
rect 56297 2932 56343 2978
rect 56413 2932 56459 2978
rect 56529 2932 56575 2978
rect 50845 2816 50891 2862
rect 50961 2816 51007 2862
rect 51077 2816 51123 2862
rect 51193 2816 51239 2862
rect 51309 2816 51355 2862
rect 51425 2816 51471 2862
rect 51541 2816 51587 2862
rect 51657 2816 51703 2862
rect 51773 2816 51819 2862
rect 51889 2816 51935 2862
rect 52005 2816 52051 2862
rect 52121 2816 52167 2862
rect 52237 2816 52283 2862
rect 52353 2816 52399 2862
rect 52469 2816 52515 2862
rect 52585 2816 52631 2862
rect 52701 2816 52747 2862
rect 52817 2816 52863 2862
rect 52933 2816 52979 2862
rect 53049 2816 53095 2862
rect 53165 2816 53211 2862
rect 53281 2816 53327 2862
rect 53397 2816 53443 2862
rect 53513 2816 53559 2862
rect 53629 2816 53675 2862
rect 53745 2816 53791 2862
rect 53861 2816 53907 2862
rect 53977 2816 54023 2862
rect 54093 2816 54139 2862
rect 54209 2816 54255 2862
rect 54325 2816 54371 2862
rect 54441 2816 54487 2862
rect 54557 2816 54603 2862
rect 54673 2816 54719 2862
rect 54789 2816 54835 2862
rect 54905 2816 54951 2862
rect 55021 2816 55067 2862
rect 55137 2816 55183 2862
rect 55253 2816 55299 2862
rect 55369 2816 55415 2862
rect 55485 2816 55531 2862
rect 55601 2816 55647 2862
rect 55717 2816 55763 2862
rect 55833 2816 55879 2862
rect 55949 2816 55995 2862
rect 56065 2816 56111 2862
rect 56181 2816 56227 2862
rect 56297 2816 56343 2862
rect 56413 2816 56459 2862
rect 56529 2816 56575 2862
rect 50845 2700 50891 2746
rect 50961 2700 51007 2746
rect 51077 2700 51123 2746
rect 51193 2700 51239 2746
rect 51309 2700 51355 2746
rect 51425 2700 51471 2746
rect 51541 2700 51587 2746
rect 51657 2700 51703 2746
rect 51773 2700 51819 2746
rect 51889 2700 51935 2746
rect 52005 2700 52051 2746
rect 52121 2700 52167 2746
rect 52237 2700 52283 2746
rect 52353 2700 52399 2746
rect 52469 2700 52515 2746
rect 52585 2700 52631 2746
rect 52701 2700 52747 2746
rect 52817 2700 52863 2746
rect 52933 2700 52979 2746
rect 53049 2700 53095 2746
rect 53165 2700 53211 2746
rect 53281 2700 53327 2746
rect 53397 2700 53443 2746
rect 53513 2700 53559 2746
rect 53629 2700 53675 2746
rect 53745 2700 53791 2746
rect 53861 2700 53907 2746
rect 53977 2700 54023 2746
rect 54093 2700 54139 2746
rect 54209 2700 54255 2746
rect 54325 2700 54371 2746
rect 54441 2700 54487 2746
rect 54557 2700 54603 2746
rect 54673 2700 54719 2746
rect 54789 2700 54835 2746
rect 54905 2700 54951 2746
rect 55021 2700 55067 2746
rect 55137 2700 55183 2746
rect 55253 2700 55299 2746
rect 55369 2700 55415 2746
rect 55485 2700 55531 2746
rect 55601 2700 55647 2746
rect 55717 2700 55763 2746
rect 55833 2700 55879 2746
rect 55949 2700 55995 2746
rect 56065 2700 56111 2746
rect 56181 2700 56227 2746
rect 56297 2700 56343 2746
rect 56413 2700 56459 2746
rect 56529 2700 56575 2746
rect 50845 2584 50891 2630
rect 50961 2584 51007 2630
rect 51077 2584 51123 2630
rect 51193 2584 51239 2630
rect 51309 2584 51355 2630
rect 51425 2584 51471 2630
rect 51541 2584 51587 2630
rect 51657 2584 51703 2630
rect 51773 2584 51819 2630
rect 51889 2584 51935 2630
rect 52005 2584 52051 2630
rect 52121 2584 52167 2630
rect 52237 2584 52283 2630
rect 52353 2584 52399 2630
rect 52469 2584 52515 2630
rect 52585 2584 52631 2630
rect 52701 2584 52747 2630
rect 52817 2584 52863 2630
rect 52933 2584 52979 2630
rect 53049 2584 53095 2630
rect 53165 2584 53211 2630
rect 53281 2584 53327 2630
rect 53397 2584 53443 2630
rect 53513 2584 53559 2630
rect 53629 2584 53675 2630
rect 53745 2584 53791 2630
rect 53861 2584 53907 2630
rect 53977 2584 54023 2630
rect 54093 2584 54139 2630
rect 54209 2584 54255 2630
rect 54325 2584 54371 2630
rect 54441 2584 54487 2630
rect 54557 2584 54603 2630
rect 54673 2584 54719 2630
rect 54789 2584 54835 2630
rect 54905 2584 54951 2630
rect 55021 2584 55067 2630
rect 55137 2584 55183 2630
rect 55253 2584 55299 2630
rect 55369 2584 55415 2630
rect 55485 2584 55531 2630
rect 55601 2584 55647 2630
rect 55717 2584 55763 2630
rect 55833 2584 55879 2630
rect 55949 2584 55995 2630
rect 56065 2584 56111 2630
rect 56181 2584 56227 2630
rect 56297 2584 56343 2630
rect 56413 2584 56459 2630
rect 56529 2584 56575 2630
rect 50845 2468 50891 2514
rect 50961 2468 51007 2514
rect 51077 2468 51123 2514
rect 51193 2468 51239 2514
rect 51309 2468 51355 2514
rect 51425 2468 51471 2514
rect 51541 2468 51587 2514
rect 51657 2468 51703 2514
rect 51773 2468 51819 2514
rect 51889 2468 51935 2514
rect 52005 2468 52051 2514
rect 52121 2468 52167 2514
rect 52237 2468 52283 2514
rect 52353 2468 52399 2514
rect 52469 2468 52515 2514
rect 52585 2468 52631 2514
rect 52701 2468 52747 2514
rect 52817 2468 52863 2514
rect 52933 2468 52979 2514
rect 53049 2468 53095 2514
rect 53165 2468 53211 2514
rect 53281 2468 53327 2514
rect 53397 2468 53443 2514
rect 53513 2468 53559 2514
rect 53629 2468 53675 2514
rect 53745 2468 53791 2514
rect 53861 2468 53907 2514
rect 53977 2468 54023 2514
rect 54093 2468 54139 2514
rect 54209 2468 54255 2514
rect 54325 2468 54371 2514
rect 54441 2468 54487 2514
rect 54557 2468 54603 2514
rect 54673 2468 54719 2514
rect 54789 2468 54835 2514
rect 54905 2468 54951 2514
rect 55021 2468 55067 2514
rect 55137 2468 55183 2514
rect 55253 2468 55299 2514
rect 55369 2468 55415 2514
rect 55485 2468 55531 2514
rect 55601 2468 55647 2514
rect 55717 2468 55763 2514
rect 55833 2468 55879 2514
rect 55949 2468 55995 2514
rect 56065 2468 56111 2514
rect 56181 2468 56227 2514
rect 56297 2468 56343 2514
rect 56413 2468 56459 2514
rect 56529 2468 56575 2514
rect 50845 2352 50891 2398
rect 50961 2352 51007 2398
rect 51077 2352 51123 2398
rect 51193 2352 51239 2398
rect 51309 2352 51355 2398
rect 51425 2352 51471 2398
rect 51541 2352 51587 2398
rect 51657 2352 51703 2398
rect 51773 2352 51819 2398
rect 51889 2352 51935 2398
rect 52005 2352 52051 2398
rect 52121 2352 52167 2398
rect 52237 2352 52283 2398
rect 52353 2352 52399 2398
rect 52469 2352 52515 2398
rect 52585 2352 52631 2398
rect 52701 2352 52747 2398
rect 52817 2352 52863 2398
rect 52933 2352 52979 2398
rect 53049 2352 53095 2398
rect 53165 2352 53211 2398
rect 53281 2352 53327 2398
rect 53397 2352 53443 2398
rect 53513 2352 53559 2398
rect 53629 2352 53675 2398
rect 53745 2352 53791 2398
rect 53861 2352 53907 2398
rect 53977 2352 54023 2398
rect 54093 2352 54139 2398
rect 54209 2352 54255 2398
rect 54325 2352 54371 2398
rect 54441 2352 54487 2398
rect 54557 2352 54603 2398
rect 54673 2352 54719 2398
rect 54789 2352 54835 2398
rect 54905 2352 54951 2398
rect 55021 2352 55067 2398
rect 55137 2352 55183 2398
rect 55253 2352 55299 2398
rect 55369 2352 55415 2398
rect 55485 2352 55531 2398
rect 55601 2352 55647 2398
rect 55717 2352 55763 2398
rect 55833 2352 55879 2398
rect 55949 2352 55995 2398
rect 56065 2352 56111 2398
rect 56181 2352 56227 2398
rect 56297 2352 56343 2398
rect 56413 2352 56459 2398
rect 56529 2352 56575 2398
rect 50845 2236 50891 2282
rect 50961 2236 51007 2282
rect 51077 2236 51123 2282
rect 51193 2236 51239 2282
rect 51309 2236 51355 2282
rect 51425 2236 51471 2282
rect 51541 2236 51587 2282
rect 51657 2236 51703 2282
rect 51773 2236 51819 2282
rect 51889 2236 51935 2282
rect 52005 2236 52051 2282
rect 52121 2236 52167 2282
rect 52237 2236 52283 2282
rect 52353 2236 52399 2282
rect 52469 2236 52515 2282
rect 52585 2236 52631 2282
rect 52701 2236 52747 2282
rect 52817 2236 52863 2282
rect 52933 2236 52979 2282
rect 53049 2236 53095 2282
rect 53165 2236 53211 2282
rect 53281 2236 53327 2282
rect 53397 2236 53443 2282
rect 53513 2236 53559 2282
rect 53629 2236 53675 2282
rect 53745 2236 53791 2282
rect 53861 2236 53907 2282
rect 53977 2236 54023 2282
rect 54093 2236 54139 2282
rect 54209 2236 54255 2282
rect 54325 2236 54371 2282
rect 54441 2236 54487 2282
rect 54557 2236 54603 2282
rect 54673 2236 54719 2282
rect 54789 2236 54835 2282
rect 54905 2236 54951 2282
rect 55021 2236 55067 2282
rect 55137 2236 55183 2282
rect 55253 2236 55299 2282
rect 55369 2236 55415 2282
rect 55485 2236 55531 2282
rect 55601 2236 55647 2282
rect 55717 2236 55763 2282
rect 55833 2236 55879 2282
rect 55949 2236 55995 2282
rect 56065 2236 56111 2282
rect 56181 2236 56227 2282
rect 56297 2236 56343 2282
rect 56413 2236 56459 2282
rect 56529 2236 56575 2282
rect 50845 2120 50891 2166
rect 50961 2120 51007 2166
rect 51077 2120 51123 2166
rect 51193 2120 51239 2166
rect 51309 2120 51355 2166
rect 51425 2120 51471 2166
rect 51541 2120 51587 2166
rect 51657 2120 51703 2166
rect 51773 2120 51819 2166
rect 51889 2120 51935 2166
rect 52005 2120 52051 2166
rect 52121 2120 52167 2166
rect 52237 2120 52283 2166
rect 52353 2120 52399 2166
rect 52469 2120 52515 2166
rect 52585 2120 52631 2166
rect 52701 2120 52747 2166
rect 52817 2120 52863 2166
rect 52933 2120 52979 2166
rect 53049 2120 53095 2166
rect 53165 2120 53211 2166
rect 53281 2120 53327 2166
rect 53397 2120 53443 2166
rect 53513 2120 53559 2166
rect 53629 2120 53675 2166
rect 53745 2120 53791 2166
rect 53861 2120 53907 2166
rect 53977 2120 54023 2166
rect 54093 2120 54139 2166
rect 54209 2120 54255 2166
rect 54325 2120 54371 2166
rect 54441 2120 54487 2166
rect 54557 2120 54603 2166
rect 54673 2120 54719 2166
rect 54789 2120 54835 2166
rect 54905 2120 54951 2166
rect 55021 2120 55067 2166
rect 55137 2120 55183 2166
rect 55253 2120 55299 2166
rect 55369 2120 55415 2166
rect 55485 2120 55531 2166
rect 55601 2120 55647 2166
rect 55717 2120 55763 2166
rect 55833 2120 55879 2166
rect 55949 2120 55995 2166
rect 56065 2120 56111 2166
rect 56181 2120 56227 2166
rect 56297 2120 56343 2166
rect 56413 2120 56459 2166
rect 56529 2120 56575 2166
rect 50845 2004 50891 2050
rect 50961 2004 51007 2050
rect 51077 2004 51123 2050
rect 51193 2004 51239 2050
rect 51309 2004 51355 2050
rect 51425 2004 51471 2050
rect 51541 2004 51587 2050
rect 51657 2004 51703 2050
rect 51773 2004 51819 2050
rect 51889 2004 51935 2050
rect 52005 2004 52051 2050
rect 52121 2004 52167 2050
rect 52237 2004 52283 2050
rect 52353 2004 52399 2050
rect 52469 2004 52515 2050
rect 52585 2004 52631 2050
rect 52701 2004 52747 2050
rect 52817 2004 52863 2050
rect 52933 2004 52979 2050
rect 53049 2004 53095 2050
rect 53165 2004 53211 2050
rect 53281 2004 53327 2050
rect 53397 2004 53443 2050
rect 53513 2004 53559 2050
rect 53629 2004 53675 2050
rect 53745 2004 53791 2050
rect 53861 2004 53907 2050
rect 53977 2004 54023 2050
rect 54093 2004 54139 2050
rect 54209 2004 54255 2050
rect 54325 2004 54371 2050
rect 54441 2004 54487 2050
rect 54557 2004 54603 2050
rect 54673 2004 54719 2050
rect 54789 2004 54835 2050
rect 54905 2004 54951 2050
rect 55021 2004 55067 2050
rect 55137 2004 55183 2050
rect 55253 2004 55299 2050
rect 55369 2004 55415 2050
rect 55485 2004 55531 2050
rect 55601 2004 55647 2050
rect 55717 2004 55763 2050
rect 55833 2004 55879 2050
rect 55949 2004 55995 2050
rect 56065 2004 56111 2050
rect 56181 2004 56227 2050
rect 56297 2004 56343 2050
rect 56413 2004 56459 2050
rect 56529 2004 56575 2050
rect 50845 1888 50891 1934
rect 50961 1888 51007 1934
rect 51077 1888 51123 1934
rect 51193 1888 51239 1934
rect 51309 1888 51355 1934
rect 51425 1888 51471 1934
rect 51541 1888 51587 1934
rect 51657 1888 51703 1934
rect 51773 1888 51819 1934
rect 51889 1888 51935 1934
rect 52005 1888 52051 1934
rect 52121 1888 52167 1934
rect 52237 1888 52283 1934
rect 52353 1888 52399 1934
rect 52469 1888 52515 1934
rect 52585 1888 52631 1934
rect 52701 1888 52747 1934
rect 52817 1888 52863 1934
rect 52933 1888 52979 1934
rect 53049 1888 53095 1934
rect 53165 1888 53211 1934
rect 53281 1888 53327 1934
rect 53397 1888 53443 1934
rect 53513 1888 53559 1934
rect 53629 1888 53675 1934
rect 53745 1888 53791 1934
rect 53861 1888 53907 1934
rect 53977 1888 54023 1934
rect 54093 1888 54139 1934
rect 54209 1888 54255 1934
rect 54325 1888 54371 1934
rect 54441 1888 54487 1934
rect 54557 1888 54603 1934
rect 54673 1888 54719 1934
rect 54789 1888 54835 1934
rect 54905 1888 54951 1934
rect 55021 1888 55067 1934
rect 55137 1888 55183 1934
rect 55253 1888 55299 1934
rect 55369 1888 55415 1934
rect 55485 1888 55531 1934
rect 55601 1888 55647 1934
rect 55717 1888 55763 1934
rect 55833 1888 55879 1934
rect 55949 1888 55995 1934
rect 56065 1888 56111 1934
rect 56181 1888 56227 1934
rect 56297 1888 56343 1934
rect 56413 1888 56459 1934
rect 56529 1888 56575 1934
rect 50845 1772 50891 1818
rect 50961 1772 51007 1818
rect 51077 1772 51123 1818
rect 51193 1772 51239 1818
rect 51309 1772 51355 1818
rect 51425 1772 51471 1818
rect 51541 1772 51587 1818
rect 51657 1772 51703 1818
rect 51773 1772 51819 1818
rect 51889 1772 51935 1818
rect 52005 1772 52051 1818
rect 52121 1772 52167 1818
rect 52237 1772 52283 1818
rect 52353 1772 52399 1818
rect 52469 1772 52515 1818
rect 52585 1772 52631 1818
rect 52701 1772 52747 1818
rect 52817 1772 52863 1818
rect 52933 1772 52979 1818
rect 53049 1772 53095 1818
rect 53165 1772 53211 1818
rect 53281 1772 53327 1818
rect 53397 1772 53443 1818
rect 53513 1772 53559 1818
rect 53629 1772 53675 1818
rect 53745 1772 53791 1818
rect 53861 1772 53907 1818
rect 53977 1772 54023 1818
rect 54093 1772 54139 1818
rect 54209 1772 54255 1818
rect 54325 1772 54371 1818
rect 54441 1772 54487 1818
rect 54557 1772 54603 1818
rect 54673 1772 54719 1818
rect 54789 1772 54835 1818
rect 54905 1772 54951 1818
rect 55021 1772 55067 1818
rect 55137 1772 55183 1818
rect 55253 1772 55299 1818
rect 55369 1772 55415 1818
rect 55485 1772 55531 1818
rect 55601 1772 55647 1818
rect 55717 1772 55763 1818
rect 55833 1772 55879 1818
rect 55949 1772 55995 1818
rect 56065 1772 56111 1818
rect 56181 1772 56227 1818
rect 56297 1772 56343 1818
rect 56413 1772 56459 1818
rect 56529 1772 56575 1818
rect 50845 1656 50891 1702
rect 50961 1656 51007 1702
rect 51077 1656 51123 1702
rect 51193 1656 51239 1702
rect 51309 1656 51355 1702
rect 51425 1656 51471 1702
rect 51541 1656 51587 1702
rect 51657 1656 51703 1702
rect 51773 1656 51819 1702
rect 51889 1656 51935 1702
rect 52005 1656 52051 1702
rect 52121 1656 52167 1702
rect 52237 1656 52283 1702
rect 52353 1656 52399 1702
rect 52469 1656 52515 1702
rect 52585 1656 52631 1702
rect 52701 1656 52747 1702
rect 52817 1656 52863 1702
rect 52933 1656 52979 1702
rect 53049 1656 53095 1702
rect 53165 1656 53211 1702
rect 53281 1656 53327 1702
rect 53397 1656 53443 1702
rect 53513 1656 53559 1702
rect 53629 1656 53675 1702
rect 53745 1656 53791 1702
rect 53861 1656 53907 1702
rect 53977 1656 54023 1702
rect 54093 1656 54139 1702
rect 54209 1656 54255 1702
rect 54325 1656 54371 1702
rect 54441 1656 54487 1702
rect 54557 1656 54603 1702
rect 54673 1656 54719 1702
rect 54789 1656 54835 1702
rect 54905 1656 54951 1702
rect 55021 1656 55067 1702
rect 55137 1656 55183 1702
rect 55253 1656 55299 1702
rect 55369 1656 55415 1702
rect 55485 1656 55531 1702
rect 55601 1656 55647 1702
rect 55717 1656 55763 1702
rect 55833 1656 55879 1702
rect 55949 1656 55995 1702
rect 56065 1656 56111 1702
rect 56181 1656 56227 1702
rect 56297 1656 56343 1702
rect 56413 1656 56459 1702
rect 56529 1656 56575 1702
<< mvnsubdiffcont >>
rect 30854 65790 30900 65836
rect 31012 65790 31058 65836
rect 31170 65790 31216 65836
rect 31328 65790 31374 65836
rect 31487 65790 31533 65836
rect 31645 65790 31691 65836
rect 31803 65790 31849 65836
rect 31961 65790 32007 65836
rect 32119 65790 32165 65836
rect 32277 65790 32323 65836
rect 32435 65790 32481 65836
rect 32593 65790 32639 65836
rect 42717 65863 42763 65909
rect 42875 65863 42921 65909
rect 43033 65863 43079 65909
rect 43191 65863 43237 65909
rect 43350 65863 43396 65909
rect 43508 65863 43554 65909
rect 30637 65676 30683 65722
rect 30854 65627 30900 65673
rect 31012 65627 31058 65673
rect 31170 65627 31216 65673
rect 31328 65627 31374 65673
rect 31487 65627 31533 65673
rect 31645 65627 31691 65673
rect 31803 65627 31849 65673
rect 31961 65627 32007 65673
rect 32119 65627 32165 65673
rect 32277 65627 32323 65673
rect 32435 65627 32481 65673
rect 32593 65627 32639 65673
rect 30637 65512 30683 65558
rect 30854 65463 30900 65509
rect 31012 65463 31058 65509
rect 31170 65463 31216 65509
rect 31328 65463 31374 65509
rect 31487 65463 31533 65509
rect 31645 65463 31691 65509
rect 31803 65463 31849 65509
rect 31961 65463 32007 65509
rect 32119 65463 32165 65509
rect 32277 65463 32323 65509
rect 32435 65463 32481 65509
rect 32593 65463 32639 65509
rect 52483 65790 52529 65836
rect 52641 65790 52687 65836
rect 52799 65790 52845 65836
rect 52957 65790 53003 65836
rect 53115 65790 53161 65836
rect 53273 65790 53319 65836
rect 53431 65790 53477 65836
rect 53589 65790 53635 65836
rect 53748 65790 53794 65836
rect 53906 65790 53952 65836
rect 54064 65790 54110 65836
rect 54222 65790 54268 65836
rect 30637 65349 30683 65395
rect 30854 65300 30900 65346
rect 31012 65300 31058 65346
rect 31170 65300 31216 65346
rect 31328 65300 31374 65346
rect 31487 65300 31533 65346
rect 31645 65300 31691 65346
rect 31803 65300 31849 65346
rect 31961 65300 32007 65346
rect 32119 65300 32165 65346
rect 32277 65300 32323 65346
rect 32435 65300 32481 65346
rect 32593 65300 32639 65346
rect 54440 65676 54486 65722
rect 52483 65627 52529 65673
rect 52641 65627 52687 65673
rect 52799 65627 52845 65673
rect 52957 65627 53003 65673
rect 53115 65627 53161 65673
rect 53273 65627 53319 65673
rect 53431 65627 53477 65673
rect 53589 65627 53635 65673
rect 53748 65627 53794 65673
rect 53906 65627 53952 65673
rect 54064 65627 54110 65673
rect 54222 65627 54268 65673
rect 54440 65512 54486 65558
rect 52483 65463 52529 65509
rect 52641 65463 52687 65509
rect 52799 65463 52845 65509
rect 52957 65463 53003 65509
rect 53115 65463 53161 65509
rect 53273 65463 53319 65509
rect 53431 65463 53477 65509
rect 53589 65463 53635 65509
rect 53748 65463 53794 65509
rect 53906 65463 53952 65509
rect 54064 65463 54110 65509
rect 54222 65463 54268 65509
rect 54440 65349 54486 65395
rect 52483 65300 52529 65346
rect 52641 65300 52687 65346
rect 52799 65300 52845 65346
rect 52957 65300 53003 65346
rect 53115 65300 53161 65346
rect 53273 65300 53319 65346
rect 53431 65300 53477 65346
rect 53589 65300 53635 65346
rect 53748 65300 53794 65346
rect 53906 65300 53952 65346
rect 54064 65300 54110 65346
rect 54222 65300 54268 65346
rect 30637 65186 30683 65232
rect 30637 65022 30683 65068
rect 54440 65186 54486 65232
rect 54440 65022 54486 65068
rect 36489 64904 36723 64950
rect 30637 64820 30683 64866
rect 30855 64780 30901 64826
rect 30637 64657 30683 64703
rect 30855 64616 30901 64662
rect 30637 64494 30683 64540
rect 30855 64453 30901 64499
rect 30637 64331 30683 64377
rect 30855 64290 30901 64336
rect 39062 64904 39108 64950
rect 39220 64904 39266 64950
rect 45619 64904 45665 64950
rect 45777 64904 45823 64950
rect 45935 64904 45981 64950
rect 46093 64904 46139 64950
rect 46251 64904 46297 64950
rect 46409 64904 46455 64950
rect 46568 64904 46614 64950
rect 46726 64904 46772 64950
rect 46884 64904 46930 64950
rect 47042 64904 47088 64950
rect 47200 64904 47246 64950
rect 47358 64904 47404 64950
rect 47516 64904 47562 64950
rect 47675 64904 47721 64950
rect 47833 64904 47879 64950
rect 47991 64904 48037 64950
rect 48149 64904 48195 64950
rect 48307 64904 48353 64950
rect 48465 64904 48511 64950
rect 45619 64740 45665 64786
rect 45777 64740 45823 64786
rect 45935 64740 45981 64786
rect 46093 64740 46139 64786
rect 46251 64740 46297 64786
rect 46409 64740 46455 64786
rect 46568 64740 46614 64786
rect 46726 64740 46772 64786
rect 46884 64740 46930 64786
rect 47042 64740 47088 64786
rect 47200 64740 47246 64786
rect 47358 64740 47404 64786
rect 47516 64740 47562 64786
rect 47675 64740 47721 64786
rect 47833 64740 47879 64786
rect 47991 64740 48037 64786
rect 48149 64740 48195 64786
rect 48307 64740 48353 64786
rect 48465 64740 48511 64786
rect 54223 64780 54269 64826
rect 54440 64820 54486 64866
rect 30637 64167 30683 64213
rect 30855 64127 30901 64173
rect 54223 64616 54269 64662
rect 54440 64657 54486 64703
rect 54440 64494 54486 64540
rect 54440 64331 54486 64377
rect 54223 64127 54269 64173
rect 54440 64167 54486 64213
rect 30637 64004 30683 64050
rect 54440 64004 54486 64050
rect 30637 63841 30683 63887
rect 30855 63881 30901 63927
rect 30637 63677 30683 63723
rect 30855 63718 30901 63764
rect 30637 63514 30683 63560
rect 30855 63555 30901 63601
rect 30637 63351 30683 63397
rect 30855 63392 30901 63438
rect 30637 63188 30683 63234
rect 30855 63228 30901 63274
rect 54223 63881 54269 63927
rect 54440 63841 54486 63887
rect 36489 63104 36723 63150
rect 30637 63020 30683 63066
rect 30855 62980 30901 63026
rect 30637 62857 30683 62903
rect 30855 62816 30901 62862
rect 30637 62694 30683 62740
rect 30855 62653 30901 62699
rect 30637 62531 30683 62577
rect 30855 62490 30901 62536
rect 39062 63104 39108 63150
rect 39220 63104 39266 63150
rect 45619 63268 45665 63314
rect 45777 63268 45823 63314
rect 45935 63268 45981 63314
rect 46093 63268 46139 63314
rect 46251 63268 46297 63314
rect 46409 63268 46455 63314
rect 46568 63268 46614 63314
rect 46726 63268 46772 63314
rect 46884 63268 46930 63314
rect 47042 63268 47088 63314
rect 47200 63268 47246 63314
rect 47358 63268 47404 63314
rect 47516 63268 47562 63314
rect 47675 63268 47721 63314
rect 47833 63268 47879 63314
rect 47991 63268 48037 63314
rect 48149 63268 48195 63314
rect 48307 63268 48353 63314
rect 48465 63268 48511 63314
rect 54440 63677 54486 63723
rect 54440 63514 54486 63560
rect 54223 63392 54269 63438
rect 54440 63351 54486 63397
rect 54223 63228 54269 63274
rect 54440 63188 54486 63234
rect 45619 63104 45665 63150
rect 45777 63104 45823 63150
rect 45935 63104 45981 63150
rect 46093 63104 46139 63150
rect 46251 63104 46297 63150
rect 46409 63104 46455 63150
rect 46568 63104 46614 63150
rect 46726 63104 46772 63150
rect 46884 63104 46930 63150
rect 47042 63104 47088 63150
rect 47200 63104 47246 63150
rect 47358 63104 47404 63150
rect 47516 63104 47562 63150
rect 47675 63104 47721 63150
rect 47833 63104 47879 63150
rect 47991 63104 48037 63150
rect 48149 63104 48195 63150
rect 48307 63104 48353 63150
rect 48465 63104 48511 63150
rect 45619 62940 45665 62986
rect 45777 62940 45823 62986
rect 45935 62940 45981 62986
rect 46093 62940 46139 62986
rect 46251 62940 46297 62986
rect 46409 62940 46455 62986
rect 46568 62940 46614 62986
rect 46726 62940 46772 62986
rect 46884 62940 46930 62986
rect 47042 62940 47088 62986
rect 47200 62940 47246 62986
rect 47358 62940 47404 62986
rect 47516 62940 47562 62986
rect 47675 62940 47721 62986
rect 47833 62940 47879 62986
rect 47991 62940 48037 62986
rect 48149 62940 48195 62986
rect 48307 62940 48353 62986
rect 48465 62940 48511 62986
rect 54223 62980 54269 63026
rect 54440 63020 54486 63066
rect 30637 62367 30683 62413
rect 30855 62327 30901 62373
rect 54223 62816 54269 62862
rect 54440 62857 54486 62903
rect 54440 62694 54486 62740
rect 54440 62531 54486 62577
rect 54223 62327 54269 62373
rect 54440 62367 54486 62413
rect 30637 62204 30683 62250
rect 54440 62204 54486 62250
rect 30637 62041 30683 62087
rect 30855 62081 30901 62127
rect 30637 61877 30683 61923
rect 30855 61918 30901 61964
rect 30637 61714 30683 61760
rect 30855 61755 30901 61801
rect 30637 61551 30683 61597
rect 30855 61592 30901 61638
rect 30637 61388 30683 61434
rect 30855 61428 30901 61474
rect 54223 62081 54269 62127
rect 54440 62041 54486 62087
rect 36489 61304 36723 61350
rect 30637 61220 30683 61266
rect 30855 61180 30901 61226
rect 30637 61057 30683 61103
rect 30855 61016 30901 61062
rect 30637 60894 30683 60940
rect 30855 60853 30901 60899
rect 30637 60731 30683 60777
rect 30855 60690 30901 60736
rect 39062 61304 39108 61350
rect 39220 61304 39266 61350
rect 45619 61468 45665 61514
rect 45777 61468 45823 61514
rect 45935 61468 45981 61514
rect 46093 61468 46139 61514
rect 46251 61468 46297 61514
rect 46409 61468 46455 61514
rect 46568 61468 46614 61514
rect 46726 61468 46772 61514
rect 46884 61468 46930 61514
rect 47042 61468 47088 61514
rect 47200 61468 47246 61514
rect 47358 61468 47404 61514
rect 47516 61468 47562 61514
rect 47675 61468 47721 61514
rect 47833 61468 47879 61514
rect 47991 61468 48037 61514
rect 48149 61468 48195 61514
rect 48307 61468 48353 61514
rect 48465 61468 48511 61514
rect 54440 61877 54486 61923
rect 54440 61714 54486 61760
rect 54223 61592 54269 61638
rect 54440 61551 54486 61597
rect 54223 61428 54269 61474
rect 54440 61388 54486 61434
rect 45619 61304 45665 61350
rect 45777 61304 45823 61350
rect 45935 61304 45981 61350
rect 46093 61304 46139 61350
rect 46251 61304 46297 61350
rect 46409 61304 46455 61350
rect 46568 61304 46614 61350
rect 46726 61304 46772 61350
rect 46884 61304 46930 61350
rect 47042 61304 47088 61350
rect 47200 61304 47246 61350
rect 47358 61304 47404 61350
rect 47516 61304 47562 61350
rect 47675 61304 47721 61350
rect 47833 61304 47879 61350
rect 47991 61304 48037 61350
rect 48149 61304 48195 61350
rect 48307 61304 48353 61350
rect 48465 61304 48511 61350
rect 45619 61140 45665 61186
rect 45777 61140 45823 61186
rect 45935 61140 45981 61186
rect 46093 61140 46139 61186
rect 46251 61140 46297 61186
rect 46409 61140 46455 61186
rect 46568 61140 46614 61186
rect 46726 61140 46772 61186
rect 46884 61140 46930 61186
rect 47042 61140 47088 61186
rect 47200 61140 47246 61186
rect 47358 61140 47404 61186
rect 47516 61140 47562 61186
rect 47675 61140 47721 61186
rect 47833 61140 47879 61186
rect 47991 61140 48037 61186
rect 48149 61140 48195 61186
rect 48307 61140 48353 61186
rect 48465 61140 48511 61186
rect 54223 61180 54269 61226
rect 54440 61220 54486 61266
rect 30637 60567 30683 60613
rect 30855 60527 30901 60573
rect 54223 61016 54269 61062
rect 54440 61057 54486 61103
rect 54440 60894 54486 60940
rect 54440 60731 54486 60777
rect 54223 60527 54269 60573
rect 54440 60567 54486 60613
rect 30637 60404 30683 60450
rect 54440 60404 54486 60450
rect 30637 60241 30683 60287
rect 30855 60281 30901 60327
rect 30637 60077 30683 60123
rect 30855 60118 30901 60164
rect 30637 59914 30683 59960
rect 30855 59955 30901 60001
rect 30637 59751 30683 59797
rect 30855 59792 30901 59838
rect 30637 59588 30683 59634
rect 30855 59628 30901 59674
rect 54223 60281 54269 60327
rect 54440 60241 54486 60287
rect 36489 59504 36723 59550
rect 30637 59420 30683 59466
rect 30855 59380 30901 59426
rect 30637 59257 30683 59303
rect 30855 59216 30901 59262
rect 30637 59094 30683 59140
rect 30855 59053 30901 59099
rect 30637 58931 30683 58977
rect 30855 58890 30901 58936
rect 39062 59504 39108 59550
rect 39220 59504 39266 59550
rect 45619 59668 45665 59714
rect 45777 59668 45823 59714
rect 45935 59668 45981 59714
rect 46093 59668 46139 59714
rect 46251 59668 46297 59714
rect 46409 59668 46455 59714
rect 46568 59668 46614 59714
rect 46726 59668 46772 59714
rect 46884 59668 46930 59714
rect 47042 59668 47088 59714
rect 47200 59668 47246 59714
rect 47358 59668 47404 59714
rect 47516 59668 47562 59714
rect 47675 59668 47721 59714
rect 47833 59668 47879 59714
rect 47991 59668 48037 59714
rect 48149 59668 48195 59714
rect 48307 59668 48353 59714
rect 48465 59668 48511 59714
rect 54440 60077 54486 60123
rect 54440 59914 54486 59960
rect 54223 59792 54269 59838
rect 54440 59751 54486 59797
rect 54223 59628 54269 59674
rect 54440 59588 54486 59634
rect 45619 59504 45665 59550
rect 45777 59504 45823 59550
rect 45935 59504 45981 59550
rect 46093 59504 46139 59550
rect 46251 59504 46297 59550
rect 46409 59504 46455 59550
rect 46568 59504 46614 59550
rect 46726 59504 46772 59550
rect 46884 59504 46930 59550
rect 47042 59504 47088 59550
rect 47200 59504 47246 59550
rect 47358 59504 47404 59550
rect 47516 59504 47562 59550
rect 47675 59504 47721 59550
rect 47833 59504 47879 59550
rect 47991 59504 48037 59550
rect 48149 59504 48195 59550
rect 48307 59504 48353 59550
rect 48465 59504 48511 59550
rect 45619 59340 45665 59386
rect 45777 59340 45823 59386
rect 45935 59340 45981 59386
rect 46093 59340 46139 59386
rect 46251 59340 46297 59386
rect 46409 59340 46455 59386
rect 46568 59340 46614 59386
rect 46726 59340 46772 59386
rect 46884 59340 46930 59386
rect 47042 59340 47088 59386
rect 47200 59340 47246 59386
rect 47358 59340 47404 59386
rect 47516 59340 47562 59386
rect 47675 59340 47721 59386
rect 47833 59340 47879 59386
rect 47991 59340 48037 59386
rect 48149 59340 48195 59386
rect 48307 59340 48353 59386
rect 48465 59340 48511 59386
rect 54223 59380 54269 59426
rect 54440 59420 54486 59466
rect 30637 58767 30683 58813
rect 30855 58727 30901 58773
rect 54223 59216 54269 59262
rect 54440 59257 54486 59303
rect 54440 59094 54486 59140
rect 54440 58931 54486 58977
rect 54223 58727 54269 58773
rect 54440 58767 54486 58813
rect 30637 58604 30683 58650
rect 54440 58604 54486 58650
rect 30637 58441 30683 58487
rect 30855 58481 30901 58527
rect 30637 58277 30683 58323
rect 30855 58318 30901 58364
rect 30637 58114 30683 58160
rect 30855 58155 30901 58201
rect 30637 57951 30683 57997
rect 30855 57992 30901 58038
rect 30637 57788 30683 57834
rect 30855 57828 30901 57874
rect 54223 58481 54269 58527
rect 54440 58441 54486 58487
rect 36489 57704 36723 57750
rect 30637 57620 30683 57666
rect 30855 57580 30901 57626
rect 30637 57457 30683 57503
rect 30855 57416 30901 57462
rect 30637 57294 30683 57340
rect 30855 57253 30901 57299
rect 30637 57131 30683 57177
rect 30855 57090 30901 57136
rect 39062 57704 39108 57750
rect 39220 57704 39266 57750
rect 45619 57868 45665 57914
rect 45777 57868 45823 57914
rect 45935 57868 45981 57914
rect 46093 57868 46139 57914
rect 46251 57868 46297 57914
rect 46409 57868 46455 57914
rect 46568 57868 46614 57914
rect 46726 57868 46772 57914
rect 46884 57868 46930 57914
rect 47042 57868 47088 57914
rect 47200 57868 47246 57914
rect 47358 57868 47404 57914
rect 47516 57868 47562 57914
rect 47675 57868 47721 57914
rect 47833 57868 47879 57914
rect 47991 57868 48037 57914
rect 48149 57868 48195 57914
rect 48307 57868 48353 57914
rect 48465 57868 48511 57914
rect 54440 58277 54486 58323
rect 54440 58114 54486 58160
rect 54223 57992 54269 58038
rect 54440 57951 54486 57997
rect 54223 57828 54269 57874
rect 54440 57788 54486 57834
rect 45619 57704 45665 57750
rect 45777 57704 45823 57750
rect 45935 57704 45981 57750
rect 46093 57704 46139 57750
rect 46251 57704 46297 57750
rect 46409 57704 46455 57750
rect 46568 57704 46614 57750
rect 46726 57704 46772 57750
rect 46884 57704 46930 57750
rect 47042 57704 47088 57750
rect 47200 57704 47246 57750
rect 47358 57704 47404 57750
rect 47516 57704 47562 57750
rect 47675 57704 47721 57750
rect 47833 57704 47879 57750
rect 47991 57704 48037 57750
rect 48149 57704 48195 57750
rect 48307 57704 48353 57750
rect 48465 57704 48511 57750
rect 45619 57540 45665 57586
rect 45777 57540 45823 57586
rect 45935 57540 45981 57586
rect 46093 57540 46139 57586
rect 46251 57540 46297 57586
rect 46409 57540 46455 57586
rect 46568 57540 46614 57586
rect 46726 57540 46772 57586
rect 46884 57540 46930 57586
rect 47042 57540 47088 57586
rect 47200 57540 47246 57586
rect 47358 57540 47404 57586
rect 47516 57540 47562 57586
rect 47675 57540 47721 57586
rect 47833 57540 47879 57586
rect 47991 57540 48037 57586
rect 48149 57540 48195 57586
rect 48307 57540 48353 57586
rect 48465 57540 48511 57586
rect 54223 57580 54269 57626
rect 54440 57620 54486 57666
rect 30637 56967 30683 57013
rect 30855 56927 30901 56973
rect 54223 57416 54269 57462
rect 54440 57457 54486 57503
rect 54440 57294 54486 57340
rect 54440 57131 54486 57177
rect 54223 56927 54269 56973
rect 54440 56967 54486 57013
rect 30637 56804 30683 56850
rect 54440 56804 54486 56850
rect 30637 56641 30683 56687
rect 30855 56681 30901 56727
rect 30637 56477 30683 56523
rect 30855 56518 30901 56564
rect 30637 56314 30683 56360
rect 30855 56355 30901 56401
rect 30637 56151 30683 56197
rect 30855 56192 30901 56238
rect 30637 55988 30683 56034
rect 30855 56028 30901 56074
rect 54223 56681 54269 56727
rect 54440 56641 54486 56687
rect 36489 55904 36723 55950
rect 30637 55820 30683 55866
rect 30855 55780 30901 55826
rect 30637 55657 30683 55703
rect 30855 55616 30901 55662
rect 30637 55494 30683 55540
rect 30855 55453 30901 55499
rect 30637 55331 30683 55377
rect 30855 55290 30901 55336
rect 39062 55904 39108 55950
rect 39220 55904 39266 55950
rect 45619 56068 45665 56114
rect 45777 56068 45823 56114
rect 45935 56068 45981 56114
rect 46093 56068 46139 56114
rect 46251 56068 46297 56114
rect 46409 56068 46455 56114
rect 46568 56068 46614 56114
rect 46726 56068 46772 56114
rect 46884 56068 46930 56114
rect 47042 56068 47088 56114
rect 47200 56068 47246 56114
rect 47358 56068 47404 56114
rect 47516 56068 47562 56114
rect 47675 56068 47721 56114
rect 47833 56068 47879 56114
rect 47991 56068 48037 56114
rect 48149 56068 48195 56114
rect 48307 56068 48353 56114
rect 48465 56068 48511 56114
rect 54440 56477 54486 56523
rect 54440 56314 54486 56360
rect 54223 56192 54269 56238
rect 54440 56151 54486 56197
rect 54223 56028 54269 56074
rect 54440 55988 54486 56034
rect 45619 55904 45665 55950
rect 45777 55904 45823 55950
rect 45935 55904 45981 55950
rect 46093 55904 46139 55950
rect 46251 55904 46297 55950
rect 46409 55904 46455 55950
rect 46568 55904 46614 55950
rect 46726 55904 46772 55950
rect 46884 55904 46930 55950
rect 47042 55904 47088 55950
rect 47200 55904 47246 55950
rect 47358 55904 47404 55950
rect 47516 55904 47562 55950
rect 47675 55904 47721 55950
rect 47833 55904 47879 55950
rect 47991 55904 48037 55950
rect 48149 55904 48195 55950
rect 48307 55904 48353 55950
rect 48465 55904 48511 55950
rect 45619 55740 45665 55786
rect 45777 55740 45823 55786
rect 45935 55740 45981 55786
rect 46093 55740 46139 55786
rect 46251 55740 46297 55786
rect 46409 55740 46455 55786
rect 46568 55740 46614 55786
rect 46726 55740 46772 55786
rect 46884 55740 46930 55786
rect 47042 55740 47088 55786
rect 47200 55740 47246 55786
rect 47358 55740 47404 55786
rect 47516 55740 47562 55786
rect 47675 55740 47721 55786
rect 47833 55740 47879 55786
rect 47991 55740 48037 55786
rect 48149 55740 48195 55786
rect 48307 55740 48353 55786
rect 48465 55740 48511 55786
rect 54223 55780 54269 55826
rect 54440 55820 54486 55866
rect 30637 55167 30683 55213
rect 30855 55127 30901 55173
rect 54223 55616 54269 55662
rect 54440 55657 54486 55703
rect 54440 55494 54486 55540
rect 54440 55331 54486 55377
rect 54223 55127 54269 55173
rect 54440 55167 54486 55213
rect 30637 55004 30683 55050
rect 54440 55004 54486 55050
rect 30637 54841 30683 54887
rect 30855 54881 30901 54927
rect 30637 54677 30683 54723
rect 30855 54718 30901 54764
rect 30637 54514 30683 54560
rect 30855 54555 30901 54601
rect 30637 54351 30683 54397
rect 30855 54392 30901 54438
rect 30637 54188 30683 54234
rect 30855 54228 30901 54274
rect 54223 54881 54269 54927
rect 54440 54841 54486 54887
rect 36489 54104 36723 54150
rect 30637 54020 30683 54066
rect 30855 53980 30901 54026
rect 30637 53857 30683 53903
rect 30855 53816 30901 53862
rect 30637 53694 30683 53740
rect 30855 53653 30901 53699
rect 30637 53531 30683 53577
rect 30855 53490 30901 53536
rect 39062 54104 39108 54150
rect 39220 54104 39266 54150
rect 45619 54268 45665 54314
rect 45777 54268 45823 54314
rect 45935 54268 45981 54314
rect 46093 54268 46139 54314
rect 46251 54268 46297 54314
rect 46409 54268 46455 54314
rect 46568 54268 46614 54314
rect 46726 54268 46772 54314
rect 46884 54268 46930 54314
rect 47042 54268 47088 54314
rect 47200 54268 47246 54314
rect 47358 54268 47404 54314
rect 47516 54268 47562 54314
rect 47675 54268 47721 54314
rect 47833 54268 47879 54314
rect 47991 54268 48037 54314
rect 48149 54268 48195 54314
rect 48307 54268 48353 54314
rect 48465 54268 48511 54314
rect 54440 54677 54486 54723
rect 54440 54514 54486 54560
rect 54223 54392 54269 54438
rect 54440 54351 54486 54397
rect 54223 54228 54269 54274
rect 54440 54188 54486 54234
rect 45619 54104 45665 54150
rect 45777 54104 45823 54150
rect 45935 54104 45981 54150
rect 46093 54104 46139 54150
rect 46251 54104 46297 54150
rect 46409 54104 46455 54150
rect 46568 54104 46614 54150
rect 46726 54104 46772 54150
rect 46884 54104 46930 54150
rect 47042 54104 47088 54150
rect 47200 54104 47246 54150
rect 47358 54104 47404 54150
rect 47516 54104 47562 54150
rect 47675 54104 47721 54150
rect 47833 54104 47879 54150
rect 47991 54104 48037 54150
rect 48149 54104 48195 54150
rect 48307 54104 48353 54150
rect 48465 54104 48511 54150
rect 45619 53940 45665 53986
rect 45777 53940 45823 53986
rect 45935 53940 45981 53986
rect 46093 53940 46139 53986
rect 46251 53940 46297 53986
rect 46409 53940 46455 53986
rect 46568 53940 46614 53986
rect 46726 53940 46772 53986
rect 46884 53940 46930 53986
rect 47042 53940 47088 53986
rect 47200 53940 47246 53986
rect 47358 53940 47404 53986
rect 47516 53940 47562 53986
rect 47675 53940 47721 53986
rect 47833 53940 47879 53986
rect 47991 53940 48037 53986
rect 48149 53940 48195 53986
rect 48307 53940 48353 53986
rect 48465 53940 48511 53986
rect 54223 53980 54269 54026
rect 54440 54020 54486 54066
rect 30637 53367 30683 53413
rect 30855 53327 30901 53373
rect 54223 53816 54269 53862
rect 54440 53857 54486 53903
rect 54440 53694 54486 53740
rect 54440 53531 54486 53577
rect 54223 53327 54269 53373
rect 54440 53367 54486 53413
rect 30637 53204 30683 53250
rect 54440 53204 54486 53250
rect 30637 53041 30683 53087
rect 30855 53081 30901 53127
rect 30637 52877 30683 52923
rect 30855 52918 30901 52964
rect 30637 52714 30683 52760
rect 30855 52755 30901 52801
rect 30637 52551 30683 52597
rect 30855 52592 30901 52638
rect 30637 52388 30683 52434
rect 30855 52428 30901 52474
rect 54223 53081 54269 53127
rect 54440 53041 54486 53087
rect 36489 52304 36723 52350
rect 30637 52220 30683 52266
rect 30855 52180 30901 52226
rect 30637 52057 30683 52103
rect 30855 52016 30901 52062
rect 30637 51894 30683 51940
rect 30855 51853 30901 51899
rect 30637 51731 30683 51777
rect 30855 51690 30901 51736
rect 39062 52304 39108 52350
rect 39220 52304 39266 52350
rect 45619 52468 45665 52514
rect 45777 52468 45823 52514
rect 45935 52468 45981 52514
rect 46093 52468 46139 52514
rect 46251 52468 46297 52514
rect 46409 52468 46455 52514
rect 46568 52468 46614 52514
rect 46726 52468 46772 52514
rect 46884 52468 46930 52514
rect 47042 52468 47088 52514
rect 47200 52468 47246 52514
rect 47358 52468 47404 52514
rect 47516 52468 47562 52514
rect 47675 52468 47721 52514
rect 47833 52468 47879 52514
rect 47991 52468 48037 52514
rect 48149 52468 48195 52514
rect 48307 52468 48353 52514
rect 48465 52468 48511 52514
rect 54440 52877 54486 52923
rect 54440 52714 54486 52760
rect 54223 52592 54269 52638
rect 54440 52551 54486 52597
rect 54223 52428 54269 52474
rect 54440 52388 54486 52434
rect 45619 52304 45665 52350
rect 45777 52304 45823 52350
rect 45935 52304 45981 52350
rect 46093 52304 46139 52350
rect 46251 52304 46297 52350
rect 46409 52304 46455 52350
rect 46568 52304 46614 52350
rect 46726 52304 46772 52350
rect 46884 52304 46930 52350
rect 47042 52304 47088 52350
rect 47200 52304 47246 52350
rect 47358 52304 47404 52350
rect 47516 52304 47562 52350
rect 47675 52304 47721 52350
rect 47833 52304 47879 52350
rect 47991 52304 48037 52350
rect 48149 52304 48195 52350
rect 48307 52304 48353 52350
rect 48465 52304 48511 52350
rect 45619 52140 45665 52186
rect 45777 52140 45823 52186
rect 45935 52140 45981 52186
rect 46093 52140 46139 52186
rect 46251 52140 46297 52186
rect 46409 52140 46455 52186
rect 46568 52140 46614 52186
rect 46726 52140 46772 52186
rect 46884 52140 46930 52186
rect 47042 52140 47088 52186
rect 47200 52140 47246 52186
rect 47358 52140 47404 52186
rect 47516 52140 47562 52186
rect 47675 52140 47721 52186
rect 47833 52140 47879 52186
rect 47991 52140 48037 52186
rect 48149 52140 48195 52186
rect 48307 52140 48353 52186
rect 48465 52140 48511 52186
rect 54223 52180 54269 52226
rect 54440 52220 54486 52266
rect 30637 51567 30683 51613
rect 30855 51527 30901 51573
rect 54223 52016 54269 52062
rect 54440 52057 54486 52103
rect 54440 51894 54486 51940
rect 54440 51731 54486 51777
rect 54223 51527 54269 51573
rect 54440 51567 54486 51613
rect 30637 51404 30683 51450
rect 54440 51404 54486 51450
rect 30637 51241 30683 51287
rect 30855 51281 30901 51327
rect 30637 51077 30683 51123
rect 30855 51118 30901 51164
rect 30637 50914 30683 50960
rect 30855 50955 30901 51001
rect 30637 50751 30683 50797
rect 30855 50792 30901 50838
rect 30637 50588 30683 50634
rect 30855 50628 30901 50674
rect 54223 51281 54269 51327
rect 54440 51241 54486 51287
rect 36489 50504 36723 50550
rect 30637 50420 30683 50466
rect 30855 50380 30901 50426
rect 30637 50257 30683 50303
rect 30855 50216 30901 50262
rect 30637 50094 30683 50140
rect 30855 50053 30901 50099
rect 30637 49931 30683 49977
rect 30855 49890 30901 49936
rect 39062 50504 39108 50550
rect 39220 50504 39266 50550
rect 45619 50668 45665 50714
rect 45777 50668 45823 50714
rect 45935 50668 45981 50714
rect 46093 50668 46139 50714
rect 46251 50668 46297 50714
rect 46409 50668 46455 50714
rect 46568 50668 46614 50714
rect 46726 50668 46772 50714
rect 46884 50668 46930 50714
rect 47042 50668 47088 50714
rect 47200 50668 47246 50714
rect 47358 50668 47404 50714
rect 47516 50668 47562 50714
rect 47675 50668 47721 50714
rect 47833 50668 47879 50714
rect 47991 50668 48037 50714
rect 48149 50668 48195 50714
rect 48307 50668 48353 50714
rect 48465 50668 48511 50714
rect 54440 51077 54486 51123
rect 54440 50914 54486 50960
rect 54223 50792 54269 50838
rect 54440 50751 54486 50797
rect 54223 50628 54269 50674
rect 54440 50588 54486 50634
rect 45619 50504 45665 50550
rect 45777 50504 45823 50550
rect 45935 50504 45981 50550
rect 46093 50504 46139 50550
rect 46251 50504 46297 50550
rect 46409 50504 46455 50550
rect 46568 50504 46614 50550
rect 46726 50504 46772 50550
rect 46884 50504 46930 50550
rect 47042 50504 47088 50550
rect 47200 50504 47246 50550
rect 47358 50504 47404 50550
rect 47516 50504 47562 50550
rect 47675 50504 47721 50550
rect 47833 50504 47879 50550
rect 47991 50504 48037 50550
rect 48149 50504 48195 50550
rect 48307 50504 48353 50550
rect 48465 50504 48511 50550
rect 45619 50340 45665 50386
rect 45777 50340 45823 50386
rect 45935 50340 45981 50386
rect 46093 50340 46139 50386
rect 46251 50340 46297 50386
rect 46409 50340 46455 50386
rect 46568 50340 46614 50386
rect 46726 50340 46772 50386
rect 46884 50340 46930 50386
rect 47042 50340 47088 50386
rect 47200 50340 47246 50386
rect 47358 50340 47404 50386
rect 47516 50340 47562 50386
rect 47675 50340 47721 50386
rect 47833 50340 47879 50386
rect 47991 50340 48037 50386
rect 48149 50340 48195 50386
rect 48307 50340 48353 50386
rect 48465 50340 48511 50386
rect 54223 50380 54269 50426
rect 54440 50420 54486 50466
rect 30637 49767 30683 49813
rect 30855 49727 30901 49773
rect 54223 50216 54269 50262
rect 54440 50257 54486 50303
rect 54440 50094 54486 50140
rect 54440 49931 54486 49977
rect 54223 49727 54269 49773
rect 54440 49767 54486 49813
rect 30637 49604 30683 49650
rect 54440 49604 54486 49650
rect 30637 49441 30683 49487
rect 30855 49481 30901 49527
rect 30637 49277 30683 49323
rect 30855 49318 30901 49364
rect 30637 49114 30683 49160
rect 30855 49155 30901 49201
rect 30637 48951 30683 48997
rect 30855 48992 30901 49038
rect 30637 48788 30683 48834
rect 30855 48828 30901 48874
rect 54223 49481 54269 49527
rect 54440 49441 54486 49487
rect 36489 48704 36723 48750
rect 30637 48620 30683 48666
rect 30855 48580 30901 48626
rect 30637 48457 30683 48503
rect 30855 48416 30901 48462
rect 30637 48294 30683 48340
rect 30855 48253 30901 48299
rect 30637 48131 30683 48177
rect 30855 48090 30901 48136
rect 39062 48704 39108 48750
rect 39220 48704 39266 48750
rect 45619 48868 45665 48914
rect 45777 48868 45823 48914
rect 45935 48868 45981 48914
rect 46093 48868 46139 48914
rect 46251 48868 46297 48914
rect 46409 48868 46455 48914
rect 46568 48868 46614 48914
rect 46726 48868 46772 48914
rect 46884 48868 46930 48914
rect 47042 48868 47088 48914
rect 47200 48868 47246 48914
rect 47358 48868 47404 48914
rect 47516 48868 47562 48914
rect 47675 48868 47721 48914
rect 47833 48868 47879 48914
rect 47991 48868 48037 48914
rect 48149 48868 48195 48914
rect 48307 48868 48353 48914
rect 48465 48868 48511 48914
rect 54440 49277 54486 49323
rect 54440 49114 54486 49160
rect 54223 48992 54269 49038
rect 54440 48951 54486 48997
rect 54223 48828 54269 48874
rect 54440 48788 54486 48834
rect 45619 48704 45665 48750
rect 45777 48704 45823 48750
rect 45935 48704 45981 48750
rect 46093 48704 46139 48750
rect 46251 48704 46297 48750
rect 46409 48704 46455 48750
rect 46568 48704 46614 48750
rect 46726 48704 46772 48750
rect 46884 48704 46930 48750
rect 47042 48704 47088 48750
rect 47200 48704 47246 48750
rect 47358 48704 47404 48750
rect 47516 48704 47562 48750
rect 47675 48704 47721 48750
rect 47833 48704 47879 48750
rect 47991 48704 48037 48750
rect 48149 48704 48195 48750
rect 48307 48704 48353 48750
rect 48465 48704 48511 48750
rect 45619 48540 45665 48586
rect 45777 48540 45823 48586
rect 45935 48540 45981 48586
rect 46093 48540 46139 48586
rect 46251 48540 46297 48586
rect 46409 48540 46455 48586
rect 46568 48540 46614 48586
rect 46726 48540 46772 48586
rect 46884 48540 46930 48586
rect 47042 48540 47088 48586
rect 47200 48540 47246 48586
rect 47358 48540 47404 48586
rect 47516 48540 47562 48586
rect 47675 48540 47721 48586
rect 47833 48540 47879 48586
rect 47991 48540 48037 48586
rect 48149 48540 48195 48586
rect 48307 48540 48353 48586
rect 48465 48540 48511 48586
rect 54223 48580 54269 48626
rect 54440 48620 54486 48666
rect 30637 47967 30683 48013
rect 30855 47927 30901 47973
rect 54223 48416 54269 48462
rect 54440 48457 54486 48503
rect 54440 48294 54486 48340
rect 54440 48131 54486 48177
rect 54223 47927 54269 47973
rect 54440 47967 54486 48013
rect 30637 47804 30683 47850
rect 54440 47804 54486 47850
rect 30637 47641 30683 47687
rect 30855 47681 30901 47727
rect 30637 47477 30683 47523
rect 30855 47518 30901 47564
rect 30637 47314 30683 47360
rect 30855 47355 30901 47401
rect 30637 47151 30683 47197
rect 30855 47192 30901 47238
rect 30637 46988 30683 47034
rect 30855 47028 30901 47074
rect 54223 47681 54269 47727
rect 54440 47641 54486 47687
rect 36489 46904 36723 46950
rect 30637 46820 30683 46866
rect 30855 46780 30901 46826
rect 30637 46657 30683 46703
rect 30855 46616 30901 46662
rect 30637 46494 30683 46540
rect 30855 46453 30901 46499
rect 30637 46331 30683 46377
rect 30855 46290 30901 46336
rect 39062 46904 39108 46950
rect 39220 46904 39266 46950
rect 45619 47068 45665 47114
rect 45777 47068 45823 47114
rect 45935 47068 45981 47114
rect 46093 47068 46139 47114
rect 46251 47068 46297 47114
rect 46409 47068 46455 47114
rect 46568 47068 46614 47114
rect 46726 47068 46772 47114
rect 46884 47068 46930 47114
rect 47042 47068 47088 47114
rect 47200 47068 47246 47114
rect 47358 47068 47404 47114
rect 47516 47068 47562 47114
rect 47675 47068 47721 47114
rect 47833 47068 47879 47114
rect 47991 47068 48037 47114
rect 48149 47068 48195 47114
rect 48307 47068 48353 47114
rect 48465 47068 48511 47114
rect 54440 47477 54486 47523
rect 54440 47314 54486 47360
rect 54223 47192 54269 47238
rect 54440 47151 54486 47197
rect 54223 47028 54269 47074
rect 54440 46988 54486 47034
rect 45619 46904 45665 46950
rect 45777 46904 45823 46950
rect 45935 46904 45981 46950
rect 46093 46904 46139 46950
rect 46251 46904 46297 46950
rect 46409 46904 46455 46950
rect 46568 46904 46614 46950
rect 46726 46904 46772 46950
rect 46884 46904 46930 46950
rect 47042 46904 47088 46950
rect 47200 46904 47246 46950
rect 47358 46904 47404 46950
rect 47516 46904 47562 46950
rect 47675 46904 47721 46950
rect 47833 46904 47879 46950
rect 47991 46904 48037 46950
rect 48149 46904 48195 46950
rect 48307 46904 48353 46950
rect 48465 46904 48511 46950
rect 45619 46740 45665 46786
rect 45777 46740 45823 46786
rect 45935 46740 45981 46786
rect 46093 46740 46139 46786
rect 46251 46740 46297 46786
rect 46409 46740 46455 46786
rect 46568 46740 46614 46786
rect 46726 46740 46772 46786
rect 46884 46740 46930 46786
rect 47042 46740 47088 46786
rect 47200 46740 47246 46786
rect 47358 46740 47404 46786
rect 47516 46740 47562 46786
rect 47675 46740 47721 46786
rect 47833 46740 47879 46786
rect 47991 46740 48037 46786
rect 48149 46740 48195 46786
rect 48307 46740 48353 46786
rect 48465 46740 48511 46786
rect 54223 46780 54269 46826
rect 54440 46820 54486 46866
rect 30637 46167 30683 46213
rect 30855 46127 30901 46173
rect 54223 46616 54269 46662
rect 54440 46657 54486 46703
rect 54440 46494 54486 46540
rect 54440 46331 54486 46377
rect 54223 46127 54269 46173
rect 54440 46167 54486 46213
rect 30637 46004 30683 46050
rect 54440 46004 54486 46050
rect 30637 45841 30683 45887
rect 30855 45881 30901 45927
rect 30637 45677 30683 45723
rect 30855 45718 30901 45764
rect 30637 45514 30683 45560
rect 30855 45555 30901 45601
rect 30637 45351 30683 45397
rect 30855 45392 30901 45438
rect 30637 45188 30683 45234
rect 30855 45228 30901 45274
rect 54223 45881 54269 45927
rect 54440 45841 54486 45887
rect 36489 45104 36723 45150
rect 30637 45020 30683 45066
rect 30855 44980 30901 45026
rect 30637 44857 30683 44903
rect 30855 44816 30901 44862
rect 30637 44694 30683 44740
rect 30855 44653 30901 44699
rect 30637 44531 30683 44577
rect 30855 44490 30901 44536
rect 39062 45104 39108 45150
rect 39220 45104 39266 45150
rect 45619 45268 45665 45314
rect 45777 45268 45823 45314
rect 45935 45268 45981 45314
rect 46093 45268 46139 45314
rect 46251 45268 46297 45314
rect 46409 45268 46455 45314
rect 46568 45268 46614 45314
rect 46726 45268 46772 45314
rect 46884 45268 46930 45314
rect 47042 45268 47088 45314
rect 47200 45268 47246 45314
rect 47358 45268 47404 45314
rect 47516 45268 47562 45314
rect 47675 45268 47721 45314
rect 47833 45268 47879 45314
rect 47991 45268 48037 45314
rect 48149 45268 48195 45314
rect 48307 45268 48353 45314
rect 48465 45268 48511 45314
rect 54440 45677 54486 45723
rect 54440 45514 54486 45560
rect 54223 45392 54269 45438
rect 54440 45351 54486 45397
rect 54223 45228 54269 45274
rect 54440 45188 54486 45234
rect 45619 45104 45665 45150
rect 45777 45104 45823 45150
rect 45935 45104 45981 45150
rect 46093 45104 46139 45150
rect 46251 45104 46297 45150
rect 46409 45104 46455 45150
rect 46568 45104 46614 45150
rect 46726 45104 46772 45150
rect 46884 45104 46930 45150
rect 47042 45104 47088 45150
rect 47200 45104 47246 45150
rect 47358 45104 47404 45150
rect 47516 45104 47562 45150
rect 47675 45104 47721 45150
rect 47833 45104 47879 45150
rect 47991 45104 48037 45150
rect 48149 45104 48195 45150
rect 48307 45104 48353 45150
rect 48465 45104 48511 45150
rect 45619 44940 45665 44986
rect 45777 44940 45823 44986
rect 45935 44940 45981 44986
rect 46093 44940 46139 44986
rect 46251 44940 46297 44986
rect 46409 44940 46455 44986
rect 46568 44940 46614 44986
rect 46726 44940 46772 44986
rect 46884 44940 46930 44986
rect 47042 44940 47088 44986
rect 47200 44940 47246 44986
rect 47358 44940 47404 44986
rect 47516 44940 47562 44986
rect 47675 44940 47721 44986
rect 47833 44940 47879 44986
rect 47991 44940 48037 44986
rect 48149 44940 48195 44986
rect 48307 44940 48353 44986
rect 48465 44940 48511 44986
rect 54223 44980 54269 45026
rect 54440 45020 54486 45066
rect 30637 44367 30683 44413
rect 30855 44327 30901 44373
rect 54223 44816 54269 44862
rect 54440 44857 54486 44903
rect 54440 44694 54486 44740
rect 54440 44531 54486 44577
rect 54223 44327 54269 44373
rect 54440 44367 54486 44413
rect 30637 44204 30683 44250
rect 54440 44204 54486 44250
rect 30637 44041 30683 44087
rect 30855 44081 30901 44127
rect 30637 43877 30683 43923
rect 30855 43918 30901 43964
rect 30637 43714 30683 43760
rect 30855 43755 30901 43801
rect 30637 43551 30683 43597
rect 30855 43592 30901 43638
rect 30637 43388 30683 43434
rect 30855 43428 30901 43474
rect 54223 44081 54269 44127
rect 54440 44041 54486 44087
rect 36489 43304 36723 43350
rect 30637 43220 30683 43266
rect 30855 43180 30901 43226
rect 30637 43057 30683 43103
rect 30855 43016 30901 43062
rect 30637 42894 30683 42940
rect 30855 42853 30901 42899
rect 30637 42731 30683 42777
rect 30855 42690 30901 42736
rect 39062 43304 39108 43350
rect 39220 43304 39266 43350
rect 45619 43468 45665 43514
rect 45777 43468 45823 43514
rect 45935 43468 45981 43514
rect 46093 43468 46139 43514
rect 46251 43468 46297 43514
rect 46409 43468 46455 43514
rect 46568 43468 46614 43514
rect 46726 43468 46772 43514
rect 46884 43468 46930 43514
rect 47042 43468 47088 43514
rect 47200 43468 47246 43514
rect 47358 43468 47404 43514
rect 47516 43468 47562 43514
rect 47675 43468 47721 43514
rect 47833 43468 47879 43514
rect 47991 43468 48037 43514
rect 48149 43468 48195 43514
rect 48307 43468 48353 43514
rect 48465 43468 48511 43514
rect 54440 43877 54486 43923
rect 54440 43714 54486 43760
rect 54223 43592 54269 43638
rect 54440 43551 54486 43597
rect 54223 43428 54269 43474
rect 54440 43388 54486 43434
rect 45619 43304 45665 43350
rect 45777 43304 45823 43350
rect 45935 43304 45981 43350
rect 46093 43304 46139 43350
rect 46251 43304 46297 43350
rect 46409 43304 46455 43350
rect 46568 43304 46614 43350
rect 46726 43304 46772 43350
rect 46884 43304 46930 43350
rect 47042 43304 47088 43350
rect 47200 43304 47246 43350
rect 47358 43304 47404 43350
rect 47516 43304 47562 43350
rect 47675 43304 47721 43350
rect 47833 43304 47879 43350
rect 47991 43304 48037 43350
rect 48149 43304 48195 43350
rect 48307 43304 48353 43350
rect 48465 43304 48511 43350
rect 45619 43140 45665 43186
rect 45777 43140 45823 43186
rect 45935 43140 45981 43186
rect 46093 43140 46139 43186
rect 46251 43140 46297 43186
rect 46409 43140 46455 43186
rect 46568 43140 46614 43186
rect 46726 43140 46772 43186
rect 46884 43140 46930 43186
rect 47042 43140 47088 43186
rect 47200 43140 47246 43186
rect 47358 43140 47404 43186
rect 47516 43140 47562 43186
rect 47675 43140 47721 43186
rect 47833 43140 47879 43186
rect 47991 43140 48037 43186
rect 48149 43140 48195 43186
rect 48307 43140 48353 43186
rect 48465 43140 48511 43186
rect 54223 43180 54269 43226
rect 54440 43220 54486 43266
rect 30637 42567 30683 42613
rect 30855 42527 30901 42573
rect 54223 43016 54269 43062
rect 54440 43057 54486 43103
rect 54440 42894 54486 42940
rect 54440 42731 54486 42777
rect 54223 42527 54269 42573
rect 54440 42567 54486 42613
rect 30637 42404 30683 42450
rect 54440 42404 54486 42450
rect 30637 42241 30683 42287
rect 30855 42281 30901 42327
rect 30637 42077 30683 42123
rect 30855 42118 30901 42164
rect 30637 41914 30683 41960
rect 30855 41955 30901 42001
rect 30637 41751 30683 41797
rect 30855 41792 30901 41838
rect 30637 41588 30683 41634
rect 30855 41628 30901 41674
rect 54223 42281 54269 42327
rect 54440 42241 54486 42287
rect 36489 41504 36723 41550
rect 30637 41420 30683 41466
rect 30855 41380 30901 41426
rect 30637 41257 30683 41303
rect 30855 41216 30901 41262
rect 30637 41094 30683 41140
rect 30855 41053 30901 41099
rect 30637 40931 30683 40977
rect 30855 40890 30901 40936
rect 39062 41504 39108 41550
rect 39220 41504 39266 41550
rect 45619 41668 45665 41714
rect 45777 41668 45823 41714
rect 45935 41668 45981 41714
rect 46093 41668 46139 41714
rect 46251 41668 46297 41714
rect 46409 41668 46455 41714
rect 46568 41668 46614 41714
rect 46726 41668 46772 41714
rect 46884 41668 46930 41714
rect 47042 41668 47088 41714
rect 47200 41668 47246 41714
rect 47358 41668 47404 41714
rect 47516 41668 47562 41714
rect 47675 41668 47721 41714
rect 47833 41668 47879 41714
rect 47991 41668 48037 41714
rect 48149 41668 48195 41714
rect 48307 41668 48353 41714
rect 48465 41668 48511 41714
rect 54440 42077 54486 42123
rect 54440 41914 54486 41960
rect 54223 41792 54269 41838
rect 54440 41751 54486 41797
rect 54223 41628 54269 41674
rect 54440 41588 54486 41634
rect 45619 41504 45665 41550
rect 45777 41504 45823 41550
rect 45935 41504 45981 41550
rect 46093 41504 46139 41550
rect 46251 41504 46297 41550
rect 46409 41504 46455 41550
rect 46568 41504 46614 41550
rect 46726 41504 46772 41550
rect 46884 41504 46930 41550
rect 47042 41504 47088 41550
rect 47200 41504 47246 41550
rect 47358 41504 47404 41550
rect 47516 41504 47562 41550
rect 47675 41504 47721 41550
rect 47833 41504 47879 41550
rect 47991 41504 48037 41550
rect 48149 41504 48195 41550
rect 48307 41504 48353 41550
rect 48465 41504 48511 41550
rect 45619 41340 45665 41386
rect 45777 41340 45823 41386
rect 45935 41340 45981 41386
rect 46093 41340 46139 41386
rect 46251 41340 46297 41386
rect 46409 41340 46455 41386
rect 46568 41340 46614 41386
rect 46726 41340 46772 41386
rect 46884 41340 46930 41386
rect 47042 41340 47088 41386
rect 47200 41340 47246 41386
rect 47358 41340 47404 41386
rect 47516 41340 47562 41386
rect 47675 41340 47721 41386
rect 47833 41340 47879 41386
rect 47991 41340 48037 41386
rect 48149 41340 48195 41386
rect 48307 41340 48353 41386
rect 48465 41340 48511 41386
rect 54223 41380 54269 41426
rect 54440 41420 54486 41466
rect 30637 40767 30683 40813
rect 30855 40727 30901 40773
rect 54223 41216 54269 41262
rect 54440 41257 54486 41303
rect 54440 41094 54486 41140
rect 54440 40931 54486 40977
rect 54223 40727 54269 40773
rect 54440 40767 54486 40813
rect 30637 40604 30683 40650
rect 54440 40604 54486 40650
rect 30637 40441 30683 40487
rect 30855 40481 30901 40527
rect 30637 40277 30683 40323
rect 30855 40318 30901 40364
rect 30637 40114 30683 40160
rect 30855 40155 30901 40201
rect 30637 39951 30683 39997
rect 30855 39992 30901 40038
rect 30637 39788 30683 39834
rect 30855 39828 30901 39874
rect 54223 40481 54269 40527
rect 54440 40441 54486 40487
rect 36489 39704 36723 39750
rect 30637 39620 30683 39666
rect 30855 39580 30901 39626
rect 30637 39457 30683 39503
rect 30855 39416 30901 39462
rect 30637 39294 30683 39340
rect 30855 39253 30901 39299
rect 30637 39131 30683 39177
rect 30855 39090 30901 39136
rect 39062 39704 39108 39750
rect 39220 39704 39266 39750
rect 45619 39868 45665 39914
rect 45777 39868 45823 39914
rect 45935 39868 45981 39914
rect 46093 39868 46139 39914
rect 46251 39868 46297 39914
rect 46409 39868 46455 39914
rect 46568 39868 46614 39914
rect 46726 39868 46772 39914
rect 46884 39868 46930 39914
rect 47042 39868 47088 39914
rect 47200 39868 47246 39914
rect 47358 39868 47404 39914
rect 47516 39868 47562 39914
rect 47675 39868 47721 39914
rect 47833 39868 47879 39914
rect 47991 39868 48037 39914
rect 48149 39868 48195 39914
rect 48307 39868 48353 39914
rect 48465 39868 48511 39914
rect 54440 40277 54486 40323
rect 54440 40114 54486 40160
rect 54223 39992 54269 40038
rect 54440 39951 54486 39997
rect 54223 39828 54269 39874
rect 54440 39788 54486 39834
rect 45619 39704 45665 39750
rect 45777 39704 45823 39750
rect 45935 39704 45981 39750
rect 46093 39704 46139 39750
rect 46251 39704 46297 39750
rect 46409 39704 46455 39750
rect 46568 39704 46614 39750
rect 46726 39704 46772 39750
rect 46884 39704 46930 39750
rect 47042 39704 47088 39750
rect 47200 39704 47246 39750
rect 47358 39704 47404 39750
rect 47516 39704 47562 39750
rect 47675 39704 47721 39750
rect 47833 39704 47879 39750
rect 47991 39704 48037 39750
rect 48149 39704 48195 39750
rect 48307 39704 48353 39750
rect 48465 39704 48511 39750
rect 45619 39540 45665 39586
rect 45777 39540 45823 39586
rect 45935 39540 45981 39586
rect 46093 39540 46139 39586
rect 46251 39540 46297 39586
rect 46409 39540 46455 39586
rect 46568 39540 46614 39586
rect 46726 39540 46772 39586
rect 46884 39540 46930 39586
rect 47042 39540 47088 39586
rect 47200 39540 47246 39586
rect 47358 39540 47404 39586
rect 47516 39540 47562 39586
rect 47675 39540 47721 39586
rect 47833 39540 47879 39586
rect 47991 39540 48037 39586
rect 48149 39540 48195 39586
rect 48307 39540 48353 39586
rect 48465 39540 48511 39586
rect 54223 39580 54269 39626
rect 54440 39620 54486 39666
rect 30637 38967 30683 39013
rect 30855 38927 30901 38973
rect 54223 39416 54269 39462
rect 54440 39457 54486 39503
rect 54440 39294 54486 39340
rect 54440 39131 54486 39177
rect 54223 38927 54269 38973
rect 54440 38967 54486 39013
rect 30637 38804 30683 38850
rect 54440 38804 54486 38850
rect 30637 38641 30683 38687
rect 30855 38681 30901 38727
rect 30637 38477 30683 38523
rect 30855 38518 30901 38564
rect 30637 38314 30683 38360
rect 30855 38355 30901 38401
rect 30637 38151 30683 38197
rect 30855 38192 30901 38238
rect 30637 37988 30683 38034
rect 30855 38028 30901 38074
rect 54223 38681 54269 38727
rect 54440 38641 54486 38687
rect 36489 37904 36723 37950
rect 30637 37820 30683 37866
rect 30855 37780 30901 37826
rect 30637 37657 30683 37703
rect 30855 37616 30901 37662
rect 30637 37494 30683 37540
rect 30855 37453 30901 37499
rect 30637 37331 30683 37377
rect 30855 37290 30901 37336
rect 39062 37904 39108 37950
rect 39220 37904 39266 37950
rect 45619 38068 45665 38114
rect 45777 38068 45823 38114
rect 45935 38068 45981 38114
rect 46093 38068 46139 38114
rect 46251 38068 46297 38114
rect 46409 38068 46455 38114
rect 46568 38068 46614 38114
rect 46726 38068 46772 38114
rect 46884 38068 46930 38114
rect 47042 38068 47088 38114
rect 47200 38068 47246 38114
rect 47358 38068 47404 38114
rect 47516 38068 47562 38114
rect 47675 38068 47721 38114
rect 47833 38068 47879 38114
rect 47991 38068 48037 38114
rect 48149 38068 48195 38114
rect 48307 38068 48353 38114
rect 48465 38068 48511 38114
rect 54440 38477 54486 38523
rect 54440 38314 54486 38360
rect 54223 38192 54269 38238
rect 54440 38151 54486 38197
rect 54223 38028 54269 38074
rect 54440 37988 54486 38034
rect 45619 37904 45665 37950
rect 45777 37904 45823 37950
rect 45935 37904 45981 37950
rect 46093 37904 46139 37950
rect 46251 37904 46297 37950
rect 46409 37904 46455 37950
rect 46568 37904 46614 37950
rect 46726 37904 46772 37950
rect 46884 37904 46930 37950
rect 47042 37904 47088 37950
rect 47200 37904 47246 37950
rect 47358 37904 47404 37950
rect 47516 37904 47562 37950
rect 47675 37904 47721 37950
rect 47833 37904 47879 37950
rect 47991 37904 48037 37950
rect 48149 37904 48195 37950
rect 48307 37904 48353 37950
rect 48465 37904 48511 37950
rect 45619 37740 45665 37786
rect 45777 37740 45823 37786
rect 45935 37740 45981 37786
rect 46093 37740 46139 37786
rect 46251 37740 46297 37786
rect 46409 37740 46455 37786
rect 46568 37740 46614 37786
rect 46726 37740 46772 37786
rect 46884 37740 46930 37786
rect 47042 37740 47088 37786
rect 47200 37740 47246 37786
rect 47358 37740 47404 37786
rect 47516 37740 47562 37786
rect 47675 37740 47721 37786
rect 47833 37740 47879 37786
rect 47991 37740 48037 37786
rect 48149 37740 48195 37786
rect 48307 37740 48353 37786
rect 48465 37740 48511 37786
rect 54223 37780 54269 37826
rect 54440 37820 54486 37866
rect 30637 37167 30683 37213
rect 30855 37127 30901 37173
rect 54223 37616 54269 37662
rect 54440 37657 54486 37703
rect 54440 37494 54486 37540
rect 54440 37331 54486 37377
rect 54223 37127 54269 37173
rect 54440 37167 54486 37213
rect 30637 37004 30683 37050
rect 54440 37004 54486 37050
rect 30637 36841 30683 36887
rect 30855 36881 30901 36927
rect 30637 36677 30683 36723
rect 30855 36718 30901 36764
rect 30637 36514 30683 36560
rect 30855 36555 30901 36601
rect 30637 36351 30683 36397
rect 30855 36392 30901 36438
rect 30637 36188 30683 36234
rect 30855 36228 30901 36274
rect 54223 36881 54269 36927
rect 54440 36841 54486 36887
rect 36489 36104 36723 36150
rect 39062 36104 39108 36150
rect 39220 36104 39266 36150
rect 45619 36268 45665 36314
rect 45777 36268 45823 36314
rect 45935 36268 45981 36314
rect 46093 36268 46139 36314
rect 46251 36268 46297 36314
rect 46409 36268 46455 36314
rect 46568 36268 46614 36314
rect 46726 36268 46772 36314
rect 46884 36268 46930 36314
rect 47042 36268 47088 36314
rect 47200 36268 47246 36314
rect 47358 36268 47404 36314
rect 47516 36268 47562 36314
rect 47675 36268 47721 36314
rect 47833 36268 47879 36314
rect 47991 36268 48037 36314
rect 48149 36268 48195 36314
rect 48307 36268 48353 36314
rect 48465 36268 48511 36314
rect 54440 36677 54486 36723
rect 54440 36514 54486 36560
rect 54223 36392 54269 36438
rect 54440 36351 54486 36397
rect 54223 36228 54269 36274
rect 54440 36188 54486 36234
rect 45619 36104 45665 36150
rect 45777 36104 45823 36150
rect 45935 36104 45981 36150
rect 46093 36104 46139 36150
rect 46251 36104 46297 36150
rect 46409 36104 46455 36150
rect 46568 36104 46614 36150
rect 46726 36104 46772 36150
rect 46884 36104 46930 36150
rect 47042 36104 47088 36150
rect 47200 36104 47246 36150
rect 47358 36104 47404 36150
rect 47516 36104 47562 36150
rect 47675 36104 47721 36150
rect 47833 36104 47879 36150
rect 47991 36104 48037 36150
rect 48149 36104 48195 36150
rect 48307 36104 48353 36150
rect 48465 36104 48511 36150
<< polysilicon >>
rect 29072 65644 29274 65771
rect 29072 65598 29116 65644
rect 29162 65598 29274 65644
rect 29072 65481 29274 65598
rect 29072 65435 29116 65481
rect 29162 65435 29274 65481
rect 29072 65317 29274 65435
rect 29072 65271 29116 65317
rect 29162 65271 29274 65317
rect 29072 65154 29274 65271
rect 29072 65108 29116 65154
rect 29162 65108 29274 65154
rect 29072 64983 29274 65108
rect 30373 64983 30444 65771
rect 42300 65843 42478 65862
rect 42300 65797 42319 65843
rect 42459 65797 42478 65843
rect 44041 65891 44144 65910
rect 44041 65845 44067 65891
rect 44113 65845 44144 65891
rect 42300 65778 42478 65797
rect 37991 65743 38125 65750
rect 35233 65623 35396 65743
rect 37922 65645 38125 65743
rect 37922 65623 38035 65645
rect 35233 65519 35336 65623
rect 37991 65519 38035 65623
rect 32932 65399 33001 65519
rect 35023 65399 35396 65519
rect 37922 65505 38035 65519
rect 38081 65505 38125 65645
rect 40675 65558 40759 65577
rect 40675 65519 40694 65558
rect 37922 65400 38125 65505
rect 37922 65399 37993 65400
rect 38292 65399 38363 65519
rect 39681 65399 40062 65519
rect 40590 65418 40694 65519
rect 40740 65418 40759 65558
rect 42341 65520 42445 65778
rect 40590 65399 40759 65418
rect 40892 65400 40963 65520
rect 42281 65400 42445 65520
rect 44041 65519 44144 65845
rect 46948 65633 47101 65743
rect 42592 65399 42663 65519
rect 43981 65399 44144 65519
rect 44260 65598 44344 65617
rect 44260 65458 44279 65598
rect 44325 65519 44344 65598
rect 44325 65458 44432 65519
rect 44260 65399 44432 65458
rect 44960 65399 45333 65519
rect 46651 65399 46722 65519
rect 46948 65493 46967 65633
rect 47013 65623 47101 65633
rect 49627 65623 49790 65743
rect 47013 65519 47032 65623
rect 49687 65519 49790 65623
rect 47013 65493 47101 65519
rect 46948 65399 47101 65493
rect 49627 65399 50001 65519
rect 52023 65399 52094 65519
rect 29072 64744 29274 64871
rect 29072 64698 29116 64744
rect 29162 64698 29274 64744
rect 29072 64581 29274 64698
rect 29072 64535 29116 64581
rect 29162 64535 29274 64581
rect 29072 64417 29274 64535
rect 29072 64371 29116 64417
rect 29162 64371 29274 64417
rect 29072 64254 29274 64371
rect 29072 64208 29116 64254
rect 29162 64208 29274 64254
rect 29072 64083 29274 64208
rect 30373 64083 30444 64871
rect 31292 64755 31336 64875
rect 33336 64784 33671 64875
rect 33336 64755 33495 64784
rect 33476 64651 33495 64755
rect 31292 64531 31336 64651
rect 33336 64531 33495 64651
rect 33458 64427 33495 64531
rect 31292 64307 31336 64427
rect 33336 64362 33495 64427
rect 33541 64755 33671 64784
rect 34671 64755 34715 64875
rect 39657 64755 39727 64875
rect 40167 64755 40346 64875
rect 44451 64864 44799 64875
rect 33541 64651 33560 64755
rect 40262 64737 40346 64755
rect 43354 64809 43695 64864
rect 43354 64763 43373 64809
rect 43513 64763 43695 64809
rect 43354 64744 43695 64763
rect 44325 64755 44799 64864
rect 45323 64755 45393 64875
rect 44325 64744 44552 64755
rect 40262 64691 40281 64737
rect 40327 64691 40346 64737
rect 40262 64672 40346 64691
rect 33541 64531 33671 64651
rect 34671 64531 34715 64651
rect 50410 64755 50454 64875
rect 51454 64755 51789 64875
rect 53789 64755 53833 64875
rect 54679 64983 54750 65771
rect 55849 65644 56051 65771
rect 55849 65598 55961 65644
rect 56007 65598 56051 65644
rect 55849 65481 56051 65598
rect 55849 65435 55961 65481
rect 56007 65435 56051 65481
rect 55849 65317 56051 65435
rect 55849 65271 55961 65317
rect 56007 65271 56051 65317
rect 55849 65154 56051 65271
rect 55849 65108 55961 65154
rect 56007 65108 56051 65154
rect 55849 64983 56051 65108
rect 33541 64362 33560 64531
rect 35133 64444 35260 64564
rect 36360 64465 36540 64564
rect 36360 64444 36475 64465
rect 35133 64395 35192 64444
rect 33336 64307 33560 64362
rect 33620 64275 33671 64395
rect 34671 64340 35192 64395
rect 36431 64340 36475 64444
rect 34671 64275 35260 64340
rect 35133 64220 35260 64275
rect 36360 64325 36475 64340
rect 36521 64325 36540 64465
rect 36360 64220 36540 64325
rect 36678 64465 36841 64564
rect 36678 64325 36697 64465
rect 36743 64444 36841 64465
rect 37501 64444 37572 64564
rect 37826 64444 37896 64564
rect 38556 64467 38734 64564
rect 43625 64531 43695 64651
rect 44325 64614 44799 64651
rect 44325 64568 44358 64614
rect 44498 64568 44799 64614
rect 44325 64531 44799 64568
rect 45323 64531 45367 64651
rect 51556 64754 51665 64755
rect 51556 64651 51600 64754
rect 38556 64444 38669 64467
rect 36743 64340 36773 64444
rect 38627 64340 38669 64444
rect 36743 64325 36841 64340
rect 36678 64220 36841 64325
rect 37501 64220 37572 64340
rect 37826 64220 37896 64340
rect 38556 64327 38669 64340
rect 38715 64327 38734 64467
rect 48603 64492 48765 64564
rect 38556 64220 38734 64327
rect 38939 64220 39008 64340
rect 39326 64220 39598 64340
rect 39730 64306 39909 64340
rect 43625 64307 43695 64427
rect 44325 64307 44799 64427
rect 45323 64383 45623 64427
rect 45323 64337 45464 64383
rect 45604 64337 45623 64383
rect 45323 64307 45623 64337
rect 48603 64352 48622 64492
rect 48668 64444 48765 64492
rect 49865 64444 49991 64564
rect 50410 64531 50454 64651
rect 51454 64531 51600 64651
rect 48668 64352 48705 64444
rect 48603 64340 48705 64352
rect 49932 64395 49991 64444
rect 49932 64340 50454 64395
rect 39730 64260 39844 64306
rect 39890 64260 39909 64306
rect 39730 64220 39909 64260
rect 48603 64220 48765 64340
rect 49865 64275 50454 64340
rect 51454 64275 51498 64395
rect 51581 64332 51600 64531
rect 51646 64651 51665 64754
rect 51646 64531 51789 64651
rect 53789 64531 53833 64651
rect 51646 64427 51667 64531
rect 51646 64332 51789 64427
rect 51581 64307 51789 64332
rect 53789 64307 53833 64427
rect 49865 64220 49991 64275
rect 29072 63844 29274 63971
rect 29072 63798 29116 63844
rect 29162 63798 29274 63844
rect 29072 63681 29274 63798
rect 29072 63635 29116 63681
rect 29162 63635 29274 63681
rect 29072 63517 29274 63635
rect 29072 63471 29116 63517
rect 29162 63471 29274 63517
rect 29072 63354 29274 63471
rect 29072 63308 29116 63354
rect 29162 63308 29274 63354
rect 29072 63183 29274 63308
rect 30373 63183 30444 63971
rect 54679 64083 54750 64871
rect 55849 64744 56051 64871
rect 55849 64698 55961 64744
rect 56007 64698 56051 64744
rect 55849 64581 56051 64698
rect 55849 64535 55961 64581
rect 56007 64535 56051 64581
rect 55849 64417 56051 64535
rect 55849 64371 55961 64417
rect 56007 64371 56051 64417
rect 55849 64254 56051 64371
rect 55849 64208 55961 64254
rect 56007 64208 56051 64254
rect 55849 64083 56051 64208
rect 35133 63779 35260 63834
rect 31292 63627 31336 63747
rect 33336 63692 33560 63747
rect 33336 63627 33495 63692
rect 33458 63523 33495 63627
rect 31292 63403 31336 63523
rect 33336 63403 33495 63523
rect 33476 63299 33495 63403
rect 29072 62944 29274 63071
rect 29072 62898 29116 62944
rect 29162 62898 29274 62944
rect 29072 62781 29274 62898
rect 29072 62735 29116 62781
rect 29162 62735 29274 62781
rect 29072 62617 29274 62735
rect 29072 62571 29116 62617
rect 29162 62571 29274 62617
rect 29072 62454 29274 62571
rect 29072 62408 29116 62454
rect 29162 62408 29274 62454
rect 29072 62283 29274 62408
rect 30373 62283 30444 63071
rect 31292 63179 31336 63299
rect 33336 63270 33495 63299
rect 33541 63523 33560 63692
rect 33620 63659 33671 63779
rect 34671 63714 35260 63779
rect 36360 63729 36540 63834
rect 36360 63714 36475 63729
rect 34671 63659 35192 63714
rect 35133 63610 35192 63659
rect 36431 63610 36475 63714
rect 33541 63403 33671 63523
rect 34671 63403 34715 63523
rect 35133 63490 35260 63610
rect 36360 63589 36475 63610
rect 36521 63589 36540 63729
rect 36360 63490 36540 63589
rect 36678 63729 36841 63834
rect 36678 63589 36697 63729
rect 36743 63714 36841 63729
rect 37501 63714 37572 63834
rect 37826 63714 37896 63834
rect 38556 63727 38734 63834
rect 38556 63714 38669 63727
rect 36743 63610 36773 63714
rect 38627 63610 38669 63714
rect 36743 63589 36841 63610
rect 36678 63490 36841 63589
rect 37501 63490 37572 63610
rect 37826 63490 37896 63610
rect 38556 63587 38669 63610
rect 38715 63587 38734 63727
rect 38939 63714 39008 63834
rect 39326 63714 39598 63834
rect 39730 63794 39909 63834
rect 39730 63748 39844 63794
rect 39890 63748 39909 63794
rect 39730 63714 39909 63748
rect 43625 63627 43695 63747
rect 44325 63627 44799 63747
rect 45323 63717 45623 63747
rect 45323 63671 45464 63717
rect 45604 63671 45623 63717
rect 45323 63627 45623 63671
rect 48603 63714 48765 63834
rect 49865 63779 49991 63834
rect 49865 63714 50454 63779
rect 48603 63702 48705 63714
rect 38556 63490 38734 63587
rect 48603 63562 48622 63702
rect 48668 63610 48705 63702
rect 49932 63659 50454 63714
rect 51454 63659 51498 63779
rect 51581 63722 51789 63747
rect 49932 63610 49991 63659
rect 48668 63562 48765 63610
rect 33541 63299 33560 63403
rect 43625 63403 43695 63523
rect 44325 63486 44799 63523
rect 44325 63440 44358 63486
rect 44498 63440 44799 63486
rect 44325 63403 44799 63440
rect 45323 63403 45367 63523
rect 48603 63490 48765 63562
rect 49865 63490 49991 63610
rect 51581 63523 51600 63722
rect 40262 63363 40346 63382
rect 40262 63317 40281 63363
rect 40327 63317 40346 63363
rect 40262 63299 40346 63317
rect 50410 63403 50454 63523
rect 51454 63403 51600 63523
rect 33541 63270 33671 63299
rect 33336 63179 33671 63270
rect 34671 63179 34715 63299
rect 31292 62955 31336 63075
rect 33336 62984 33671 63075
rect 33336 62955 33495 62984
rect 33476 62851 33495 62955
rect 31292 62731 31336 62851
rect 33336 62731 33495 62851
rect 33458 62627 33495 62731
rect 31292 62507 31336 62627
rect 33336 62562 33495 62627
rect 33541 62955 33671 62984
rect 34671 62955 34715 63075
rect 39657 63179 39727 63299
rect 40167 63179 40346 63299
rect 43354 63291 43695 63310
rect 43354 63245 43373 63291
rect 43513 63245 43695 63291
rect 43354 63190 43695 63245
rect 44325 63299 44552 63310
rect 44325 63190 44799 63299
rect 39657 62955 39727 63075
rect 40167 62955 40346 63075
rect 44451 63179 44799 63190
rect 45323 63179 45393 63299
rect 51556 63300 51600 63403
rect 51646 63627 51789 63722
rect 53789 63627 53833 63747
rect 51646 63523 51667 63627
rect 51646 63403 51789 63523
rect 53789 63403 53833 63523
rect 51646 63300 51665 63403
rect 51556 63299 51665 63300
rect 50410 63179 50454 63299
rect 51454 63179 51789 63299
rect 53789 63179 53833 63299
rect 44451 63064 44799 63075
rect 33541 62851 33560 62955
rect 40262 62937 40346 62955
rect 43354 63009 43695 63064
rect 43354 62963 43373 63009
rect 43513 62963 43695 63009
rect 43354 62944 43695 62963
rect 44325 62955 44799 63064
rect 45323 62955 45393 63075
rect 44325 62944 44552 62955
rect 40262 62891 40281 62937
rect 40327 62891 40346 62937
rect 40262 62872 40346 62891
rect 33541 62731 33671 62851
rect 34671 62731 34715 62851
rect 50410 62955 50454 63075
rect 51454 62955 51789 63075
rect 53789 62955 53833 63075
rect 54679 63183 54750 63971
rect 55849 63844 56051 63971
rect 55849 63798 55961 63844
rect 56007 63798 56051 63844
rect 55849 63681 56051 63798
rect 55849 63635 55961 63681
rect 56007 63635 56051 63681
rect 55849 63517 56051 63635
rect 55849 63471 55961 63517
rect 56007 63471 56051 63517
rect 55849 63354 56051 63471
rect 55849 63308 55961 63354
rect 56007 63308 56051 63354
rect 55849 63183 56051 63308
rect 33541 62562 33560 62731
rect 35133 62644 35260 62764
rect 36360 62665 36540 62764
rect 36360 62644 36475 62665
rect 35133 62595 35192 62644
rect 33336 62507 33560 62562
rect 33620 62475 33671 62595
rect 34671 62540 35192 62595
rect 36431 62540 36475 62644
rect 34671 62475 35260 62540
rect 35133 62420 35260 62475
rect 36360 62525 36475 62540
rect 36521 62525 36540 62665
rect 36360 62420 36540 62525
rect 36678 62665 36841 62764
rect 36678 62525 36697 62665
rect 36743 62644 36841 62665
rect 37501 62644 37572 62764
rect 37826 62644 37896 62764
rect 38556 62667 38734 62764
rect 43625 62731 43695 62851
rect 44325 62814 44799 62851
rect 44325 62768 44358 62814
rect 44498 62768 44799 62814
rect 44325 62731 44799 62768
rect 45323 62731 45367 62851
rect 51556 62954 51665 62955
rect 51556 62851 51600 62954
rect 38556 62644 38669 62667
rect 36743 62540 36773 62644
rect 38627 62540 38669 62644
rect 36743 62525 36841 62540
rect 36678 62420 36841 62525
rect 37501 62420 37572 62540
rect 37826 62420 37896 62540
rect 38556 62527 38669 62540
rect 38715 62527 38734 62667
rect 48603 62692 48765 62764
rect 38556 62420 38734 62527
rect 38939 62420 39008 62540
rect 39326 62420 39598 62540
rect 39730 62506 39909 62540
rect 43625 62507 43695 62627
rect 44325 62507 44799 62627
rect 45323 62583 45623 62627
rect 45323 62537 45464 62583
rect 45604 62537 45623 62583
rect 45323 62507 45623 62537
rect 48603 62552 48622 62692
rect 48668 62644 48765 62692
rect 49865 62644 49991 62764
rect 50410 62731 50454 62851
rect 51454 62731 51600 62851
rect 48668 62552 48705 62644
rect 48603 62540 48705 62552
rect 49932 62595 49991 62644
rect 49932 62540 50454 62595
rect 39730 62460 39844 62506
rect 39890 62460 39909 62506
rect 39730 62420 39909 62460
rect 48603 62420 48765 62540
rect 49865 62475 50454 62540
rect 51454 62475 51498 62595
rect 51581 62532 51600 62731
rect 51646 62851 51665 62954
rect 51646 62731 51789 62851
rect 53789 62731 53833 62851
rect 51646 62627 51667 62731
rect 51646 62532 51789 62627
rect 51581 62507 51789 62532
rect 53789 62507 53833 62627
rect 49865 62420 49991 62475
rect 29072 62044 29274 62171
rect 29072 61998 29116 62044
rect 29162 61998 29274 62044
rect 29072 61881 29274 61998
rect 29072 61835 29116 61881
rect 29162 61835 29274 61881
rect 29072 61717 29274 61835
rect 29072 61671 29116 61717
rect 29162 61671 29274 61717
rect 29072 61554 29274 61671
rect 29072 61508 29116 61554
rect 29162 61508 29274 61554
rect 29072 61383 29274 61508
rect 30373 61383 30444 62171
rect 54679 62283 54750 63071
rect 55849 62944 56051 63071
rect 55849 62898 55961 62944
rect 56007 62898 56051 62944
rect 55849 62781 56051 62898
rect 55849 62735 55961 62781
rect 56007 62735 56051 62781
rect 55849 62617 56051 62735
rect 55849 62571 55961 62617
rect 56007 62571 56051 62617
rect 55849 62454 56051 62571
rect 55849 62408 55961 62454
rect 56007 62408 56051 62454
rect 55849 62283 56051 62408
rect 35133 61979 35260 62034
rect 31292 61827 31336 61947
rect 33336 61892 33560 61947
rect 33336 61827 33495 61892
rect 33458 61723 33495 61827
rect 31292 61603 31336 61723
rect 33336 61603 33495 61723
rect 33476 61499 33495 61603
rect 29072 61144 29274 61271
rect 29072 61098 29116 61144
rect 29162 61098 29274 61144
rect 29072 60981 29274 61098
rect 29072 60935 29116 60981
rect 29162 60935 29274 60981
rect 29072 60817 29274 60935
rect 29072 60771 29116 60817
rect 29162 60771 29274 60817
rect 29072 60654 29274 60771
rect 29072 60608 29116 60654
rect 29162 60608 29274 60654
rect 29072 60483 29274 60608
rect 30373 60483 30444 61271
rect 31292 61379 31336 61499
rect 33336 61470 33495 61499
rect 33541 61723 33560 61892
rect 33620 61859 33671 61979
rect 34671 61914 35260 61979
rect 36360 61929 36540 62034
rect 36360 61914 36475 61929
rect 34671 61859 35192 61914
rect 35133 61810 35192 61859
rect 36431 61810 36475 61914
rect 33541 61603 33671 61723
rect 34671 61603 34715 61723
rect 35133 61690 35260 61810
rect 36360 61789 36475 61810
rect 36521 61789 36540 61929
rect 36360 61690 36540 61789
rect 36678 61929 36841 62034
rect 36678 61789 36697 61929
rect 36743 61914 36841 61929
rect 37501 61914 37572 62034
rect 37826 61914 37896 62034
rect 38556 61927 38734 62034
rect 38556 61914 38669 61927
rect 36743 61810 36773 61914
rect 38627 61810 38669 61914
rect 36743 61789 36841 61810
rect 36678 61690 36841 61789
rect 37501 61690 37572 61810
rect 37826 61690 37896 61810
rect 38556 61787 38669 61810
rect 38715 61787 38734 61927
rect 38939 61914 39008 62034
rect 39326 61914 39598 62034
rect 39730 61994 39909 62034
rect 39730 61948 39844 61994
rect 39890 61948 39909 61994
rect 39730 61914 39909 61948
rect 43625 61827 43695 61947
rect 44325 61827 44799 61947
rect 45323 61917 45623 61947
rect 45323 61871 45464 61917
rect 45604 61871 45623 61917
rect 45323 61827 45623 61871
rect 48603 61914 48765 62034
rect 49865 61979 49991 62034
rect 49865 61914 50454 61979
rect 48603 61902 48705 61914
rect 38556 61690 38734 61787
rect 48603 61762 48622 61902
rect 48668 61810 48705 61902
rect 49932 61859 50454 61914
rect 51454 61859 51498 61979
rect 51581 61922 51789 61947
rect 49932 61810 49991 61859
rect 48668 61762 48765 61810
rect 33541 61499 33560 61603
rect 43625 61603 43695 61723
rect 44325 61686 44799 61723
rect 44325 61640 44358 61686
rect 44498 61640 44799 61686
rect 44325 61603 44799 61640
rect 45323 61603 45367 61723
rect 48603 61690 48765 61762
rect 49865 61690 49991 61810
rect 51581 61723 51600 61922
rect 40262 61563 40346 61582
rect 40262 61517 40281 61563
rect 40327 61517 40346 61563
rect 40262 61499 40346 61517
rect 50410 61603 50454 61723
rect 51454 61603 51600 61723
rect 33541 61470 33671 61499
rect 33336 61379 33671 61470
rect 34671 61379 34715 61499
rect 31292 61155 31336 61275
rect 33336 61184 33671 61275
rect 33336 61155 33495 61184
rect 33476 61051 33495 61155
rect 31292 60931 31336 61051
rect 33336 60931 33495 61051
rect 33458 60827 33495 60931
rect 31292 60707 31336 60827
rect 33336 60762 33495 60827
rect 33541 61155 33671 61184
rect 34671 61155 34715 61275
rect 39657 61379 39727 61499
rect 40167 61379 40346 61499
rect 43354 61491 43695 61510
rect 43354 61445 43373 61491
rect 43513 61445 43695 61491
rect 43354 61390 43695 61445
rect 44325 61499 44552 61510
rect 44325 61390 44799 61499
rect 39657 61155 39727 61275
rect 40167 61155 40346 61275
rect 44451 61379 44799 61390
rect 45323 61379 45393 61499
rect 51556 61500 51600 61603
rect 51646 61827 51789 61922
rect 53789 61827 53833 61947
rect 51646 61723 51667 61827
rect 51646 61603 51789 61723
rect 53789 61603 53833 61723
rect 51646 61500 51665 61603
rect 51556 61499 51665 61500
rect 50410 61379 50454 61499
rect 51454 61379 51789 61499
rect 53789 61379 53833 61499
rect 44451 61264 44799 61275
rect 33541 61051 33560 61155
rect 40262 61137 40346 61155
rect 43354 61209 43695 61264
rect 43354 61163 43373 61209
rect 43513 61163 43695 61209
rect 43354 61144 43695 61163
rect 44325 61155 44799 61264
rect 45323 61155 45393 61275
rect 44325 61144 44552 61155
rect 40262 61091 40281 61137
rect 40327 61091 40346 61137
rect 40262 61072 40346 61091
rect 33541 60931 33671 61051
rect 34671 60931 34715 61051
rect 50410 61155 50454 61275
rect 51454 61155 51789 61275
rect 53789 61155 53833 61275
rect 54679 61383 54750 62171
rect 55849 62044 56051 62171
rect 55849 61998 55961 62044
rect 56007 61998 56051 62044
rect 55849 61881 56051 61998
rect 55849 61835 55961 61881
rect 56007 61835 56051 61881
rect 55849 61717 56051 61835
rect 55849 61671 55961 61717
rect 56007 61671 56051 61717
rect 55849 61554 56051 61671
rect 55849 61508 55961 61554
rect 56007 61508 56051 61554
rect 55849 61383 56051 61508
rect 33541 60762 33560 60931
rect 35133 60844 35260 60964
rect 36360 60865 36540 60964
rect 36360 60844 36475 60865
rect 35133 60795 35192 60844
rect 33336 60707 33560 60762
rect 33620 60675 33671 60795
rect 34671 60740 35192 60795
rect 36431 60740 36475 60844
rect 34671 60675 35260 60740
rect 35133 60620 35260 60675
rect 36360 60725 36475 60740
rect 36521 60725 36540 60865
rect 36360 60620 36540 60725
rect 36678 60865 36841 60964
rect 36678 60725 36697 60865
rect 36743 60844 36841 60865
rect 37501 60844 37572 60964
rect 37826 60844 37896 60964
rect 38556 60867 38734 60964
rect 43625 60931 43695 61051
rect 44325 61014 44799 61051
rect 44325 60968 44358 61014
rect 44498 60968 44799 61014
rect 44325 60931 44799 60968
rect 45323 60931 45367 61051
rect 51556 61154 51665 61155
rect 51556 61051 51600 61154
rect 38556 60844 38669 60867
rect 36743 60740 36773 60844
rect 38627 60740 38669 60844
rect 36743 60725 36841 60740
rect 36678 60620 36841 60725
rect 37501 60620 37572 60740
rect 37826 60620 37896 60740
rect 38556 60727 38669 60740
rect 38715 60727 38734 60867
rect 48603 60892 48765 60964
rect 38556 60620 38734 60727
rect 38939 60620 39008 60740
rect 39326 60620 39598 60740
rect 39730 60706 39909 60740
rect 43625 60707 43695 60827
rect 44325 60707 44799 60827
rect 45323 60783 45623 60827
rect 45323 60737 45464 60783
rect 45604 60737 45623 60783
rect 45323 60707 45623 60737
rect 48603 60752 48622 60892
rect 48668 60844 48765 60892
rect 49865 60844 49991 60964
rect 50410 60931 50454 61051
rect 51454 60931 51600 61051
rect 48668 60752 48705 60844
rect 48603 60740 48705 60752
rect 49932 60795 49991 60844
rect 49932 60740 50454 60795
rect 39730 60660 39844 60706
rect 39890 60660 39909 60706
rect 39730 60620 39909 60660
rect 48603 60620 48765 60740
rect 49865 60675 50454 60740
rect 51454 60675 51498 60795
rect 51581 60732 51600 60931
rect 51646 61051 51665 61154
rect 51646 60931 51789 61051
rect 53789 60931 53833 61051
rect 51646 60827 51667 60931
rect 51646 60732 51789 60827
rect 51581 60707 51789 60732
rect 53789 60707 53833 60827
rect 49865 60620 49991 60675
rect 29072 60244 29274 60371
rect 29072 60198 29116 60244
rect 29162 60198 29274 60244
rect 29072 60081 29274 60198
rect 29072 60035 29116 60081
rect 29162 60035 29274 60081
rect 29072 59917 29274 60035
rect 29072 59871 29116 59917
rect 29162 59871 29274 59917
rect 29072 59754 29274 59871
rect 29072 59708 29116 59754
rect 29162 59708 29274 59754
rect 29072 59583 29274 59708
rect 30373 59583 30444 60371
rect 54679 60483 54750 61271
rect 55849 61144 56051 61271
rect 55849 61098 55961 61144
rect 56007 61098 56051 61144
rect 55849 60981 56051 61098
rect 55849 60935 55961 60981
rect 56007 60935 56051 60981
rect 55849 60817 56051 60935
rect 55849 60771 55961 60817
rect 56007 60771 56051 60817
rect 55849 60654 56051 60771
rect 55849 60608 55961 60654
rect 56007 60608 56051 60654
rect 55849 60483 56051 60608
rect 35133 60179 35260 60234
rect 31292 60027 31336 60147
rect 33336 60092 33560 60147
rect 33336 60027 33495 60092
rect 33458 59923 33495 60027
rect 31292 59803 31336 59923
rect 33336 59803 33495 59923
rect 33476 59699 33495 59803
rect 29072 59344 29274 59471
rect 29072 59298 29116 59344
rect 29162 59298 29274 59344
rect 29072 59181 29274 59298
rect 29072 59135 29116 59181
rect 29162 59135 29274 59181
rect 29072 59017 29274 59135
rect 29072 58971 29116 59017
rect 29162 58971 29274 59017
rect 29072 58854 29274 58971
rect 29072 58808 29116 58854
rect 29162 58808 29274 58854
rect 29072 58683 29274 58808
rect 30373 58683 30444 59471
rect 31292 59579 31336 59699
rect 33336 59670 33495 59699
rect 33541 59923 33560 60092
rect 33620 60059 33671 60179
rect 34671 60114 35260 60179
rect 36360 60129 36540 60234
rect 36360 60114 36475 60129
rect 34671 60059 35192 60114
rect 35133 60010 35192 60059
rect 36431 60010 36475 60114
rect 33541 59803 33671 59923
rect 34671 59803 34715 59923
rect 35133 59890 35260 60010
rect 36360 59989 36475 60010
rect 36521 59989 36540 60129
rect 36360 59890 36540 59989
rect 36678 60129 36841 60234
rect 36678 59989 36697 60129
rect 36743 60114 36841 60129
rect 37501 60114 37572 60234
rect 37826 60114 37896 60234
rect 38556 60127 38734 60234
rect 38556 60114 38669 60127
rect 36743 60010 36773 60114
rect 38627 60010 38669 60114
rect 36743 59989 36841 60010
rect 36678 59890 36841 59989
rect 37501 59890 37572 60010
rect 37826 59890 37896 60010
rect 38556 59987 38669 60010
rect 38715 59987 38734 60127
rect 38939 60114 39008 60234
rect 39326 60114 39598 60234
rect 39730 60194 39909 60234
rect 39730 60148 39844 60194
rect 39890 60148 39909 60194
rect 39730 60114 39909 60148
rect 43625 60027 43695 60147
rect 44325 60027 44799 60147
rect 45323 60117 45623 60147
rect 45323 60071 45464 60117
rect 45604 60071 45623 60117
rect 45323 60027 45623 60071
rect 48603 60114 48765 60234
rect 49865 60179 49991 60234
rect 49865 60114 50454 60179
rect 48603 60102 48705 60114
rect 38556 59890 38734 59987
rect 48603 59962 48622 60102
rect 48668 60010 48705 60102
rect 49932 60059 50454 60114
rect 51454 60059 51498 60179
rect 51581 60122 51789 60147
rect 49932 60010 49991 60059
rect 48668 59962 48765 60010
rect 33541 59699 33560 59803
rect 43625 59803 43695 59923
rect 44325 59886 44799 59923
rect 44325 59840 44358 59886
rect 44498 59840 44799 59886
rect 44325 59803 44799 59840
rect 45323 59803 45367 59923
rect 48603 59890 48765 59962
rect 49865 59890 49991 60010
rect 51581 59923 51600 60122
rect 40262 59763 40346 59782
rect 40262 59717 40281 59763
rect 40327 59717 40346 59763
rect 40262 59699 40346 59717
rect 50410 59803 50454 59923
rect 51454 59803 51600 59923
rect 33541 59670 33671 59699
rect 33336 59579 33671 59670
rect 34671 59579 34715 59699
rect 31292 59355 31336 59475
rect 33336 59384 33671 59475
rect 33336 59355 33495 59384
rect 33476 59251 33495 59355
rect 31292 59131 31336 59251
rect 33336 59131 33495 59251
rect 33458 59027 33495 59131
rect 31292 58907 31336 59027
rect 33336 58962 33495 59027
rect 33541 59355 33671 59384
rect 34671 59355 34715 59475
rect 39657 59579 39727 59699
rect 40167 59579 40346 59699
rect 43354 59691 43695 59710
rect 43354 59645 43373 59691
rect 43513 59645 43695 59691
rect 43354 59590 43695 59645
rect 44325 59699 44552 59710
rect 44325 59590 44799 59699
rect 39657 59355 39727 59475
rect 40167 59355 40346 59475
rect 44451 59579 44799 59590
rect 45323 59579 45393 59699
rect 51556 59700 51600 59803
rect 51646 60027 51789 60122
rect 53789 60027 53833 60147
rect 51646 59923 51667 60027
rect 51646 59803 51789 59923
rect 53789 59803 53833 59923
rect 51646 59700 51665 59803
rect 51556 59699 51665 59700
rect 50410 59579 50454 59699
rect 51454 59579 51789 59699
rect 53789 59579 53833 59699
rect 44451 59464 44799 59475
rect 33541 59251 33560 59355
rect 40262 59337 40346 59355
rect 43354 59409 43695 59464
rect 43354 59363 43373 59409
rect 43513 59363 43695 59409
rect 43354 59344 43695 59363
rect 44325 59355 44799 59464
rect 45323 59355 45393 59475
rect 44325 59344 44552 59355
rect 40262 59291 40281 59337
rect 40327 59291 40346 59337
rect 40262 59272 40346 59291
rect 33541 59131 33671 59251
rect 34671 59131 34715 59251
rect 50410 59355 50454 59475
rect 51454 59355 51789 59475
rect 53789 59355 53833 59475
rect 54679 59583 54750 60371
rect 55849 60244 56051 60371
rect 55849 60198 55961 60244
rect 56007 60198 56051 60244
rect 55849 60081 56051 60198
rect 55849 60035 55961 60081
rect 56007 60035 56051 60081
rect 55849 59917 56051 60035
rect 55849 59871 55961 59917
rect 56007 59871 56051 59917
rect 55849 59754 56051 59871
rect 55849 59708 55961 59754
rect 56007 59708 56051 59754
rect 55849 59583 56051 59708
rect 33541 58962 33560 59131
rect 35133 59044 35260 59164
rect 36360 59065 36540 59164
rect 36360 59044 36475 59065
rect 35133 58995 35192 59044
rect 33336 58907 33560 58962
rect 33620 58875 33671 58995
rect 34671 58940 35192 58995
rect 36431 58940 36475 59044
rect 34671 58875 35260 58940
rect 35133 58820 35260 58875
rect 36360 58925 36475 58940
rect 36521 58925 36540 59065
rect 36360 58820 36540 58925
rect 36678 59065 36841 59164
rect 36678 58925 36697 59065
rect 36743 59044 36841 59065
rect 37501 59044 37572 59164
rect 37826 59044 37896 59164
rect 38556 59067 38734 59164
rect 43625 59131 43695 59251
rect 44325 59214 44799 59251
rect 44325 59168 44358 59214
rect 44498 59168 44799 59214
rect 44325 59131 44799 59168
rect 45323 59131 45367 59251
rect 51556 59354 51665 59355
rect 51556 59251 51600 59354
rect 38556 59044 38669 59067
rect 36743 58940 36773 59044
rect 38627 58940 38669 59044
rect 36743 58925 36841 58940
rect 36678 58820 36841 58925
rect 37501 58820 37572 58940
rect 37826 58820 37896 58940
rect 38556 58927 38669 58940
rect 38715 58927 38734 59067
rect 48603 59092 48765 59164
rect 38556 58820 38734 58927
rect 38939 58820 39008 58940
rect 39326 58820 39598 58940
rect 39730 58906 39909 58940
rect 43625 58907 43695 59027
rect 44325 58907 44799 59027
rect 45323 58983 45623 59027
rect 45323 58937 45464 58983
rect 45604 58937 45623 58983
rect 45323 58907 45623 58937
rect 48603 58952 48622 59092
rect 48668 59044 48765 59092
rect 49865 59044 49991 59164
rect 50410 59131 50454 59251
rect 51454 59131 51600 59251
rect 48668 58952 48705 59044
rect 48603 58940 48705 58952
rect 49932 58995 49991 59044
rect 49932 58940 50454 58995
rect 39730 58860 39844 58906
rect 39890 58860 39909 58906
rect 39730 58820 39909 58860
rect 48603 58820 48765 58940
rect 49865 58875 50454 58940
rect 51454 58875 51498 58995
rect 51581 58932 51600 59131
rect 51646 59251 51665 59354
rect 51646 59131 51789 59251
rect 53789 59131 53833 59251
rect 51646 59027 51667 59131
rect 51646 58932 51789 59027
rect 51581 58907 51789 58932
rect 53789 58907 53833 59027
rect 49865 58820 49991 58875
rect 29072 58444 29274 58571
rect 29072 58398 29116 58444
rect 29162 58398 29274 58444
rect 29072 58281 29274 58398
rect 29072 58235 29116 58281
rect 29162 58235 29274 58281
rect 29072 58117 29274 58235
rect 29072 58071 29116 58117
rect 29162 58071 29274 58117
rect 29072 57954 29274 58071
rect 29072 57908 29116 57954
rect 29162 57908 29274 57954
rect 29072 57783 29274 57908
rect 30373 57783 30444 58571
rect 54679 58683 54750 59471
rect 55849 59344 56051 59471
rect 55849 59298 55961 59344
rect 56007 59298 56051 59344
rect 55849 59181 56051 59298
rect 55849 59135 55961 59181
rect 56007 59135 56051 59181
rect 55849 59017 56051 59135
rect 55849 58971 55961 59017
rect 56007 58971 56051 59017
rect 55849 58854 56051 58971
rect 55849 58808 55961 58854
rect 56007 58808 56051 58854
rect 55849 58683 56051 58808
rect 35133 58379 35260 58434
rect 31292 58227 31336 58347
rect 33336 58292 33560 58347
rect 33336 58227 33495 58292
rect 33458 58123 33495 58227
rect 31292 58003 31336 58123
rect 33336 58003 33495 58123
rect 33476 57899 33495 58003
rect 29072 57544 29274 57671
rect 29072 57498 29116 57544
rect 29162 57498 29274 57544
rect 29072 57381 29274 57498
rect 29072 57335 29116 57381
rect 29162 57335 29274 57381
rect 29072 57217 29274 57335
rect 29072 57171 29116 57217
rect 29162 57171 29274 57217
rect 29072 57054 29274 57171
rect 29072 57008 29116 57054
rect 29162 57008 29274 57054
rect 29072 56883 29274 57008
rect 30373 56883 30444 57671
rect 31292 57779 31336 57899
rect 33336 57870 33495 57899
rect 33541 58123 33560 58292
rect 33620 58259 33671 58379
rect 34671 58314 35260 58379
rect 36360 58329 36540 58434
rect 36360 58314 36475 58329
rect 34671 58259 35192 58314
rect 35133 58210 35192 58259
rect 36431 58210 36475 58314
rect 33541 58003 33671 58123
rect 34671 58003 34715 58123
rect 35133 58090 35260 58210
rect 36360 58189 36475 58210
rect 36521 58189 36540 58329
rect 36360 58090 36540 58189
rect 36678 58329 36841 58434
rect 36678 58189 36697 58329
rect 36743 58314 36841 58329
rect 37501 58314 37572 58434
rect 37826 58314 37896 58434
rect 38556 58327 38734 58434
rect 38556 58314 38669 58327
rect 36743 58210 36773 58314
rect 38627 58210 38669 58314
rect 36743 58189 36841 58210
rect 36678 58090 36841 58189
rect 37501 58090 37572 58210
rect 37826 58090 37896 58210
rect 38556 58187 38669 58210
rect 38715 58187 38734 58327
rect 38939 58314 39008 58434
rect 39326 58314 39598 58434
rect 39730 58394 39909 58434
rect 39730 58348 39844 58394
rect 39890 58348 39909 58394
rect 39730 58314 39909 58348
rect 43625 58227 43695 58347
rect 44325 58227 44799 58347
rect 45323 58317 45623 58347
rect 45323 58271 45464 58317
rect 45604 58271 45623 58317
rect 45323 58227 45623 58271
rect 48603 58314 48765 58434
rect 49865 58379 49991 58434
rect 49865 58314 50454 58379
rect 48603 58302 48705 58314
rect 38556 58090 38734 58187
rect 48603 58162 48622 58302
rect 48668 58210 48705 58302
rect 49932 58259 50454 58314
rect 51454 58259 51498 58379
rect 51581 58322 51789 58347
rect 49932 58210 49991 58259
rect 48668 58162 48765 58210
rect 33541 57899 33560 58003
rect 43625 58003 43695 58123
rect 44325 58086 44799 58123
rect 44325 58040 44358 58086
rect 44498 58040 44799 58086
rect 44325 58003 44799 58040
rect 45323 58003 45367 58123
rect 48603 58090 48765 58162
rect 49865 58090 49991 58210
rect 51581 58123 51600 58322
rect 40262 57963 40346 57982
rect 40262 57917 40281 57963
rect 40327 57917 40346 57963
rect 40262 57899 40346 57917
rect 50410 58003 50454 58123
rect 51454 58003 51600 58123
rect 33541 57870 33671 57899
rect 33336 57779 33671 57870
rect 34671 57779 34715 57899
rect 31292 57555 31336 57675
rect 33336 57584 33671 57675
rect 33336 57555 33495 57584
rect 33476 57451 33495 57555
rect 31292 57331 31336 57451
rect 33336 57331 33495 57451
rect 33458 57227 33495 57331
rect 31292 57107 31336 57227
rect 33336 57162 33495 57227
rect 33541 57555 33671 57584
rect 34671 57555 34715 57675
rect 39657 57779 39727 57899
rect 40167 57779 40346 57899
rect 43354 57891 43695 57910
rect 43354 57845 43373 57891
rect 43513 57845 43695 57891
rect 43354 57790 43695 57845
rect 44325 57899 44552 57910
rect 44325 57790 44799 57899
rect 39657 57555 39727 57675
rect 40167 57555 40346 57675
rect 44451 57779 44799 57790
rect 45323 57779 45393 57899
rect 51556 57900 51600 58003
rect 51646 58227 51789 58322
rect 53789 58227 53833 58347
rect 51646 58123 51667 58227
rect 51646 58003 51789 58123
rect 53789 58003 53833 58123
rect 51646 57900 51665 58003
rect 51556 57899 51665 57900
rect 50410 57779 50454 57899
rect 51454 57779 51789 57899
rect 53789 57779 53833 57899
rect 44451 57664 44799 57675
rect 33541 57451 33560 57555
rect 40262 57537 40346 57555
rect 43354 57609 43695 57664
rect 43354 57563 43373 57609
rect 43513 57563 43695 57609
rect 43354 57544 43695 57563
rect 44325 57555 44799 57664
rect 45323 57555 45393 57675
rect 44325 57544 44552 57555
rect 40262 57491 40281 57537
rect 40327 57491 40346 57537
rect 40262 57472 40346 57491
rect 33541 57331 33671 57451
rect 34671 57331 34715 57451
rect 50410 57555 50454 57675
rect 51454 57555 51789 57675
rect 53789 57555 53833 57675
rect 54679 57783 54750 58571
rect 55849 58444 56051 58571
rect 55849 58398 55961 58444
rect 56007 58398 56051 58444
rect 55849 58281 56051 58398
rect 55849 58235 55961 58281
rect 56007 58235 56051 58281
rect 55849 58117 56051 58235
rect 55849 58071 55961 58117
rect 56007 58071 56051 58117
rect 55849 57954 56051 58071
rect 55849 57908 55961 57954
rect 56007 57908 56051 57954
rect 55849 57783 56051 57908
rect 33541 57162 33560 57331
rect 35133 57244 35260 57364
rect 36360 57265 36540 57364
rect 36360 57244 36475 57265
rect 35133 57195 35192 57244
rect 33336 57107 33560 57162
rect 33620 57075 33671 57195
rect 34671 57140 35192 57195
rect 36431 57140 36475 57244
rect 34671 57075 35260 57140
rect 35133 57020 35260 57075
rect 36360 57125 36475 57140
rect 36521 57125 36540 57265
rect 36360 57020 36540 57125
rect 36678 57265 36841 57364
rect 36678 57125 36697 57265
rect 36743 57244 36841 57265
rect 37501 57244 37572 57364
rect 37826 57244 37896 57364
rect 38556 57267 38734 57364
rect 43625 57331 43695 57451
rect 44325 57414 44799 57451
rect 44325 57368 44358 57414
rect 44498 57368 44799 57414
rect 44325 57331 44799 57368
rect 45323 57331 45367 57451
rect 51556 57554 51665 57555
rect 51556 57451 51600 57554
rect 38556 57244 38669 57267
rect 36743 57140 36773 57244
rect 38627 57140 38669 57244
rect 36743 57125 36841 57140
rect 36678 57020 36841 57125
rect 37501 57020 37572 57140
rect 37826 57020 37896 57140
rect 38556 57127 38669 57140
rect 38715 57127 38734 57267
rect 48603 57292 48765 57364
rect 38556 57020 38734 57127
rect 38939 57020 39008 57140
rect 39326 57020 39598 57140
rect 39730 57106 39909 57140
rect 43625 57107 43695 57227
rect 44325 57107 44799 57227
rect 45323 57183 45623 57227
rect 45323 57137 45464 57183
rect 45604 57137 45623 57183
rect 45323 57107 45623 57137
rect 48603 57152 48622 57292
rect 48668 57244 48765 57292
rect 49865 57244 49991 57364
rect 50410 57331 50454 57451
rect 51454 57331 51600 57451
rect 48668 57152 48705 57244
rect 48603 57140 48705 57152
rect 49932 57195 49991 57244
rect 49932 57140 50454 57195
rect 39730 57060 39844 57106
rect 39890 57060 39909 57106
rect 39730 57020 39909 57060
rect 48603 57020 48765 57140
rect 49865 57075 50454 57140
rect 51454 57075 51498 57195
rect 51581 57132 51600 57331
rect 51646 57451 51665 57554
rect 51646 57331 51789 57451
rect 53789 57331 53833 57451
rect 51646 57227 51667 57331
rect 51646 57132 51789 57227
rect 51581 57107 51789 57132
rect 53789 57107 53833 57227
rect 49865 57020 49991 57075
rect 29072 56644 29274 56771
rect 29072 56598 29116 56644
rect 29162 56598 29274 56644
rect 29072 56481 29274 56598
rect 29072 56435 29116 56481
rect 29162 56435 29274 56481
rect 29072 56317 29274 56435
rect 29072 56271 29116 56317
rect 29162 56271 29274 56317
rect 29072 56154 29274 56271
rect 29072 56108 29116 56154
rect 29162 56108 29274 56154
rect 29072 55983 29274 56108
rect 30373 55983 30444 56771
rect 54679 56883 54750 57671
rect 55849 57544 56051 57671
rect 55849 57498 55961 57544
rect 56007 57498 56051 57544
rect 55849 57381 56051 57498
rect 55849 57335 55961 57381
rect 56007 57335 56051 57381
rect 55849 57217 56051 57335
rect 55849 57171 55961 57217
rect 56007 57171 56051 57217
rect 55849 57054 56051 57171
rect 55849 57008 55961 57054
rect 56007 57008 56051 57054
rect 55849 56883 56051 57008
rect 35133 56579 35260 56634
rect 31292 56427 31336 56547
rect 33336 56492 33560 56547
rect 33336 56427 33495 56492
rect 33458 56323 33495 56427
rect 31292 56203 31336 56323
rect 33336 56203 33495 56323
rect 33476 56099 33495 56203
rect 29072 55744 29274 55871
rect 29072 55698 29116 55744
rect 29162 55698 29274 55744
rect 29072 55581 29274 55698
rect 29072 55535 29116 55581
rect 29162 55535 29274 55581
rect 29072 55417 29274 55535
rect 29072 55371 29116 55417
rect 29162 55371 29274 55417
rect 29072 55254 29274 55371
rect 29072 55208 29116 55254
rect 29162 55208 29274 55254
rect 29072 55083 29274 55208
rect 30373 55083 30444 55871
rect 31292 55979 31336 56099
rect 33336 56070 33495 56099
rect 33541 56323 33560 56492
rect 33620 56459 33671 56579
rect 34671 56514 35260 56579
rect 36360 56529 36540 56634
rect 36360 56514 36475 56529
rect 34671 56459 35192 56514
rect 35133 56410 35192 56459
rect 36431 56410 36475 56514
rect 33541 56203 33671 56323
rect 34671 56203 34715 56323
rect 35133 56290 35260 56410
rect 36360 56389 36475 56410
rect 36521 56389 36540 56529
rect 36360 56290 36540 56389
rect 36678 56529 36841 56634
rect 36678 56389 36697 56529
rect 36743 56514 36841 56529
rect 37501 56514 37572 56634
rect 37826 56514 37896 56634
rect 38556 56527 38734 56634
rect 38556 56514 38669 56527
rect 36743 56410 36773 56514
rect 38627 56410 38669 56514
rect 36743 56389 36841 56410
rect 36678 56290 36841 56389
rect 37501 56290 37572 56410
rect 37826 56290 37896 56410
rect 38556 56387 38669 56410
rect 38715 56387 38734 56527
rect 38939 56514 39008 56634
rect 39326 56514 39598 56634
rect 39730 56594 39909 56634
rect 39730 56548 39844 56594
rect 39890 56548 39909 56594
rect 39730 56514 39909 56548
rect 43625 56427 43695 56547
rect 44325 56427 44799 56547
rect 45323 56517 45623 56547
rect 45323 56471 45464 56517
rect 45604 56471 45623 56517
rect 45323 56427 45623 56471
rect 48603 56514 48765 56634
rect 49865 56579 49991 56634
rect 49865 56514 50454 56579
rect 48603 56502 48705 56514
rect 38556 56290 38734 56387
rect 48603 56362 48622 56502
rect 48668 56410 48705 56502
rect 49932 56459 50454 56514
rect 51454 56459 51498 56579
rect 51581 56522 51789 56547
rect 49932 56410 49991 56459
rect 48668 56362 48765 56410
rect 33541 56099 33560 56203
rect 43625 56203 43695 56323
rect 44325 56286 44799 56323
rect 44325 56240 44358 56286
rect 44498 56240 44799 56286
rect 44325 56203 44799 56240
rect 45323 56203 45367 56323
rect 48603 56290 48765 56362
rect 49865 56290 49991 56410
rect 51581 56323 51600 56522
rect 40262 56163 40346 56182
rect 40262 56117 40281 56163
rect 40327 56117 40346 56163
rect 40262 56099 40346 56117
rect 50410 56203 50454 56323
rect 51454 56203 51600 56323
rect 33541 56070 33671 56099
rect 33336 55979 33671 56070
rect 34671 55979 34715 56099
rect 31292 55755 31336 55875
rect 33336 55784 33671 55875
rect 33336 55755 33495 55784
rect 33476 55651 33495 55755
rect 31292 55531 31336 55651
rect 33336 55531 33495 55651
rect 33458 55427 33495 55531
rect 31292 55307 31336 55427
rect 33336 55362 33495 55427
rect 33541 55755 33671 55784
rect 34671 55755 34715 55875
rect 39657 55979 39727 56099
rect 40167 55979 40346 56099
rect 43354 56091 43695 56110
rect 43354 56045 43373 56091
rect 43513 56045 43695 56091
rect 43354 55990 43695 56045
rect 44325 56099 44552 56110
rect 44325 55990 44799 56099
rect 39657 55755 39727 55875
rect 40167 55755 40346 55875
rect 44451 55979 44799 55990
rect 45323 55979 45393 56099
rect 51556 56100 51600 56203
rect 51646 56427 51789 56522
rect 53789 56427 53833 56547
rect 51646 56323 51667 56427
rect 51646 56203 51789 56323
rect 53789 56203 53833 56323
rect 51646 56100 51665 56203
rect 51556 56099 51665 56100
rect 50410 55979 50454 56099
rect 51454 55979 51789 56099
rect 53789 55979 53833 56099
rect 44451 55864 44799 55875
rect 33541 55651 33560 55755
rect 40262 55737 40346 55755
rect 43354 55809 43695 55864
rect 43354 55763 43373 55809
rect 43513 55763 43695 55809
rect 43354 55744 43695 55763
rect 44325 55755 44799 55864
rect 45323 55755 45393 55875
rect 44325 55744 44552 55755
rect 40262 55691 40281 55737
rect 40327 55691 40346 55737
rect 40262 55672 40346 55691
rect 33541 55531 33671 55651
rect 34671 55531 34715 55651
rect 50410 55755 50454 55875
rect 51454 55755 51789 55875
rect 53789 55755 53833 55875
rect 54679 55983 54750 56771
rect 55849 56644 56051 56771
rect 55849 56598 55961 56644
rect 56007 56598 56051 56644
rect 55849 56481 56051 56598
rect 55849 56435 55961 56481
rect 56007 56435 56051 56481
rect 55849 56317 56051 56435
rect 55849 56271 55961 56317
rect 56007 56271 56051 56317
rect 55849 56154 56051 56271
rect 55849 56108 55961 56154
rect 56007 56108 56051 56154
rect 55849 55983 56051 56108
rect 33541 55362 33560 55531
rect 35133 55444 35260 55564
rect 36360 55465 36540 55564
rect 36360 55444 36475 55465
rect 35133 55395 35192 55444
rect 33336 55307 33560 55362
rect 33620 55275 33671 55395
rect 34671 55340 35192 55395
rect 36431 55340 36475 55444
rect 34671 55275 35260 55340
rect 35133 55220 35260 55275
rect 36360 55325 36475 55340
rect 36521 55325 36540 55465
rect 36360 55220 36540 55325
rect 36678 55465 36841 55564
rect 36678 55325 36697 55465
rect 36743 55444 36841 55465
rect 37501 55444 37572 55564
rect 37826 55444 37896 55564
rect 38556 55467 38734 55564
rect 43625 55531 43695 55651
rect 44325 55614 44799 55651
rect 44325 55568 44358 55614
rect 44498 55568 44799 55614
rect 44325 55531 44799 55568
rect 45323 55531 45367 55651
rect 51556 55754 51665 55755
rect 51556 55651 51600 55754
rect 38556 55444 38669 55467
rect 36743 55340 36773 55444
rect 38627 55340 38669 55444
rect 36743 55325 36841 55340
rect 36678 55220 36841 55325
rect 37501 55220 37572 55340
rect 37826 55220 37896 55340
rect 38556 55327 38669 55340
rect 38715 55327 38734 55467
rect 48603 55492 48765 55564
rect 38556 55220 38734 55327
rect 38939 55220 39008 55340
rect 39326 55220 39598 55340
rect 39730 55306 39909 55340
rect 43625 55307 43695 55427
rect 44325 55307 44799 55427
rect 45323 55383 45623 55427
rect 45323 55337 45464 55383
rect 45604 55337 45623 55383
rect 45323 55307 45623 55337
rect 48603 55352 48622 55492
rect 48668 55444 48765 55492
rect 49865 55444 49991 55564
rect 50410 55531 50454 55651
rect 51454 55531 51600 55651
rect 48668 55352 48705 55444
rect 48603 55340 48705 55352
rect 49932 55395 49991 55444
rect 49932 55340 50454 55395
rect 39730 55260 39844 55306
rect 39890 55260 39909 55306
rect 39730 55220 39909 55260
rect 48603 55220 48765 55340
rect 49865 55275 50454 55340
rect 51454 55275 51498 55395
rect 51581 55332 51600 55531
rect 51646 55651 51665 55754
rect 51646 55531 51789 55651
rect 53789 55531 53833 55651
rect 51646 55427 51667 55531
rect 51646 55332 51789 55427
rect 51581 55307 51789 55332
rect 53789 55307 53833 55427
rect 49865 55220 49991 55275
rect 29072 54844 29274 54971
rect 29072 54798 29116 54844
rect 29162 54798 29274 54844
rect 29072 54681 29274 54798
rect 29072 54635 29116 54681
rect 29162 54635 29274 54681
rect 29072 54517 29274 54635
rect 29072 54471 29116 54517
rect 29162 54471 29274 54517
rect 29072 54354 29274 54471
rect 29072 54308 29116 54354
rect 29162 54308 29274 54354
rect 29072 54183 29274 54308
rect 30373 54183 30444 54971
rect 54679 55083 54750 55871
rect 55849 55744 56051 55871
rect 55849 55698 55961 55744
rect 56007 55698 56051 55744
rect 55849 55581 56051 55698
rect 55849 55535 55961 55581
rect 56007 55535 56051 55581
rect 55849 55417 56051 55535
rect 55849 55371 55961 55417
rect 56007 55371 56051 55417
rect 55849 55254 56051 55371
rect 55849 55208 55961 55254
rect 56007 55208 56051 55254
rect 55849 55083 56051 55208
rect 35133 54779 35260 54834
rect 31292 54627 31336 54747
rect 33336 54692 33560 54747
rect 33336 54627 33495 54692
rect 33458 54523 33495 54627
rect 31292 54403 31336 54523
rect 33336 54403 33495 54523
rect 33476 54299 33495 54403
rect 29072 53944 29274 54071
rect 29072 53898 29116 53944
rect 29162 53898 29274 53944
rect 29072 53781 29274 53898
rect 29072 53735 29116 53781
rect 29162 53735 29274 53781
rect 29072 53617 29274 53735
rect 29072 53571 29116 53617
rect 29162 53571 29274 53617
rect 29072 53454 29274 53571
rect 29072 53408 29116 53454
rect 29162 53408 29274 53454
rect 29072 53283 29274 53408
rect 30373 53283 30444 54071
rect 31292 54179 31336 54299
rect 33336 54270 33495 54299
rect 33541 54523 33560 54692
rect 33620 54659 33671 54779
rect 34671 54714 35260 54779
rect 36360 54729 36540 54834
rect 36360 54714 36475 54729
rect 34671 54659 35192 54714
rect 35133 54610 35192 54659
rect 36431 54610 36475 54714
rect 33541 54403 33671 54523
rect 34671 54403 34715 54523
rect 35133 54490 35260 54610
rect 36360 54589 36475 54610
rect 36521 54589 36540 54729
rect 36360 54490 36540 54589
rect 36678 54729 36841 54834
rect 36678 54589 36697 54729
rect 36743 54714 36841 54729
rect 37501 54714 37572 54834
rect 37826 54714 37896 54834
rect 38556 54727 38734 54834
rect 38556 54714 38669 54727
rect 36743 54610 36773 54714
rect 38627 54610 38669 54714
rect 36743 54589 36841 54610
rect 36678 54490 36841 54589
rect 37501 54490 37572 54610
rect 37826 54490 37896 54610
rect 38556 54587 38669 54610
rect 38715 54587 38734 54727
rect 38939 54714 39008 54834
rect 39326 54714 39598 54834
rect 39730 54794 39909 54834
rect 39730 54748 39844 54794
rect 39890 54748 39909 54794
rect 39730 54714 39909 54748
rect 43625 54627 43695 54747
rect 44325 54627 44799 54747
rect 45323 54717 45623 54747
rect 45323 54671 45464 54717
rect 45604 54671 45623 54717
rect 45323 54627 45623 54671
rect 48603 54714 48765 54834
rect 49865 54779 49991 54834
rect 49865 54714 50454 54779
rect 48603 54702 48705 54714
rect 38556 54490 38734 54587
rect 48603 54562 48622 54702
rect 48668 54610 48705 54702
rect 49932 54659 50454 54714
rect 51454 54659 51498 54779
rect 51581 54722 51789 54747
rect 49932 54610 49991 54659
rect 48668 54562 48765 54610
rect 33541 54299 33560 54403
rect 43625 54403 43695 54523
rect 44325 54486 44799 54523
rect 44325 54440 44358 54486
rect 44498 54440 44799 54486
rect 44325 54403 44799 54440
rect 45323 54403 45367 54523
rect 48603 54490 48765 54562
rect 49865 54490 49991 54610
rect 51581 54523 51600 54722
rect 40262 54363 40346 54382
rect 40262 54317 40281 54363
rect 40327 54317 40346 54363
rect 40262 54299 40346 54317
rect 50410 54403 50454 54523
rect 51454 54403 51600 54523
rect 33541 54270 33671 54299
rect 33336 54179 33671 54270
rect 34671 54179 34715 54299
rect 31292 53955 31336 54075
rect 33336 53984 33671 54075
rect 33336 53955 33495 53984
rect 33476 53851 33495 53955
rect 31292 53731 31336 53851
rect 33336 53731 33495 53851
rect 33458 53627 33495 53731
rect 31292 53507 31336 53627
rect 33336 53562 33495 53627
rect 33541 53955 33671 53984
rect 34671 53955 34715 54075
rect 39657 54179 39727 54299
rect 40167 54179 40346 54299
rect 43354 54291 43695 54310
rect 43354 54245 43373 54291
rect 43513 54245 43695 54291
rect 43354 54190 43695 54245
rect 44325 54299 44552 54310
rect 44325 54190 44799 54299
rect 39657 53955 39727 54075
rect 40167 53955 40346 54075
rect 44451 54179 44799 54190
rect 45323 54179 45393 54299
rect 51556 54300 51600 54403
rect 51646 54627 51789 54722
rect 53789 54627 53833 54747
rect 51646 54523 51667 54627
rect 51646 54403 51789 54523
rect 53789 54403 53833 54523
rect 51646 54300 51665 54403
rect 51556 54299 51665 54300
rect 50410 54179 50454 54299
rect 51454 54179 51789 54299
rect 53789 54179 53833 54299
rect 44451 54064 44799 54075
rect 33541 53851 33560 53955
rect 40262 53937 40346 53955
rect 43354 54009 43695 54064
rect 43354 53963 43373 54009
rect 43513 53963 43695 54009
rect 43354 53944 43695 53963
rect 44325 53955 44799 54064
rect 45323 53955 45393 54075
rect 44325 53944 44552 53955
rect 40262 53891 40281 53937
rect 40327 53891 40346 53937
rect 40262 53872 40346 53891
rect 33541 53731 33671 53851
rect 34671 53731 34715 53851
rect 50410 53955 50454 54075
rect 51454 53955 51789 54075
rect 53789 53955 53833 54075
rect 54679 54183 54750 54971
rect 55849 54844 56051 54971
rect 55849 54798 55961 54844
rect 56007 54798 56051 54844
rect 55849 54681 56051 54798
rect 55849 54635 55961 54681
rect 56007 54635 56051 54681
rect 55849 54517 56051 54635
rect 55849 54471 55961 54517
rect 56007 54471 56051 54517
rect 55849 54354 56051 54471
rect 55849 54308 55961 54354
rect 56007 54308 56051 54354
rect 55849 54183 56051 54308
rect 33541 53562 33560 53731
rect 35133 53644 35260 53764
rect 36360 53665 36540 53764
rect 36360 53644 36475 53665
rect 35133 53595 35192 53644
rect 33336 53507 33560 53562
rect 33620 53475 33671 53595
rect 34671 53540 35192 53595
rect 36431 53540 36475 53644
rect 34671 53475 35260 53540
rect 35133 53420 35260 53475
rect 36360 53525 36475 53540
rect 36521 53525 36540 53665
rect 36360 53420 36540 53525
rect 36678 53665 36841 53764
rect 36678 53525 36697 53665
rect 36743 53644 36841 53665
rect 37501 53644 37572 53764
rect 37826 53644 37896 53764
rect 38556 53667 38734 53764
rect 43625 53731 43695 53851
rect 44325 53814 44799 53851
rect 44325 53768 44358 53814
rect 44498 53768 44799 53814
rect 44325 53731 44799 53768
rect 45323 53731 45367 53851
rect 51556 53954 51665 53955
rect 51556 53851 51600 53954
rect 38556 53644 38669 53667
rect 36743 53540 36773 53644
rect 38627 53540 38669 53644
rect 36743 53525 36841 53540
rect 36678 53420 36841 53525
rect 37501 53420 37572 53540
rect 37826 53420 37896 53540
rect 38556 53527 38669 53540
rect 38715 53527 38734 53667
rect 48603 53692 48765 53764
rect 38556 53420 38734 53527
rect 38939 53420 39008 53540
rect 39326 53420 39598 53540
rect 39730 53506 39909 53540
rect 43625 53507 43695 53627
rect 44325 53507 44799 53627
rect 45323 53583 45623 53627
rect 45323 53537 45464 53583
rect 45604 53537 45623 53583
rect 45323 53507 45623 53537
rect 48603 53552 48622 53692
rect 48668 53644 48765 53692
rect 49865 53644 49991 53764
rect 50410 53731 50454 53851
rect 51454 53731 51600 53851
rect 48668 53552 48705 53644
rect 48603 53540 48705 53552
rect 49932 53595 49991 53644
rect 49932 53540 50454 53595
rect 39730 53460 39844 53506
rect 39890 53460 39909 53506
rect 39730 53420 39909 53460
rect 48603 53420 48765 53540
rect 49865 53475 50454 53540
rect 51454 53475 51498 53595
rect 51581 53532 51600 53731
rect 51646 53851 51665 53954
rect 51646 53731 51789 53851
rect 53789 53731 53833 53851
rect 51646 53627 51667 53731
rect 51646 53532 51789 53627
rect 51581 53507 51789 53532
rect 53789 53507 53833 53627
rect 49865 53420 49991 53475
rect 29072 53044 29274 53171
rect 29072 52998 29116 53044
rect 29162 52998 29274 53044
rect 29072 52881 29274 52998
rect 29072 52835 29116 52881
rect 29162 52835 29274 52881
rect 29072 52717 29274 52835
rect 29072 52671 29116 52717
rect 29162 52671 29274 52717
rect 29072 52554 29274 52671
rect 29072 52508 29116 52554
rect 29162 52508 29274 52554
rect 29072 52383 29274 52508
rect 30373 52383 30444 53171
rect 54679 53283 54750 54071
rect 55849 53944 56051 54071
rect 55849 53898 55961 53944
rect 56007 53898 56051 53944
rect 55849 53781 56051 53898
rect 55849 53735 55961 53781
rect 56007 53735 56051 53781
rect 55849 53617 56051 53735
rect 55849 53571 55961 53617
rect 56007 53571 56051 53617
rect 55849 53454 56051 53571
rect 55849 53408 55961 53454
rect 56007 53408 56051 53454
rect 55849 53283 56051 53408
rect 35133 52979 35260 53034
rect 31292 52827 31336 52947
rect 33336 52892 33560 52947
rect 33336 52827 33495 52892
rect 33458 52723 33495 52827
rect 31292 52603 31336 52723
rect 33336 52603 33495 52723
rect 33476 52499 33495 52603
rect 29072 52144 29274 52271
rect 29072 52098 29116 52144
rect 29162 52098 29274 52144
rect 29072 51981 29274 52098
rect 29072 51935 29116 51981
rect 29162 51935 29274 51981
rect 29072 51817 29274 51935
rect 29072 51771 29116 51817
rect 29162 51771 29274 51817
rect 29072 51654 29274 51771
rect 29072 51608 29116 51654
rect 29162 51608 29274 51654
rect 29072 51483 29274 51608
rect 30373 51483 30444 52271
rect 31292 52379 31336 52499
rect 33336 52470 33495 52499
rect 33541 52723 33560 52892
rect 33620 52859 33671 52979
rect 34671 52914 35260 52979
rect 36360 52929 36540 53034
rect 36360 52914 36475 52929
rect 34671 52859 35192 52914
rect 35133 52810 35192 52859
rect 36431 52810 36475 52914
rect 33541 52603 33671 52723
rect 34671 52603 34715 52723
rect 35133 52690 35260 52810
rect 36360 52789 36475 52810
rect 36521 52789 36540 52929
rect 36360 52690 36540 52789
rect 36678 52929 36841 53034
rect 36678 52789 36697 52929
rect 36743 52914 36841 52929
rect 37501 52914 37572 53034
rect 37826 52914 37896 53034
rect 38556 52927 38734 53034
rect 38556 52914 38669 52927
rect 36743 52810 36773 52914
rect 38627 52810 38669 52914
rect 36743 52789 36841 52810
rect 36678 52690 36841 52789
rect 37501 52690 37572 52810
rect 37826 52690 37896 52810
rect 38556 52787 38669 52810
rect 38715 52787 38734 52927
rect 38939 52914 39008 53034
rect 39326 52914 39598 53034
rect 39730 52994 39909 53034
rect 39730 52948 39844 52994
rect 39890 52948 39909 52994
rect 39730 52914 39909 52948
rect 43625 52827 43695 52947
rect 44325 52827 44799 52947
rect 45323 52917 45623 52947
rect 45323 52871 45464 52917
rect 45604 52871 45623 52917
rect 45323 52827 45623 52871
rect 48603 52914 48765 53034
rect 49865 52979 49991 53034
rect 49865 52914 50454 52979
rect 48603 52902 48705 52914
rect 38556 52690 38734 52787
rect 48603 52762 48622 52902
rect 48668 52810 48705 52902
rect 49932 52859 50454 52914
rect 51454 52859 51498 52979
rect 51581 52922 51789 52947
rect 49932 52810 49991 52859
rect 48668 52762 48765 52810
rect 33541 52499 33560 52603
rect 43625 52603 43695 52723
rect 44325 52686 44799 52723
rect 44325 52640 44358 52686
rect 44498 52640 44799 52686
rect 44325 52603 44799 52640
rect 45323 52603 45367 52723
rect 48603 52690 48765 52762
rect 49865 52690 49991 52810
rect 51581 52723 51600 52922
rect 40262 52563 40346 52582
rect 40262 52517 40281 52563
rect 40327 52517 40346 52563
rect 40262 52499 40346 52517
rect 50410 52603 50454 52723
rect 51454 52603 51600 52723
rect 33541 52470 33671 52499
rect 33336 52379 33671 52470
rect 34671 52379 34715 52499
rect 31292 52155 31336 52275
rect 33336 52184 33671 52275
rect 33336 52155 33495 52184
rect 33476 52051 33495 52155
rect 31292 51931 31336 52051
rect 33336 51931 33495 52051
rect 33458 51827 33495 51931
rect 31292 51707 31336 51827
rect 33336 51762 33495 51827
rect 33541 52155 33671 52184
rect 34671 52155 34715 52275
rect 39657 52379 39727 52499
rect 40167 52379 40346 52499
rect 43354 52491 43695 52510
rect 43354 52445 43373 52491
rect 43513 52445 43695 52491
rect 43354 52390 43695 52445
rect 44325 52499 44552 52510
rect 44325 52390 44799 52499
rect 39657 52155 39727 52275
rect 40167 52155 40346 52275
rect 44451 52379 44799 52390
rect 45323 52379 45393 52499
rect 51556 52500 51600 52603
rect 51646 52827 51789 52922
rect 53789 52827 53833 52947
rect 51646 52723 51667 52827
rect 51646 52603 51789 52723
rect 53789 52603 53833 52723
rect 51646 52500 51665 52603
rect 51556 52499 51665 52500
rect 50410 52379 50454 52499
rect 51454 52379 51789 52499
rect 53789 52379 53833 52499
rect 44451 52264 44799 52275
rect 33541 52051 33560 52155
rect 40262 52137 40346 52155
rect 43354 52209 43695 52264
rect 43354 52163 43373 52209
rect 43513 52163 43695 52209
rect 43354 52144 43695 52163
rect 44325 52155 44799 52264
rect 45323 52155 45393 52275
rect 44325 52144 44552 52155
rect 40262 52091 40281 52137
rect 40327 52091 40346 52137
rect 40262 52072 40346 52091
rect 33541 51931 33671 52051
rect 34671 51931 34715 52051
rect 50410 52155 50454 52275
rect 51454 52155 51789 52275
rect 53789 52155 53833 52275
rect 54679 52383 54750 53171
rect 55849 53044 56051 53171
rect 55849 52998 55961 53044
rect 56007 52998 56051 53044
rect 55849 52881 56051 52998
rect 55849 52835 55961 52881
rect 56007 52835 56051 52881
rect 55849 52717 56051 52835
rect 55849 52671 55961 52717
rect 56007 52671 56051 52717
rect 55849 52554 56051 52671
rect 55849 52508 55961 52554
rect 56007 52508 56051 52554
rect 55849 52383 56051 52508
rect 33541 51762 33560 51931
rect 35133 51844 35260 51964
rect 36360 51865 36540 51964
rect 36360 51844 36475 51865
rect 35133 51795 35192 51844
rect 33336 51707 33560 51762
rect 33620 51675 33671 51795
rect 34671 51740 35192 51795
rect 36431 51740 36475 51844
rect 34671 51675 35260 51740
rect 35133 51620 35260 51675
rect 36360 51725 36475 51740
rect 36521 51725 36540 51865
rect 36360 51620 36540 51725
rect 36678 51865 36841 51964
rect 36678 51725 36697 51865
rect 36743 51844 36841 51865
rect 37501 51844 37572 51964
rect 37826 51844 37896 51964
rect 38556 51867 38734 51964
rect 43625 51931 43695 52051
rect 44325 52014 44799 52051
rect 44325 51968 44358 52014
rect 44498 51968 44799 52014
rect 44325 51931 44799 51968
rect 45323 51931 45367 52051
rect 51556 52154 51665 52155
rect 51556 52051 51600 52154
rect 38556 51844 38669 51867
rect 36743 51740 36773 51844
rect 38627 51740 38669 51844
rect 36743 51725 36841 51740
rect 36678 51620 36841 51725
rect 37501 51620 37572 51740
rect 37826 51620 37896 51740
rect 38556 51727 38669 51740
rect 38715 51727 38734 51867
rect 48603 51892 48765 51964
rect 38556 51620 38734 51727
rect 38939 51620 39008 51740
rect 39326 51620 39598 51740
rect 39730 51706 39909 51740
rect 43625 51707 43695 51827
rect 44325 51707 44799 51827
rect 45323 51783 45623 51827
rect 45323 51737 45464 51783
rect 45604 51737 45623 51783
rect 45323 51707 45623 51737
rect 48603 51752 48622 51892
rect 48668 51844 48765 51892
rect 49865 51844 49991 51964
rect 50410 51931 50454 52051
rect 51454 51931 51600 52051
rect 48668 51752 48705 51844
rect 48603 51740 48705 51752
rect 49932 51795 49991 51844
rect 49932 51740 50454 51795
rect 39730 51660 39844 51706
rect 39890 51660 39909 51706
rect 39730 51620 39909 51660
rect 48603 51620 48765 51740
rect 49865 51675 50454 51740
rect 51454 51675 51498 51795
rect 51581 51732 51600 51931
rect 51646 52051 51665 52154
rect 51646 51931 51789 52051
rect 53789 51931 53833 52051
rect 51646 51827 51667 51931
rect 51646 51732 51789 51827
rect 51581 51707 51789 51732
rect 53789 51707 53833 51827
rect 49865 51620 49991 51675
rect 29072 51244 29274 51371
rect 29072 51198 29116 51244
rect 29162 51198 29274 51244
rect 29072 51081 29274 51198
rect 29072 51035 29116 51081
rect 29162 51035 29274 51081
rect 29072 50917 29274 51035
rect 29072 50871 29116 50917
rect 29162 50871 29274 50917
rect 29072 50754 29274 50871
rect 29072 50708 29116 50754
rect 29162 50708 29274 50754
rect 29072 50583 29274 50708
rect 30373 50583 30444 51371
rect 54679 51483 54750 52271
rect 55849 52144 56051 52271
rect 55849 52098 55961 52144
rect 56007 52098 56051 52144
rect 55849 51981 56051 52098
rect 55849 51935 55961 51981
rect 56007 51935 56051 51981
rect 55849 51817 56051 51935
rect 55849 51771 55961 51817
rect 56007 51771 56051 51817
rect 55849 51654 56051 51771
rect 55849 51608 55961 51654
rect 56007 51608 56051 51654
rect 55849 51483 56051 51608
rect 35133 51179 35260 51234
rect 31292 51027 31336 51147
rect 33336 51092 33560 51147
rect 33336 51027 33495 51092
rect 33458 50923 33495 51027
rect 31292 50803 31336 50923
rect 33336 50803 33495 50923
rect 33476 50699 33495 50803
rect 29072 50344 29274 50471
rect 29072 50298 29116 50344
rect 29162 50298 29274 50344
rect 29072 50181 29274 50298
rect 29072 50135 29116 50181
rect 29162 50135 29274 50181
rect 29072 50017 29274 50135
rect 29072 49971 29116 50017
rect 29162 49971 29274 50017
rect 29072 49854 29274 49971
rect 29072 49808 29116 49854
rect 29162 49808 29274 49854
rect 29072 49683 29274 49808
rect 30373 49683 30444 50471
rect 31292 50579 31336 50699
rect 33336 50670 33495 50699
rect 33541 50923 33560 51092
rect 33620 51059 33671 51179
rect 34671 51114 35260 51179
rect 36360 51129 36540 51234
rect 36360 51114 36475 51129
rect 34671 51059 35192 51114
rect 35133 51010 35192 51059
rect 36431 51010 36475 51114
rect 33541 50803 33671 50923
rect 34671 50803 34715 50923
rect 35133 50890 35260 51010
rect 36360 50989 36475 51010
rect 36521 50989 36540 51129
rect 36360 50890 36540 50989
rect 36678 51129 36841 51234
rect 36678 50989 36697 51129
rect 36743 51114 36841 51129
rect 37501 51114 37572 51234
rect 37826 51114 37896 51234
rect 38556 51127 38734 51234
rect 38556 51114 38669 51127
rect 36743 51010 36773 51114
rect 38627 51010 38669 51114
rect 36743 50989 36841 51010
rect 36678 50890 36841 50989
rect 37501 50890 37572 51010
rect 37826 50890 37896 51010
rect 38556 50987 38669 51010
rect 38715 50987 38734 51127
rect 38939 51114 39008 51234
rect 39326 51114 39598 51234
rect 39730 51194 39909 51234
rect 39730 51148 39844 51194
rect 39890 51148 39909 51194
rect 39730 51114 39909 51148
rect 43625 51027 43695 51147
rect 44325 51027 44799 51147
rect 45323 51117 45623 51147
rect 45323 51071 45464 51117
rect 45604 51071 45623 51117
rect 45323 51027 45623 51071
rect 48603 51114 48765 51234
rect 49865 51179 49991 51234
rect 49865 51114 50454 51179
rect 48603 51102 48705 51114
rect 38556 50890 38734 50987
rect 48603 50962 48622 51102
rect 48668 51010 48705 51102
rect 49932 51059 50454 51114
rect 51454 51059 51498 51179
rect 51581 51122 51789 51147
rect 49932 51010 49991 51059
rect 48668 50962 48765 51010
rect 33541 50699 33560 50803
rect 43625 50803 43695 50923
rect 44325 50886 44799 50923
rect 44325 50840 44358 50886
rect 44498 50840 44799 50886
rect 44325 50803 44799 50840
rect 45323 50803 45367 50923
rect 48603 50890 48765 50962
rect 49865 50890 49991 51010
rect 51581 50923 51600 51122
rect 40262 50763 40346 50782
rect 40262 50717 40281 50763
rect 40327 50717 40346 50763
rect 40262 50699 40346 50717
rect 50410 50803 50454 50923
rect 51454 50803 51600 50923
rect 33541 50670 33671 50699
rect 33336 50579 33671 50670
rect 34671 50579 34715 50699
rect 31292 50355 31336 50475
rect 33336 50384 33671 50475
rect 33336 50355 33495 50384
rect 33476 50251 33495 50355
rect 31292 50131 31336 50251
rect 33336 50131 33495 50251
rect 33458 50027 33495 50131
rect 31292 49907 31336 50027
rect 33336 49962 33495 50027
rect 33541 50355 33671 50384
rect 34671 50355 34715 50475
rect 39657 50579 39727 50699
rect 40167 50579 40346 50699
rect 43354 50691 43695 50710
rect 43354 50645 43373 50691
rect 43513 50645 43695 50691
rect 43354 50590 43695 50645
rect 44325 50699 44552 50710
rect 44325 50590 44799 50699
rect 39657 50355 39727 50475
rect 40167 50355 40346 50475
rect 44451 50579 44799 50590
rect 45323 50579 45393 50699
rect 51556 50700 51600 50803
rect 51646 51027 51789 51122
rect 53789 51027 53833 51147
rect 51646 50923 51667 51027
rect 51646 50803 51789 50923
rect 53789 50803 53833 50923
rect 51646 50700 51665 50803
rect 51556 50699 51665 50700
rect 50410 50579 50454 50699
rect 51454 50579 51789 50699
rect 53789 50579 53833 50699
rect 44451 50464 44799 50475
rect 33541 50251 33560 50355
rect 40262 50337 40346 50355
rect 43354 50409 43695 50464
rect 43354 50363 43373 50409
rect 43513 50363 43695 50409
rect 43354 50344 43695 50363
rect 44325 50355 44799 50464
rect 45323 50355 45393 50475
rect 44325 50344 44552 50355
rect 40262 50291 40281 50337
rect 40327 50291 40346 50337
rect 40262 50272 40346 50291
rect 33541 50131 33671 50251
rect 34671 50131 34715 50251
rect 50410 50355 50454 50475
rect 51454 50355 51789 50475
rect 53789 50355 53833 50475
rect 54679 50583 54750 51371
rect 55849 51244 56051 51371
rect 55849 51198 55961 51244
rect 56007 51198 56051 51244
rect 55849 51081 56051 51198
rect 55849 51035 55961 51081
rect 56007 51035 56051 51081
rect 55849 50917 56051 51035
rect 55849 50871 55961 50917
rect 56007 50871 56051 50917
rect 55849 50754 56051 50871
rect 55849 50708 55961 50754
rect 56007 50708 56051 50754
rect 55849 50583 56051 50708
rect 33541 49962 33560 50131
rect 35133 50044 35260 50164
rect 36360 50065 36540 50164
rect 36360 50044 36475 50065
rect 35133 49995 35192 50044
rect 33336 49907 33560 49962
rect 33620 49875 33671 49995
rect 34671 49940 35192 49995
rect 36431 49940 36475 50044
rect 34671 49875 35260 49940
rect 35133 49820 35260 49875
rect 36360 49925 36475 49940
rect 36521 49925 36540 50065
rect 36360 49820 36540 49925
rect 36678 50065 36841 50164
rect 36678 49925 36697 50065
rect 36743 50044 36841 50065
rect 37501 50044 37572 50164
rect 37826 50044 37896 50164
rect 38556 50067 38734 50164
rect 43625 50131 43695 50251
rect 44325 50214 44799 50251
rect 44325 50168 44358 50214
rect 44498 50168 44799 50214
rect 44325 50131 44799 50168
rect 45323 50131 45367 50251
rect 51556 50354 51665 50355
rect 51556 50251 51600 50354
rect 38556 50044 38669 50067
rect 36743 49940 36773 50044
rect 38627 49940 38669 50044
rect 36743 49925 36841 49940
rect 36678 49820 36841 49925
rect 37501 49820 37572 49940
rect 37826 49820 37896 49940
rect 38556 49927 38669 49940
rect 38715 49927 38734 50067
rect 48603 50092 48765 50164
rect 38556 49820 38734 49927
rect 38939 49820 39008 49940
rect 39326 49820 39598 49940
rect 39730 49906 39909 49940
rect 43625 49907 43695 50027
rect 44325 49907 44799 50027
rect 45323 49983 45623 50027
rect 45323 49937 45464 49983
rect 45604 49937 45623 49983
rect 45323 49907 45623 49937
rect 48603 49952 48622 50092
rect 48668 50044 48765 50092
rect 49865 50044 49991 50164
rect 50410 50131 50454 50251
rect 51454 50131 51600 50251
rect 48668 49952 48705 50044
rect 48603 49940 48705 49952
rect 49932 49995 49991 50044
rect 49932 49940 50454 49995
rect 39730 49860 39844 49906
rect 39890 49860 39909 49906
rect 39730 49820 39909 49860
rect 48603 49820 48765 49940
rect 49865 49875 50454 49940
rect 51454 49875 51498 49995
rect 51581 49932 51600 50131
rect 51646 50251 51665 50354
rect 51646 50131 51789 50251
rect 53789 50131 53833 50251
rect 51646 50027 51667 50131
rect 51646 49932 51789 50027
rect 51581 49907 51789 49932
rect 53789 49907 53833 50027
rect 49865 49820 49991 49875
rect 29072 49444 29274 49571
rect 29072 49398 29116 49444
rect 29162 49398 29274 49444
rect 29072 49281 29274 49398
rect 29072 49235 29116 49281
rect 29162 49235 29274 49281
rect 29072 49117 29274 49235
rect 29072 49071 29116 49117
rect 29162 49071 29274 49117
rect 29072 48954 29274 49071
rect 29072 48908 29116 48954
rect 29162 48908 29274 48954
rect 29072 48783 29274 48908
rect 30373 48783 30444 49571
rect 54679 49683 54750 50471
rect 55849 50344 56051 50471
rect 55849 50298 55961 50344
rect 56007 50298 56051 50344
rect 55849 50181 56051 50298
rect 55849 50135 55961 50181
rect 56007 50135 56051 50181
rect 55849 50017 56051 50135
rect 55849 49971 55961 50017
rect 56007 49971 56051 50017
rect 55849 49854 56051 49971
rect 55849 49808 55961 49854
rect 56007 49808 56051 49854
rect 55849 49683 56051 49808
rect 35133 49379 35260 49434
rect 31292 49227 31336 49347
rect 33336 49292 33560 49347
rect 33336 49227 33495 49292
rect 33458 49123 33495 49227
rect 31292 49003 31336 49123
rect 33336 49003 33495 49123
rect 33476 48899 33495 49003
rect 29072 48544 29274 48671
rect 29072 48498 29116 48544
rect 29162 48498 29274 48544
rect 29072 48381 29274 48498
rect 29072 48335 29116 48381
rect 29162 48335 29274 48381
rect 29072 48217 29274 48335
rect 29072 48171 29116 48217
rect 29162 48171 29274 48217
rect 29072 48054 29274 48171
rect 29072 48008 29116 48054
rect 29162 48008 29274 48054
rect 29072 47883 29274 48008
rect 30373 47883 30444 48671
rect 31292 48779 31336 48899
rect 33336 48870 33495 48899
rect 33541 49123 33560 49292
rect 33620 49259 33671 49379
rect 34671 49314 35260 49379
rect 36360 49329 36540 49434
rect 36360 49314 36475 49329
rect 34671 49259 35192 49314
rect 35133 49210 35192 49259
rect 36431 49210 36475 49314
rect 33541 49003 33671 49123
rect 34671 49003 34715 49123
rect 35133 49090 35260 49210
rect 36360 49189 36475 49210
rect 36521 49189 36540 49329
rect 36360 49090 36540 49189
rect 36678 49329 36841 49434
rect 36678 49189 36697 49329
rect 36743 49314 36841 49329
rect 37501 49314 37572 49434
rect 37826 49314 37896 49434
rect 38556 49327 38734 49434
rect 38556 49314 38669 49327
rect 36743 49210 36773 49314
rect 38627 49210 38669 49314
rect 36743 49189 36841 49210
rect 36678 49090 36841 49189
rect 37501 49090 37572 49210
rect 37826 49090 37896 49210
rect 38556 49187 38669 49210
rect 38715 49187 38734 49327
rect 38939 49314 39008 49434
rect 39326 49314 39598 49434
rect 39730 49394 39909 49434
rect 39730 49348 39844 49394
rect 39890 49348 39909 49394
rect 39730 49314 39909 49348
rect 43625 49227 43695 49347
rect 44325 49227 44799 49347
rect 45323 49317 45623 49347
rect 45323 49271 45464 49317
rect 45604 49271 45623 49317
rect 45323 49227 45623 49271
rect 48603 49314 48765 49434
rect 49865 49379 49991 49434
rect 49865 49314 50454 49379
rect 48603 49302 48705 49314
rect 38556 49090 38734 49187
rect 48603 49162 48622 49302
rect 48668 49210 48705 49302
rect 49932 49259 50454 49314
rect 51454 49259 51498 49379
rect 51581 49322 51789 49347
rect 49932 49210 49991 49259
rect 48668 49162 48765 49210
rect 33541 48899 33560 49003
rect 43625 49003 43695 49123
rect 44325 49086 44799 49123
rect 44325 49040 44358 49086
rect 44498 49040 44799 49086
rect 44325 49003 44799 49040
rect 45323 49003 45367 49123
rect 48603 49090 48765 49162
rect 49865 49090 49991 49210
rect 51581 49123 51600 49322
rect 40262 48963 40346 48982
rect 40262 48917 40281 48963
rect 40327 48917 40346 48963
rect 40262 48899 40346 48917
rect 50410 49003 50454 49123
rect 51454 49003 51600 49123
rect 33541 48870 33671 48899
rect 33336 48779 33671 48870
rect 34671 48779 34715 48899
rect 31292 48555 31336 48675
rect 33336 48584 33671 48675
rect 33336 48555 33495 48584
rect 33476 48451 33495 48555
rect 31292 48331 31336 48451
rect 33336 48331 33495 48451
rect 33458 48227 33495 48331
rect 31292 48107 31336 48227
rect 33336 48162 33495 48227
rect 33541 48555 33671 48584
rect 34671 48555 34715 48675
rect 39657 48779 39727 48899
rect 40167 48779 40346 48899
rect 43354 48891 43695 48910
rect 43354 48845 43373 48891
rect 43513 48845 43695 48891
rect 43354 48790 43695 48845
rect 44325 48899 44552 48910
rect 44325 48790 44799 48899
rect 39657 48555 39727 48675
rect 40167 48555 40346 48675
rect 44451 48779 44799 48790
rect 45323 48779 45393 48899
rect 51556 48900 51600 49003
rect 51646 49227 51789 49322
rect 53789 49227 53833 49347
rect 51646 49123 51667 49227
rect 51646 49003 51789 49123
rect 53789 49003 53833 49123
rect 51646 48900 51665 49003
rect 51556 48899 51665 48900
rect 50410 48779 50454 48899
rect 51454 48779 51789 48899
rect 53789 48779 53833 48899
rect 44451 48664 44799 48675
rect 33541 48451 33560 48555
rect 40262 48537 40346 48555
rect 43354 48609 43695 48664
rect 43354 48563 43373 48609
rect 43513 48563 43695 48609
rect 43354 48544 43695 48563
rect 44325 48555 44799 48664
rect 45323 48555 45393 48675
rect 44325 48544 44552 48555
rect 40262 48491 40281 48537
rect 40327 48491 40346 48537
rect 40262 48472 40346 48491
rect 33541 48331 33671 48451
rect 34671 48331 34715 48451
rect 50410 48555 50454 48675
rect 51454 48555 51789 48675
rect 53789 48555 53833 48675
rect 54679 48783 54750 49571
rect 55849 49444 56051 49571
rect 55849 49398 55961 49444
rect 56007 49398 56051 49444
rect 55849 49281 56051 49398
rect 55849 49235 55961 49281
rect 56007 49235 56051 49281
rect 55849 49117 56051 49235
rect 55849 49071 55961 49117
rect 56007 49071 56051 49117
rect 55849 48954 56051 49071
rect 55849 48908 55961 48954
rect 56007 48908 56051 48954
rect 55849 48783 56051 48908
rect 33541 48162 33560 48331
rect 35133 48244 35260 48364
rect 36360 48265 36540 48364
rect 36360 48244 36475 48265
rect 35133 48195 35192 48244
rect 33336 48107 33560 48162
rect 33620 48075 33671 48195
rect 34671 48140 35192 48195
rect 36431 48140 36475 48244
rect 34671 48075 35260 48140
rect 35133 48020 35260 48075
rect 36360 48125 36475 48140
rect 36521 48125 36540 48265
rect 36360 48020 36540 48125
rect 36678 48265 36841 48364
rect 36678 48125 36697 48265
rect 36743 48244 36841 48265
rect 37501 48244 37572 48364
rect 37826 48244 37896 48364
rect 38556 48267 38734 48364
rect 43625 48331 43695 48451
rect 44325 48414 44799 48451
rect 44325 48368 44358 48414
rect 44498 48368 44799 48414
rect 44325 48331 44799 48368
rect 45323 48331 45367 48451
rect 51556 48554 51665 48555
rect 51556 48451 51600 48554
rect 38556 48244 38669 48267
rect 36743 48140 36773 48244
rect 38627 48140 38669 48244
rect 36743 48125 36841 48140
rect 36678 48020 36841 48125
rect 37501 48020 37572 48140
rect 37826 48020 37896 48140
rect 38556 48127 38669 48140
rect 38715 48127 38734 48267
rect 48603 48292 48765 48364
rect 38556 48020 38734 48127
rect 38939 48020 39008 48140
rect 39326 48020 39598 48140
rect 39730 48106 39909 48140
rect 43625 48107 43695 48227
rect 44325 48107 44799 48227
rect 45323 48183 45623 48227
rect 45323 48137 45464 48183
rect 45604 48137 45623 48183
rect 45323 48107 45623 48137
rect 48603 48152 48622 48292
rect 48668 48244 48765 48292
rect 49865 48244 49991 48364
rect 50410 48331 50454 48451
rect 51454 48331 51600 48451
rect 48668 48152 48705 48244
rect 48603 48140 48705 48152
rect 49932 48195 49991 48244
rect 49932 48140 50454 48195
rect 39730 48060 39844 48106
rect 39890 48060 39909 48106
rect 39730 48020 39909 48060
rect 48603 48020 48765 48140
rect 49865 48075 50454 48140
rect 51454 48075 51498 48195
rect 51581 48132 51600 48331
rect 51646 48451 51665 48554
rect 51646 48331 51789 48451
rect 53789 48331 53833 48451
rect 51646 48227 51667 48331
rect 51646 48132 51789 48227
rect 51581 48107 51789 48132
rect 53789 48107 53833 48227
rect 49865 48020 49991 48075
rect 29072 47644 29274 47771
rect 29072 47598 29116 47644
rect 29162 47598 29274 47644
rect 29072 47481 29274 47598
rect 29072 47435 29116 47481
rect 29162 47435 29274 47481
rect 29072 47317 29274 47435
rect 29072 47271 29116 47317
rect 29162 47271 29274 47317
rect 29072 47154 29274 47271
rect 29072 47108 29116 47154
rect 29162 47108 29274 47154
rect 29072 46983 29274 47108
rect 30373 46983 30444 47771
rect 54679 47883 54750 48671
rect 55849 48544 56051 48671
rect 55849 48498 55961 48544
rect 56007 48498 56051 48544
rect 55849 48381 56051 48498
rect 55849 48335 55961 48381
rect 56007 48335 56051 48381
rect 55849 48217 56051 48335
rect 55849 48171 55961 48217
rect 56007 48171 56051 48217
rect 55849 48054 56051 48171
rect 55849 48008 55961 48054
rect 56007 48008 56051 48054
rect 55849 47883 56051 48008
rect 35133 47579 35260 47634
rect 31292 47427 31336 47547
rect 33336 47492 33560 47547
rect 33336 47427 33495 47492
rect 33458 47323 33495 47427
rect 31292 47203 31336 47323
rect 33336 47203 33495 47323
rect 33476 47099 33495 47203
rect 29072 46744 29274 46871
rect 29072 46698 29116 46744
rect 29162 46698 29274 46744
rect 29072 46581 29274 46698
rect 29072 46535 29116 46581
rect 29162 46535 29274 46581
rect 29072 46417 29274 46535
rect 29072 46371 29116 46417
rect 29162 46371 29274 46417
rect 29072 46254 29274 46371
rect 29072 46208 29116 46254
rect 29162 46208 29274 46254
rect 29072 46083 29274 46208
rect 30373 46083 30444 46871
rect 31292 46979 31336 47099
rect 33336 47070 33495 47099
rect 33541 47323 33560 47492
rect 33620 47459 33671 47579
rect 34671 47514 35260 47579
rect 36360 47529 36540 47634
rect 36360 47514 36475 47529
rect 34671 47459 35192 47514
rect 35133 47410 35192 47459
rect 36431 47410 36475 47514
rect 33541 47203 33671 47323
rect 34671 47203 34715 47323
rect 35133 47290 35260 47410
rect 36360 47389 36475 47410
rect 36521 47389 36540 47529
rect 36360 47290 36540 47389
rect 36678 47529 36841 47634
rect 36678 47389 36697 47529
rect 36743 47514 36841 47529
rect 37501 47514 37572 47634
rect 37826 47514 37896 47634
rect 38556 47527 38734 47634
rect 38556 47514 38669 47527
rect 36743 47410 36773 47514
rect 38627 47410 38669 47514
rect 36743 47389 36841 47410
rect 36678 47290 36841 47389
rect 37501 47290 37572 47410
rect 37826 47290 37896 47410
rect 38556 47387 38669 47410
rect 38715 47387 38734 47527
rect 38939 47514 39008 47634
rect 39326 47514 39598 47634
rect 39730 47594 39909 47634
rect 39730 47548 39844 47594
rect 39890 47548 39909 47594
rect 39730 47514 39909 47548
rect 43625 47427 43695 47547
rect 44325 47427 44799 47547
rect 45323 47517 45623 47547
rect 45323 47471 45464 47517
rect 45604 47471 45623 47517
rect 45323 47427 45623 47471
rect 48603 47514 48765 47634
rect 49865 47579 49991 47634
rect 49865 47514 50454 47579
rect 48603 47502 48705 47514
rect 38556 47290 38734 47387
rect 48603 47362 48622 47502
rect 48668 47410 48705 47502
rect 49932 47459 50454 47514
rect 51454 47459 51498 47579
rect 51581 47522 51789 47547
rect 49932 47410 49991 47459
rect 48668 47362 48765 47410
rect 33541 47099 33560 47203
rect 43625 47203 43695 47323
rect 44325 47286 44799 47323
rect 44325 47240 44358 47286
rect 44498 47240 44799 47286
rect 44325 47203 44799 47240
rect 45323 47203 45367 47323
rect 48603 47290 48765 47362
rect 49865 47290 49991 47410
rect 51581 47323 51600 47522
rect 40262 47163 40346 47182
rect 40262 47117 40281 47163
rect 40327 47117 40346 47163
rect 40262 47099 40346 47117
rect 50410 47203 50454 47323
rect 51454 47203 51600 47323
rect 33541 47070 33671 47099
rect 33336 46979 33671 47070
rect 34671 46979 34715 47099
rect 31292 46755 31336 46875
rect 33336 46784 33671 46875
rect 33336 46755 33495 46784
rect 33476 46651 33495 46755
rect 31292 46531 31336 46651
rect 33336 46531 33495 46651
rect 33458 46427 33495 46531
rect 31292 46307 31336 46427
rect 33336 46362 33495 46427
rect 33541 46755 33671 46784
rect 34671 46755 34715 46875
rect 39657 46979 39727 47099
rect 40167 46979 40346 47099
rect 43354 47091 43695 47110
rect 43354 47045 43373 47091
rect 43513 47045 43695 47091
rect 43354 46990 43695 47045
rect 44325 47099 44552 47110
rect 44325 46990 44799 47099
rect 39657 46755 39727 46875
rect 40167 46755 40346 46875
rect 44451 46979 44799 46990
rect 45323 46979 45393 47099
rect 51556 47100 51600 47203
rect 51646 47427 51789 47522
rect 53789 47427 53833 47547
rect 51646 47323 51667 47427
rect 51646 47203 51789 47323
rect 53789 47203 53833 47323
rect 51646 47100 51665 47203
rect 51556 47099 51665 47100
rect 50410 46979 50454 47099
rect 51454 46979 51789 47099
rect 53789 46979 53833 47099
rect 44451 46864 44799 46875
rect 33541 46651 33560 46755
rect 40262 46737 40346 46755
rect 43354 46809 43695 46864
rect 43354 46763 43373 46809
rect 43513 46763 43695 46809
rect 43354 46744 43695 46763
rect 44325 46755 44799 46864
rect 45323 46755 45393 46875
rect 44325 46744 44552 46755
rect 40262 46691 40281 46737
rect 40327 46691 40346 46737
rect 40262 46672 40346 46691
rect 33541 46531 33671 46651
rect 34671 46531 34715 46651
rect 50410 46755 50454 46875
rect 51454 46755 51789 46875
rect 53789 46755 53833 46875
rect 54679 46983 54750 47771
rect 55849 47644 56051 47771
rect 55849 47598 55961 47644
rect 56007 47598 56051 47644
rect 55849 47481 56051 47598
rect 55849 47435 55961 47481
rect 56007 47435 56051 47481
rect 55849 47317 56051 47435
rect 55849 47271 55961 47317
rect 56007 47271 56051 47317
rect 55849 47154 56051 47271
rect 55849 47108 55961 47154
rect 56007 47108 56051 47154
rect 55849 46983 56051 47108
rect 33541 46362 33560 46531
rect 35133 46444 35260 46564
rect 36360 46465 36540 46564
rect 36360 46444 36475 46465
rect 35133 46395 35192 46444
rect 33336 46307 33560 46362
rect 33620 46275 33671 46395
rect 34671 46340 35192 46395
rect 36431 46340 36475 46444
rect 34671 46275 35260 46340
rect 35133 46220 35260 46275
rect 36360 46325 36475 46340
rect 36521 46325 36540 46465
rect 36360 46220 36540 46325
rect 36678 46465 36841 46564
rect 36678 46325 36697 46465
rect 36743 46444 36841 46465
rect 37501 46444 37572 46564
rect 37826 46444 37896 46564
rect 38556 46467 38734 46564
rect 43625 46531 43695 46651
rect 44325 46614 44799 46651
rect 44325 46568 44358 46614
rect 44498 46568 44799 46614
rect 44325 46531 44799 46568
rect 45323 46531 45367 46651
rect 51556 46754 51665 46755
rect 51556 46651 51600 46754
rect 38556 46444 38669 46467
rect 36743 46340 36773 46444
rect 38627 46340 38669 46444
rect 36743 46325 36841 46340
rect 36678 46220 36841 46325
rect 37501 46220 37572 46340
rect 37826 46220 37896 46340
rect 38556 46327 38669 46340
rect 38715 46327 38734 46467
rect 48603 46492 48765 46564
rect 38556 46220 38734 46327
rect 38939 46220 39008 46340
rect 39326 46220 39598 46340
rect 39730 46306 39909 46340
rect 43625 46307 43695 46427
rect 44325 46307 44799 46427
rect 45323 46383 45623 46427
rect 45323 46337 45464 46383
rect 45604 46337 45623 46383
rect 45323 46307 45623 46337
rect 48603 46352 48622 46492
rect 48668 46444 48765 46492
rect 49865 46444 49991 46564
rect 50410 46531 50454 46651
rect 51454 46531 51600 46651
rect 48668 46352 48705 46444
rect 48603 46340 48705 46352
rect 49932 46395 49991 46444
rect 49932 46340 50454 46395
rect 39730 46260 39844 46306
rect 39890 46260 39909 46306
rect 39730 46220 39909 46260
rect 48603 46220 48765 46340
rect 49865 46275 50454 46340
rect 51454 46275 51498 46395
rect 51581 46332 51600 46531
rect 51646 46651 51665 46754
rect 51646 46531 51789 46651
rect 53789 46531 53833 46651
rect 51646 46427 51667 46531
rect 51646 46332 51789 46427
rect 51581 46307 51789 46332
rect 53789 46307 53833 46427
rect 49865 46220 49991 46275
rect 29072 45844 29274 45971
rect 29072 45798 29116 45844
rect 29162 45798 29274 45844
rect 29072 45681 29274 45798
rect 29072 45635 29116 45681
rect 29162 45635 29274 45681
rect 29072 45517 29274 45635
rect 29072 45471 29116 45517
rect 29162 45471 29274 45517
rect 29072 45354 29274 45471
rect 29072 45308 29116 45354
rect 29162 45308 29274 45354
rect 29072 45183 29274 45308
rect 30373 45183 30444 45971
rect 54679 46083 54750 46871
rect 55849 46744 56051 46871
rect 55849 46698 55961 46744
rect 56007 46698 56051 46744
rect 55849 46581 56051 46698
rect 55849 46535 55961 46581
rect 56007 46535 56051 46581
rect 55849 46417 56051 46535
rect 55849 46371 55961 46417
rect 56007 46371 56051 46417
rect 55849 46254 56051 46371
rect 55849 46208 55961 46254
rect 56007 46208 56051 46254
rect 55849 46083 56051 46208
rect 35133 45779 35260 45834
rect 31292 45627 31336 45747
rect 33336 45692 33560 45747
rect 33336 45627 33495 45692
rect 33458 45523 33495 45627
rect 31292 45403 31336 45523
rect 33336 45403 33495 45523
rect 33476 45299 33495 45403
rect 29072 44944 29274 45071
rect 29072 44898 29116 44944
rect 29162 44898 29274 44944
rect 29072 44781 29274 44898
rect 29072 44735 29116 44781
rect 29162 44735 29274 44781
rect 29072 44617 29274 44735
rect 29072 44571 29116 44617
rect 29162 44571 29274 44617
rect 29072 44454 29274 44571
rect 29072 44408 29116 44454
rect 29162 44408 29274 44454
rect 29072 44283 29274 44408
rect 30373 44283 30444 45071
rect 31292 45179 31336 45299
rect 33336 45270 33495 45299
rect 33541 45523 33560 45692
rect 33620 45659 33671 45779
rect 34671 45714 35260 45779
rect 36360 45729 36540 45834
rect 36360 45714 36475 45729
rect 34671 45659 35192 45714
rect 35133 45610 35192 45659
rect 36431 45610 36475 45714
rect 33541 45403 33671 45523
rect 34671 45403 34715 45523
rect 35133 45490 35260 45610
rect 36360 45589 36475 45610
rect 36521 45589 36540 45729
rect 36360 45490 36540 45589
rect 36678 45729 36841 45834
rect 36678 45589 36697 45729
rect 36743 45714 36841 45729
rect 37501 45714 37572 45834
rect 37826 45714 37896 45834
rect 38556 45727 38734 45834
rect 38556 45714 38669 45727
rect 36743 45610 36773 45714
rect 38627 45610 38669 45714
rect 36743 45589 36841 45610
rect 36678 45490 36841 45589
rect 37501 45490 37572 45610
rect 37826 45490 37896 45610
rect 38556 45587 38669 45610
rect 38715 45587 38734 45727
rect 38939 45714 39008 45834
rect 39326 45714 39598 45834
rect 39730 45794 39909 45834
rect 39730 45748 39844 45794
rect 39890 45748 39909 45794
rect 39730 45714 39909 45748
rect 43625 45627 43695 45747
rect 44325 45627 44799 45747
rect 45323 45717 45623 45747
rect 45323 45671 45464 45717
rect 45604 45671 45623 45717
rect 45323 45627 45623 45671
rect 48603 45714 48765 45834
rect 49865 45779 49991 45834
rect 49865 45714 50454 45779
rect 48603 45702 48705 45714
rect 38556 45490 38734 45587
rect 48603 45562 48622 45702
rect 48668 45610 48705 45702
rect 49932 45659 50454 45714
rect 51454 45659 51498 45779
rect 51581 45722 51789 45747
rect 49932 45610 49991 45659
rect 48668 45562 48765 45610
rect 33541 45299 33560 45403
rect 43625 45403 43695 45523
rect 44325 45486 44799 45523
rect 44325 45440 44358 45486
rect 44498 45440 44799 45486
rect 44325 45403 44799 45440
rect 45323 45403 45367 45523
rect 48603 45490 48765 45562
rect 49865 45490 49991 45610
rect 51581 45523 51600 45722
rect 40262 45363 40346 45382
rect 40262 45317 40281 45363
rect 40327 45317 40346 45363
rect 40262 45299 40346 45317
rect 50410 45403 50454 45523
rect 51454 45403 51600 45523
rect 33541 45270 33671 45299
rect 33336 45179 33671 45270
rect 34671 45179 34715 45299
rect 31292 44955 31336 45075
rect 33336 44984 33671 45075
rect 33336 44955 33495 44984
rect 33476 44851 33495 44955
rect 31292 44731 31336 44851
rect 33336 44731 33495 44851
rect 33458 44627 33495 44731
rect 31292 44507 31336 44627
rect 33336 44562 33495 44627
rect 33541 44955 33671 44984
rect 34671 44955 34715 45075
rect 39657 45179 39727 45299
rect 40167 45179 40346 45299
rect 43354 45291 43695 45310
rect 43354 45245 43373 45291
rect 43513 45245 43695 45291
rect 43354 45190 43695 45245
rect 44325 45299 44552 45310
rect 44325 45190 44799 45299
rect 39657 44955 39727 45075
rect 40167 44955 40346 45075
rect 44451 45179 44799 45190
rect 45323 45179 45393 45299
rect 51556 45300 51600 45403
rect 51646 45627 51789 45722
rect 53789 45627 53833 45747
rect 51646 45523 51667 45627
rect 51646 45403 51789 45523
rect 53789 45403 53833 45523
rect 51646 45300 51665 45403
rect 51556 45299 51665 45300
rect 50410 45179 50454 45299
rect 51454 45179 51789 45299
rect 53789 45179 53833 45299
rect 44451 45064 44799 45075
rect 33541 44851 33560 44955
rect 40262 44937 40346 44955
rect 43354 45009 43695 45064
rect 43354 44963 43373 45009
rect 43513 44963 43695 45009
rect 43354 44944 43695 44963
rect 44325 44955 44799 45064
rect 45323 44955 45393 45075
rect 44325 44944 44552 44955
rect 40262 44891 40281 44937
rect 40327 44891 40346 44937
rect 40262 44872 40346 44891
rect 33541 44731 33671 44851
rect 34671 44731 34715 44851
rect 50410 44955 50454 45075
rect 51454 44955 51789 45075
rect 53789 44955 53833 45075
rect 54679 45183 54750 45971
rect 55849 45844 56051 45971
rect 55849 45798 55961 45844
rect 56007 45798 56051 45844
rect 55849 45681 56051 45798
rect 55849 45635 55961 45681
rect 56007 45635 56051 45681
rect 55849 45517 56051 45635
rect 55849 45471 55961 45517
rect 56007 45471 56051 45517
rect 55849 45354 56051 45471
rect 55849 45308 55961 45354
rect 56007 45308 56051 45354
rect 55849 45183 56051 45308
rect 33541 44562 33560 44731
rect 35133 44644 35260 44764
rect 36360 44665 36540 44764
rect 36360 44644 36475 44665
rect 35133 44595 35192 44644
rect 33336 44507 33560 44562
rect 33620 44475 33671 44595
rect 34671 44540 35192 44595
rect 36431 44540 36475 44644
rect 34671 44475 35260 44540
rect 35133 44420 35260 44475
rect 36360 44525 36475 44540
rect 36521 44525 36540 44665
rect 36360 44420 36540 44525
rect 36678 44665 36841 44764
rect 36678 44525 36697 44665
rect 36743 44644 36841 44665
rect 37501 44644 37572 44764
rect 37826 44644 37896 44764
rect 38556 44667 38734 44764
rect 43625 44731 43695 44851
rect 44325 44814 44799 44851
rect 44325 44768 44358 44814
rect 44498 44768 44799 44814
rect 44325 44731 44799 44768
rect 45323 44731 45367 44851
rect 51556 44954 51665 44955
rect 51556 44851 51600 44954
rect 38556 44644 38669 44667
rect 36743 44540 36773 44644
rect 38627 44540 38669 44644
rect 36743 44525 36841 44540
rect 36678 44420 36841 44525
rect 37501 44420 37572 44540
rect 37826 44420 37896 44540
rect 38556 44527 38669 44540
rect 38715 44527 38734 44667
rect 48603 44692 48765 44764
rect 38556 44420 38734 44527
rect 38939 44420 39008 44540
rect 39326 44420 39598 44540
rect 39730 44506 39909 44540
rect 43625 44507 43695 44627
rect 44325 44507 44799 44627
rect 45323 44583 45623 44627
rect 45323 44537 45464 44583
rect 45604 44537 45623 44583
rect 45323 44507 45623 44537
rect 48603 44552 48622 44692
rect 48668 44644 48765 44692
rect 49865 44644 49991 44764
rect 50410 44731 50454 44851
rect 51454 44731 51600 44851
rect 48668 44552 48705 44644
rect 48603 44540 48705 44552
rect 49932 44595 49991 44644
rect 49932 44540 50454 44595
rect 39730 44460 39844 44506
rect 39890 44460 39909 44506
rect 39730 44420 39909 44460
rect 48603 44420 48765 44540
rect 49865 44475 50454 44540
rect 51454 44475 51498 44595
rect 51581 44532 51600 44731
rect 51646 44851 51665 44954
rect 51646 44731 51789 44851
rect 53789 44731 53833 44851
rect 51646 44627 51667 44731
rect 51646 44532 51789 44627
rect 51581 44507 51789 44532
rect 53789 44507 53833 44627
rect 49865 44420 49991 44475
rect 29072 44044 29274 44171
rect 29072 43998 29116 44044
rect 29162 43998 29274 44044
rect 29072 43881 29274 43998
rect 29072 43835 29116 43881
rect 29162 43835 29274 43881
rect 29072 43717 29274 43835
rect 29072 43671 29116 43717
rect 29162 43671 29274 43717
rect 29072 43554 29274 43671
rect 29072 43508 29116 43554
rect 29162 43508 29274 43554
rect 29072 43383 29274 43508
rect 30373 43383 30444 44171
rect 54679 44283 54750 45071
rect 55849 44944 56051 45071
rect 55849 44898 55961 44944
rect 56007 44898 56051 44944
rect 55849 44781 56051 44898
rect 55849 44735 55961 44781
rect 56007 44735 56051 44781
rect 55849 44617 56051 44735
rect 55849 44571 55961 44617
rect 56007 44571 56051 44617
rect 55849 44454 56051 44571
rect 55849 44408 55961 44454
rect 56007 44408 56051 44454
rect 55849 44283 56051 44408
rect 35133 43979 35260 44034
rect 31292 43827 31336 43947
rect 33336 43892 33560 43947
rect 33336 43827 33495 43892
rect 33458 43723 33495 43827
rect 31292 43603 31336 43723
rect 33336 43603 33495 43723
rect 33476 43499 33495 43603
rect 29072 43144 29274 43271
rect 29072 43098 29116 43144
rect 29162 43098 29274 43144
rect 29072 42981 29274 43098
rect 29072 42935 29116 42981
rect 29162 42935 29274 42981
rect 29072 42817 29274 42935
rect 29072 42771 29116 42817
rect 29162 42771 29274 42817
rect 29072 42654 29274 42771
rect 29072 42608 29116 42654
rect 29162 42608 29274 42654
rect 29072 42483 29274 42608
rect 30373 42483 30444 43271
rect 31292 43379 31336 43499
rect 33336 43470 33495 43499
rect 33541 43723 33560 43892
rect 33620 43859 33671 43979
rect 34671 43914 35260 43979
rect 36360 43929 36540 44034
rect 36360 43914 36475 43929
rect 34671 43859 35192 43914
rect 35133 43810 35192 43859
rect 36431 43810 36475 43914
rect 33541 43603 33671 43723
rect 34671 43603 34715 43723
rect 35133 43690 35260 43810
rect 36360 43789 36475 43810
rect 36521 43789 36540 43929
rect 36360 43690 36540 43789
rect 36678 43929 36841 44034
rect 36678 43789 36697 43929
rect 36743 43914 36841 43929
rect 37501 43914 37572 44034
rect 37826 43914 37896 44034
rect 38556 43927 38734 44034
rect 38556 43914 38669 43927
rect 36743 43810 36773 43914
rect 38627 43810 38669 43914
rect 36743 43789 36841 43810
rect 36678 43690 36841 43789
rect 37501 43690 37572 43810
rect 37826 43690 37896 43810
rect 38556 43787 38669 43810
rect 38715 43787 38734 43927
rect 38939 43914 39008 44034
rect 39326 43914 39598 44034
rect 39730 43994 39909 44034
rect 39730 43948 39844 43994
rect 39890 43948 39909 43994
rect 39730 43914 39909 43948
rect 43625 43827 43695 43947
rect 44325 43827 44799 43947
rect 45323 43917 45623 43947
rect 45323 43871 45464 43917
rect 45604 43871 45623 43917
rect 45323 43827 45623 43871
rect 48603 43914 48765 44034
rect 49865 43979 49991 44034
rect 49865 43914 50454 43979
rect 48603 43902 48705 43914
rect 38556 43690 38734 43787
rect 48603 43762 48622 43902
rect 48668 43810 48705 43902
rect 49932 43859 50454 43914
rect 51454 43859 51498 43979
rect 51581 43922 51789 43947
rect 49932 43810 49991 43859
rect 48668 43762 48765 43810
rect 33541 43499 33560 43603
rect 43625 43603 43695 43723
rect 44325 43686 44799 43723
rect 44325 43640 44358 43686
rect 44498 43640 44799 43686
rect 44325 43603 44799 43640
rect 45323 43603 45367 43723
rect 48603 43690 48765 43762
rect 49865 43690 49991 43810
rect 51581 43723 51600 43922
rect 40262 43563 40346 43582
rect 40262 43517 40281 43563
rect 40327 43517 40346 43563
rect 40262 43499 40346 43517
rect 50410 43603 50454 43723
rect 51454 43603 51600 43723
rect 33541 43470 33671 43499
rect 33336 43379 33671 43470
rect 34671 43379 34715 43499
rect 31292 43155 31336 43275
rect 33336 43184 33671 43275
rect 33336 43155 33495 43184
rect 33476 43051 33495 43155
rect 31292 42931 31336 43051
rect 33336 42931 33495 43051
rect 33458 42827 33495 42931
rect 31292 42707 31336 42827
rect 33336 42762 33495 42827
rect 33541 43155 33671 43184
rect 34671 43155 34715 43275
rect 39657 43379 39727 43499
rect 40167 43379 40346 43499
rect 43354 43491 43695 43510
rect 43354 43445 43373 43491
rect 43513 43445 43695 43491
rect 43354 43390 43695 43445
rect 44325 43499 44552 43510
rect 44325 43390 44799 43499
rect 39657 43155 39727 43275
rect 40167 43155 40346 43275
rect 44451 43379 44799 43390
rect 45323 43379 45393 43499
rect 51556 43500 51600 43603
rect 51646 43827 51789 43922
rect 53789 43827 53833 43947
rect 51646 43723 51667 43827
rect 51646 43603 51789 43723
rect 53789 43603 53833 43723
rect 51646 43500 51665 43603
rect 51556 43499 51665 43500
rect 50410 43379 50454 43499
rect 51454 43379 51789 43499
rect 53789 43379 53833 43499
rect 44451 43264 44799 43275
rect 33541 43051 33560 43155
rect 40262 43137 40346 43155
rect 43354 43209 43695 43264
rect 43354 43163 43373 43209
rect 43513 43163 43695 43209
rect 43354 43144 43695 43163
rect 44325 43155 44799 43264
rect 45323 43155 45393 43275
rect 44325 43144 44552 43155
rect 40262 43091 40281 43137
rect 40327 43091 40346 43137
rect 40262 43072 40346 43091
rect 33541 42931 33671 43051
rect 34671 42931 34715 43051
rect 50410 43155 50454 43275
rect 51454 43155 51789 43275
rect 53789 43155 53833 43275
rect 54679 43383 54750 44171
rect 55849 44044 56051 44171
rect 55849 43998 55961 44044
rect 56007 43998 56051 44044
rect 55849 43881 56051 43998
rect 55849 43835 55961 43881
rect 56007 43835 56051 43881
rect 55849 43717 56051 43835
rect 55849 43671 55961 43717
rect 56007 43671 56051 43717
rect 55849 43554 56051 43671
rect 55849 43508 55961 43554
rect 56007 43508 56051 43554
rect 55849 43383 56051 43508
rect 33541 42762 33560 42931
rect 35133 42844 35260 42964
rect 36360 42865 36540 42964
rect 36360 42844 36475 42865
rect 35133 42795 35192 42844
rect 33336 42707 33560 42762
rect 33620 42675 33671 42795
rect 34671 42740 35192 42795
rect 36431 42740 36475 42844
rect 34671 42675 35260 42740
rect 35133 42620 35260 42675
rect 36360 42725 36475 42740
rect 36521 42725 36540 42865
rect 36360 42620 36540 42725
rect 36678 42865 36841 42964
rect 36678 42725 36697 42865
rect 36743 42844 36841 42865
rect 37501 42844 37572 42964
rect 37826 42844 37896 42964
rect 38556 42867 38734 42964
rect 43625 42931 43695 43051
rect 44325 43014 44799 43051
rect 44325 42968 44358 43014
rect 44498 42968 44799 43014
rect 44325 42931 44799 42968
rect 45323 42931 45367 43051
rect 51556 43154 51665 43155
rect 51556 43051 51600 43154
rect 38556 42844 38669 42867
rect 36743 42740 36773 42844
rect 38627 42740 38669 42844
rect 36743 42725 36841 42740
rect 36678 42620 36841 42725
rect 37501 42620 37572 42740
rect 37826 42620 37896 42740
rect 38556 42727 38669 42740
rect 38715 42727 38734 42867
rect 48603 42892 48765 42964
rect 38556 42620 38734 42727
rect 38939 42620 39008 42740
rect 39326 42620 39598 42740
rect 39730 42706 39909 42740
rect 43625 42707 43695 42827
rect 44325 42707 44799 42827
rect 45323 42783 45623 42827
rect 45323 42737 45464 42783
rect 45604 42737 45623 42783
rect 45323 42707 45623 42737
rect 48603 42752 48622 42892
rect 48668 42844 48765 42892
rect 49865 42844 49991 42964
rect 50410 42931 50454 43051
rect 51454 42931 51600 43051
rect 48668 42752 48705 42844
rect 48603 42740 48705 42752
rect 49932 42795 49991 42844
rect 49932 42740 50454 42795
rect 39730 42660 39844 42706
rect 39890 42660 39909 42706
rect 39730 42620 39909 42660
rect 48603 42620 48765 42740
rect 49865 42675 50454 42740
rect 51454 42675 51498 42795
rect 51581 42732 51600 42931
rect 51646 43051 51665 43154
rect 51646 42931 51789 43051
rect 53789 42931 53833 43051
rect 51646 42827 51667 42931
rect 51646 42732 51789 42827
rect 51581 42707 51789 42732
rect 53789 42707 53833 42827
rect 49865 42620 49991 42675
rect 29072 42244 29274 42371
rect 29072 42198 29116 42244
rect 29162 42198 29274 42244
rect 29072 42081 29274 42198
rect 29072 42035 29116 42081
rect 29162 42035 29274 42081
rect 29072 41917 29274 42035
rect 29072 41871 29116 41917
rect 29162 41871 29274 41917
rect 29072 41754 29274 41871
rect 29072 41708 29116 41754
rect 29162 41708 29274 41754
rect 29072 41583 29274 41708
rect 30373 41583 30444 42371
rect 54679 42483 54750 43271
rect 55849 43144 56051 43271
rect 55849 43098 55961 43144
rect 56007 43098 56051 43144
rect 55849 42981 56051 43098
rect 55849 42935 55961 42981
rect 56007 42935 56051 42981
rect 55849 42817 56051 42935
rect 55849 42771 55961 42817
rect 56007 42771 56051 42817
rect 55849 42654 56051 42771
rect 55849 42608 55961 42654
rect 56007 42608 56051 42654
rect 55849 42483 56051 42608
rect 35133 42179 35260 42234
rect 31292 42027 31336 42147
rect 33336 42092 33560 42147
rect 33336 42027 33495 42092
rect 33458 41923 33495 42027
rect 31292 41803 31336 41923
rect 33336 41803 33495 41923
rect 33476 41699 33495 41803
rect 29072 41344 29274 41471
rect 29072 41298 29116 41344
rect 29162 41298 29274 41344
rect 29072 41181 29274 41298
rect 29072 41135 29116 41181
rect 29162 41135 29274 41181
rect 29072 41017 29274 41135
rect 29072 40971 29116 41017
rect 29162 40971 29274 41017
rect 29072 40854 29274 40971
rect 29072 40808 29116 40854
rect 29162 40808 29274 40854
rect 29072 40683 29274 40808
rect 30373 40683 30444 41471
rect 31292 41579 31336 41699
rect 33336 41670 33495 41699
rect 33541 41923 33560 42092
rect 33620 42059 33671 42179
rect 34671 42114 35260 42179
rect 36360 42129 36540 42234
rect 36360 42114 36475 42129
rect 34671 42059 35192 42114
rect 35133 42010 35192 42059
rect 36431 42010 36475 42114
rect 33541 41803 33671 41923
rect 34671 41803 34715 41923
rect 35133 41890 35260 42010
rect 36360 41989 36475 42010
rect 36521 41989 36540 42129
rect 36360 41890 36540 41989
rect 36678 42129 36841 42234
rect 36678 41989 36697 42129
rect 36743 42114 36841 42129
rect 37501 42114 37572 42234
rect 37826 42114 37896 42234
rect 38556 42127 38734 42234
rect 38556 42114 38669 42127
rect 36743 42010 36773 42114
rect 38627 42010 38669 42114
rect 36743 41989 36841 42010
rect 36678 41890 36841 41989
rect 37501 41890 37572 42010
rect 37826 41890 37896 42010
rect 38556 41987 38669 42010
rect 38715 41987 38734 42127
rect 38939 42114 39008 42234
rect 39326 42114 39598 42234
rect 39730 42194 39909 42234
rect 39730 42148 39844 42194
rect 39890 42148 39909 42194
rect 39730 42114 39909 42148
rect 43625 42027 43695 42147
rect 44325 42027 44799 42147
rect 45323 42117 45623 42147
rect 45323 42071 45464 42117
rect 45604 42071 45623 42117
rect 45323 42027 45623 42071
rect 48603 42114 48765 42234
rect 49865 42179 49991 42234
rect 49865 42114 50454 42179
rect 48603 42102 48705 42114
rect 38556 41890 38734 41987
rect 48603 41962 48622 42102
rect 48668 42010 48705 42102
rect 49932 42059 50454 42114
rect 51454 42059 51498 42179
rect 51581 42122 51789 42147
rect 49932 42010 49991 42059
rect 48668 41962 48765 42010
rect 33541 41699 33560 41803
rect 43625 41803 43695 41923
rect 44325 41886 44799 41923
rect 44325 41840 44358 41886
rect 44498 41840 44799 41886
rect 44325 41803 44799 41840
rect 45323 41803 45367 41923
rect 48603 41890 48765 41962
rect 49865 41890 49991 42010
rect 51581 41923 51600 42122
rect 40262 41763 40346 41782
rect 40262 41717 40281 41763
rect 40327 41717 40346 41763
rect 40262 41699 40346 41717
rect 50410 41803 50454 41923
rect 51454 41803 51600 41923
rect 33541 41670 33671 41699
rect 33336 41579 33671 41670
rect 34671 41579 34715 41699
rect 31292 41355 31336 41475
rect 33336 41384 33671 41475
rect 33336 41355 33495 41384
rect 33476 41251 33495 41355
rect 31292 41131 31336 41251
rect 33336 41131 33495 41251
rect 33458 41027 33495 41131
rect 31292 40907 31336 41027
rect 33336 40962 33495 41027
rect 33541 41355 33671 41384
rect 34671 41355 34715 41475
rect 39657 41579 39727 41699
rect 40167 41579 40346 41699
rect 43354 41691 43695 41710
rect 43354 41645 43373 41691
rect 43513 41645 43695 41691
rect 43354 41590 43695 41645
rect 44325 41699 44552 41710
rect 44325 41590 44799 41699
rect 39657 41355 39727 41475
rect 40167 41355 40346 41475
rect 44451 41579 44799 41590
rect 45323 41579 45393 41699
rect 51556 41700 51600 41803
rect 51646 42027 51789 42122
rect 53789 42027 53833 42147
rect 51646 41923 51667 42027
rect 51646 41803 51789 41923
rect 53789 41803 53833 41923
rect 51646 41700 51665 41803
rect 51556 41699 51665 41700
rect 50410 41579 50454 41699
rect 51454 41579 51789 41699
rect 53789 41579 53833 41699
rect 44451 41464 44799 41475
rect 33541 41251 33560 41355
rect 40262 41337 40346 41355
rect 43354 41409 43695 41464
rect 43354 41363 43373 41409
rect 43513 41363 43695 41409
rect 43354 41344 43695 41363
rect 44325 41355 44799 41464
rect 45323 41355 45393 41475
rect 44325 41344 44552 41355
rect 40262 41291 40281 41337
rect 40327 41291 40346 41337
rect 40262 41272 40346 41291
rect 33541 41131 33671 41251
rect 34671 41131 34715 41251
rect 50410 41355 50454 41475
rect 51454 41355 51789 41475
rect 53789 41355 53833 41475
rect 54679 41583 54750 42371
rect 55849 42244 56051 42371
rect 55849 42198 55961 42244
rect 56007 42198 56051 42244
rect 55849 42081 56051 42198
rect 55849 42035 55961 42081
rect 56007 42035 56051 42081
rect 55849 41917 56051 42035
rect 55849 41871 55961 41917
rect 56007 41871 56051 41917
rect 55849 41754 56051 41871
rect 55849 41708 55961 41754
rect 56007 41708 56051 41754
rect 55849 41583 56051 41708
rect 33541 40962 33560 41131
rect 35133 41044 35260 41164
rect 36360 41065 36540 41164
rect 36360 41044 36475 41065
rect 35133 40995 35192 41044
rect 33336 40907 33560 40962
rect 33620 40875 33671 40995
rect 34671 40940 35192 40995
rect 36431 40940 36475 41044
rect 34671 40875 35260 40940
rect 35133 40820 35260 40875
rect 36360 40925 36475 40940
rect 36521 40925 36540 41065
rect 36360 40820 36540 40925
rect 36678 41065 36841 41164
rect 36678 40925 36697 41065
rect 36743 41044 36841 41065
rect 37501 41044 37572 41164
rect 37826 41044 37896 41164
rect 38556 41067 38734 41164
rect 43625 41131 43695 41251
rect 44325 41214 44799 41251
rect 44325 41168 44358 41214
rect 44498 41168 44799 41214
rect 44325 41131 44799 41168
rect 45323 41131 45367 41251
rect 51556 41354 51665 41355
rect 51556 41251 51600 41354
rect 38556 41044 38669 41067
rect 36743 40940 36773 41044
rect 38627 40940 38669 41044
rect 36743 40925 36841 40940
rect 36678 40820 36841 40925
rect 37501 40820 37572 40940
rect 37826 40820 37896 40940
rect 38556 40927 38669 40940
rect 38715 40927 38734 41067
rect 48603 41092 48765 41164
rect 38556 40820 38734 40927
rect 38939 40820 39008 40940
rect 39326 40820 39598 40940
rect 39730 40906 39909 40940
rect 43625 40907 43695 41027
rect 44325 40907 44799 41027
rect 45323 40983 45623 41027
rect 45323 40937 45464 40983
rect 45604 40937 45623 40983
rect 45323 40907 45623 40937
rect 48603 40952 48622 41092
rect 48668 41044 48765 41092
rect 49865 41044 49991 41164
rect 50410 41131 50454 41251
rect 51454 41131 51600 41251
rect 48668 40952 48705 41044
rect 48603 40940 48705 40952
rect 49932 40995 49991 41044
rect 49932 40940 50454 40995
rect 39730 40860 39844 40906
rect 39890 40860 39909 40906
rect 39730 40820 39909 40860
rect 48603 40820 48765 40940
rect 49865 40875 50454 40940
rect 51454 40875 51498 40995
rect 51581 40932 51600 41131
rect 51646 41251 51665 41354
rect 51646 41131 51789 41251
rect 53789 41131 53833 41251
rect 51646 41027 51667 41131
rect 51646 40932 51789 41027
rect 51581 40907 51789 40932
rect 53789 40907 53833 41027
rect 49865 40820 49991 40875
rect 29072 40444 29274 40571
rect 29072 40398 29116 40444
rect 29162 40398 29274 40444
rect 29072 40281 29274 40398
rect 29072 40235 29116 40281
rect 29162 40235 29274 40281
rect 29072 40117 29274 40235
rect 29072 40071 29116 40117
rect 29162 40071 29274 40117
rect 29072 39954 29274 40071
rect 29072 39908 29116 39954
rect 29162 39908 29274 39954
rect 29072 39783 29274 39908
rect 30373 39783 30444 40571
rect 54679 40683 54750 41471
rect 55849 41344 56051 41471
rect 55849 41298 55961 41344
rect 56007 41298 56051 41344
rect 55849 41181 56051 41298
rect 55849 41135 55961 41181
rect 56007 41135 56051 41181
rect 55849 41017 56051 41135
rect 55849 40971 55961 41017
rect 56007 40971 56051 41017
rect 55849 40854 56051 40971
rect 55849 40808 55961 40854
rect 56007 40808 56051 40854
rect 55849 40683 56051 40808
rect 35133 40379 35260 40434
rect 31292 40227 31336 40347
rect 33336 40292 33560 40347
rect 33336 40227 33495 40292
rect 33458 40123 33495 40227
rect 31292 40003 31336 40123
rect 33336 40003 33495 40123
rect 33476 39899 33495 40003
rect 29072 39544 29274 39671
rect 29072 39498 29116 39544
rect 29162 39498 29274 39544
rect 29072 39381 29274 39498
rect 29072 39335 29116 39381
rect 29162 39335 29274 39381
rect 29072 39217 29274 39335
rect 29072 39171 29116 39217
rect 29162 39171 29274 39217
rect 29072 39054 29274 39171
rect 29072 39008 29116 39054
rect 29162 39008 29274 39054
rect 29072 38883 29274 39008
rect 30373 38883 30444 39671
rect 31292 39779 31336 39899
rect 33336 39870 33495 39899
rect 33541 40123 33560 40292
rect 33620 40259 33671 40379
rect 34671 40314 35260 40379
rect 36360 40329 36540 40434
rect 36360 40314 36475 40329
rect 34671 40259 35192 40314
rect 35133 40210 35192 40259
rect 36431 40210 36475 40314
rect 33541 40003 33671 40123
rect 34671 40003 34715 40123
rect 35133 40090 35260 40210
rect 36360 40189 36475 40210
rect 36521 40189 36540 40329
rect 36360 40090 36540 40189
rect 36678 40329 36841 40434
rect 36678 40189 36697 40329
rect 36743 40314 36841 40329
rect 37501 40314 37572 40434
rect 37826 40314 37896 40434
rect 38556 40327 38734 40434
rect 38556 40314 38669 40327
rect 36743 40210 36773 40314
rect 38627 40210 38669 40314
rect 36743 40189 36841 40210
rect 36678 40090 36841 40189
rect 37501 40090 37572 40210
rect 37826 40090 37896 40210
rect 38556 40187 38669 40210
rect 38715 40187 38734 40327
rect 38939 40314 39008 40434
rect 39326 40314 39598 40434
rect 39730 40394 39909 40434
rect 39730 40348 39844 40394
rect 39890 40348 39909 40394
rect 39730 40314 39909 40348
rect 43625 40227 43695 40347
rect 44325 40227 44799 40347
rect 45323 40317 45623 40347
rect 45323 40271 45464 40317
rect 45604 40271 45623 40317
rect 45323 40227 45623 40271
rect 48603 40314 48765 40434
rect 49865 40379 49991 40434
rect 49865 40314 50454 40379
rect 48603 40302 48705 40314
rect 38556 40090 38734 40187
rect 48603 40162 48622 40302
rect 48668 40210 48705 40302
rect 49932 40259 50454 40314
rect 51454 40259 51498 40379
rect 51581 40322 51789 40347
rect 49932 40210 49991 40259
rect 48668 40162 48765 40210
rect 33541 39899 33560 40003
rect 43625 40003 43695 40123
rect 44325 40086 44799 40123
rect 44325 40040 44358 40086
rect 44498 40040 44799 40086
rect 44325 40003 44799 40040
rect 45323 40003 45367 40123
rect 48603 40090 48765 40162
rect 49865 40090 49991 40210
rect 51581 40123 51600 40322
rect 40262 39963 40346 39982
rect 40262 39917 40281 39963
rect 40327 39917 40346 39963
rect 40262 39899 40346 39917
rect 50410 40003 50454 40123
rect 51454 40003 51600 40123
rect 33541 39870 33671 39899
rect 33336 39779 33671 39870
rect 34671 39779 34715 39899
rect 31292 39555 31336 39675
rect 33336 39584 33671 39675
rect 33336 39555 33495 39584
rect 33476 39451 33495 39555
rect 31292 39331 31336 39451
rect 33336 39331 33495 39451
rect 33458 39227 33495 39331
rect 31292 39107 31336 39227
rect 33336 39162 33495 39227
rect 33541 39555 33671 39584
rect 34671 39555 34715 39675
rect 39657 39779 39727 39899
rect 40167 39779 40346 39899
rect 43354 39891 43695 39910
rect 43354 39845 43373 39891
rect 43513 39845 43695 39891
rect 43354 39790 43695 39845
rect 44325 39899 44552 39910
rect 44325 39790 44799 39899
rect 39657 39555 39727 39675
rect 40167 39555 40346 39675
rect 44451 39779 44799 39790
rect 45323 39779 45393 39899
rect 51556 39900 51600 40003
rect 51646 40227 51789 40322
rect 53789 40227 53833 40347
rect 51646 40123 51667 40227
rect 51646 40003 51789 40123
rect 53789 40003 53833 40123
rect 51646 39900 51665 40003
rect 51556 39899 51665 39900
rect 50410 39779 50454 39899
rect 51454 39779 51789 39899
rect 53789 39779 53833 39899
rect 44451 39664 44799 39675
rect 33541 39451 33560 39555
rect 40262 39537 40346 39555
rect 43354 39609 43695 39664
rect 43354 39563 43373 39609
rect 43513 39563 43695 39609
rect 43354 39544 43695 39563
rect 44325 39555 44799 39664
rect 45323 39555 45393 39675
rect 44325 39544 44552 39555
rect 40262 39491 40281 39537
rect 40327 39491 40346 39537
rect 40262 39472 40346 39491
rect 33541 39331 33671 39451
rect 34671 39331 34715 39451
rect 50410 39555 50454 39675
rect 51454 39555 51789 39675
rect 53789 39555 53833 39675
rect 54679 39783 54750 40571
rect 55849 40444 56051 40571
rect 55849 40398 55961 40444
rect 56007 40398 56051 40444
rect 55849 40281 56051 40398
rect 55849 40235 55961 40281
rect 56007 40235 56051 40281
rect 55849 40117 56051 40235
rect 55849 40071 55961 40117
rect 56007 40071 56051 40117
rect 55849 39954 56051 40071
rect 55849 39908 55961 39954
rect 56007 39908 56051 39954
rect 55849 39783 56051 39908
rect 33541 39162 33560 39331
rect 35133 39244 35260 39364
rect 36360 39265 36540 39364
rect 36360 39244 36475 39265
rect 35133 39195 35192 39244
rect 33336 39107 33560 39162
rect 33620 39075 33671 39195
rect 34671 39140 35192 39195
rect 36431 39140 36475 39244
rect 34671 39075 35260 39140
rect 35133 39020 35260 39075
rect 36360 39125 36475 39140
rect 36521 39125 36540 39265
rect 36360 39020 36540 39125
rect 36678 39265 36841 39364
rect 36678 39125 36697 39265
rect 36743 39244 36841 39265
rect 37501 39244 37572 39364
rect 37826 39244 37896 39364
rect 38556 39267 38734 39364
rect 43625 39331 43695 39451
rect 44325 39414 44799 39451
rect 44325 39368 44358 39414
rect 44498 39368 44799 39414
rect 44325 39331 44799 39368
rect 45323 39331 45367 39451
rect 51556 39554 51665 39555
rect 51556 39451 51600 39554
rect 38556 39244 38669 39267
rect 36743 39140 36773 39244
rect 38627 39140 38669 39244
rect 36743 39125 36841 39140
rect 36678 39020 36841 39125
rect 37501 39020 37572 39140
rect 37826 39020 37896 39140
rect 38556 39127 38669 39140
rect 38715 39127 38734 39267
rect 48603 39292 48765 39364
rect 38556 39020 38734 39127
rect 38939 39020 39008 39140
rect 39326 39020 39598 39140
rect 39730 39106 39909 39140
rect 43625 39107 43695 39227
rect 44325 39107 44799 39227
rect 45323 39183 45623 39227
rect 45323 39137 45464 39183
rect 45604 39137 45623 39183
rect 45323 39107 45623 39137
rect 48603 39152 48622 39292
rect 48668 39244 48765 39292
rect 49865 39244 49991 39364
rect 50410 39331 50454 39451
rect 51454 39331 51600 39451
rect 48668 39152 48705 39244
rect 48603 39140 48705 39152
rect 49932 39195 49991 39244
rect 49932 39140 50454 39195
rect 39730 39060 39844 39106
rect 39890 39060 39909 39106
rect 39730 39020 39909 39060
rect 48603 39020 48765 39140
rect 49865 39075 50454 39140
rect 51454 39075 51498 39195
rect 51581 39132 51600 39331
rect 51646 39451 51665 39554
rect 51646 39331 51789 39451
rect 53789 39331 53833 39451
rect 51646 39227 51667 39331
rect 51646 39132 51789 39227
rect 51581 39107 51789 39132
rect 53789 39107 53833 39227
rect 49865 39020 49991 39075
rect 29072 38644 29274 38771
rect 29072 38598 29116 38644
rect 29162 38598 29274 38644
rect 29072 38481 29274 38598
rect 29072 38435 29116 38481
rect 29162 38435 29274 38481
rect 29072 38317 29274 38435
rect 29072 38271 29116 38317
rect 29162 38271 29274 38317
rect 29072 38154 29274 38271
rect 29072 38108 29116 38154
rect 29162 38108 29274 38154
rect 29072 37983 29274 38108
rect 30373 37983 30444 38771
rect 54679 38883 54750 39671
rect 55849 39544 56051 39671
rect 55849 39498 55961 39544
rect 56007 39498 56051 39544
rect 55849 39381 56051 39498
rect 55849 39335 55961 39381
rect 56007 39335 56051 39381
rect 55849 39217 56051 39335
rect 55849 39171 55961 39217
rect 56007 39171 56051 39217
rect 55849 39054 56051 39171
rect 55849 39008 55961 39054
rect 56007 39008 56051 39054
rect 55849 38883 56051 39008
rect 35133 38579 35260 38634
rect 31292 38427 31336 38547
rect 33336 38492 33560 38547
rect 33336 38427 33495 38492
rect 33458 38323 33495 38427
rect 31292 38203 31336 38323
rect 33336 38203 33495 38323
rect 33476 38099 33495 38203
rect 29072 37744 29274 37871
rect 29072 37698 29116 37744
rect 29162 37698 29274 37744
rect 29072 37581 29274 37698
rect 29072 37535 29116 37581
rect 29162 37535 29274 37581
rect 29072 37417 29274 37535
rect 29072 37371 29116 37417
rect 29162 37371 29274 37417
rect 29072 37254 29274 37371
rect 29072 37208 29116 37254
rect 29162 37208 29274 37254
rect 29072 37083 29274 37208
rect 30373 37083 30444 37871
rect 31292 37979 31336 38099
rect 33336 38070 33495 38099
rect 33541 38323 33560 38492
rect 33620 38459 33671 38579
rect 34671 38514 35260 38579
rect 36360 38529 36540 38634
rect 36360 38514 36475 38529
rect 34671 38459 35192 38514
rect 35133 38410 35192 38459
rect 36431 38410 36475 38514
rect 33541 38203 33671 38323
rect 34671 38203 34715 38323
rect 35133 38290 35260 38410
rect 36360 38389 36475 38410
rect 36521 38389 36540 38529
rect 36360 38290 36540 38389
rect 36678 38529 36841 38634
rect 36678 38389 36697 38529
rect 36743 38514 36841 38529
rect 37501 38514 37572 38634
rect 37826 38514 37896 38634
rect 38556 38527 38734 38634
rect 38556 38514 38669 38527
rect 36743 38410 36773 38514
rect 38627 38410 38669 38514
rect 36743 38389 36841 38410
rect 36678 38290 36841 38389
rect 37501 38290 37572 38410
rect 37826 38290 37896 38410
rect 38556 38387 38669 38410
rect 38715 38387 38734 38527
rect 38939 38514 39008 38634
rect 39326 38514 39598 38634
rect 39730 38594 39909 38634
rect 39730 38548 39844 38594
rect 39890 38548 39909 38594
rect 39730 38514 39909 38548
rect 43625 38427 43695 38547
rect 44325 38427 44799 38547
rect 45323 38517 45623 38547
rect 45323 38471 45464 38517
rect 45604 38471 45623 38517
rect 45323 38427 45623 38471
rect 48603 38514 48765 38634
rect 49865 38579 49991 38634
rect 49865 38514 50454 38579
rect 48603 38502 48705 38514
rect 38556 38290 38734 38387
rect 48603 38362 48622 38502
rect 48668 38410 48705 38502
rect 49932 38459 50454 38514
rect 51454 38459 51498 38579
rect 51581 38522 51789 38547
rect 49932 38410 49991 38459
rect 48668 38362 48765 38410
rect 33541 38099 33560 38203
rect 43625 38203 43695 38323
rect 44325 38286 44799 38323
rect 44325 38240 44358 38286
rect 44498 38240 44799 38286
rect 44325 38203 44799 38240
rect 45323 38203 45367 38323
rect 48603 38290 48765 38362
rect 49865 38290 49991 38410
rect 51581 38323 51600 38522
rect 40262 38163 40346 38182
rect 40262 38117 40281 38163
rect 40327 38117 40346 38163
rect 40262 38099 40346 38117
rect 50410 38203 50454 38323
rect 51454 38203 51600 38323
rect 33541 38070 33671 38099
rect 33336 37979 33671 38070
rect 34671 37979 34715 38099
rect 31292 37755 31336 37875
rect 33336 37784 33671 37875
rect 33336 37755 33495 37784
rect 33476 37651 33495 37755
rect 31292 37531 31336 37651
rect 33336 37531 33495 37651
rect 33458 37427 33495 37531
rect 31292 37307 31336 37427
rect 33336 37362 33495 37427
rect 33541 37755 33671 37784
rect 34671 37755 34715 37875
rect 39657 37979 39727 38099
rect 40167 37979 40346 38099
rect 43354 38091 43695 38110
rect 43354 38045 43373 38091
rect 43513 38045 43695 38091
rect 43354 37990 43695 38045
rect 44325 38099 44552 38110
rect 44325 37990 44799 38099
rect 39657 37755 39727 37875
rect 40167 37755 40346 37875
rect 44451 37979 44799 37990
rect 45323 37979 45393 38099
rect 51556 38100 51600 38203
rect 51646 38427 51789 38522
rect 53789 38427 53833 38547
rect 51646 38323 51667 38427
rect 51646 38203 51789 38323
rect 53789 38203 53833 38323
rect 51646 38100 51665 38203
rect 51556 38099 51665 38100
rect 50410 37979 50454 38099
rect 51454 37979 51789 38099
rect 53789 37979 53833 38099
rect 44451 37864 44799 37875
rect 33541 37651 33560 37755
rect 40262 37737 40346 37755
rect 43354 37809 43695 37864
rect 43354 37763 43373 37809
rect 43513 37763 43695 37809
rect 43354 37744 43695 37763
rect 44325 37755 44799 37864
rect 45323 37755 45393 37875
rect 44325 37744 44552 37755
rect 40262 37691 40281 37737
rect 40327 37691 40346 37737
rect 40262 37672 40346 37691
rect 33541 37531 33671 37651
rect 34671 37531 34715 37651
rect 50410 37755 50454 37875
rect 51454 37755 51789 37875
rect 53789 37755 53833 37875
rect 54679 37983 54750 38771
rect 55849 38644 56051 38771
rect 55849 38598 55961 38644
rect 56007 38598 56051 38644
rect 55849 38481 56051 38598
rect 55849 38435 55961 38481
rect 56007 38435 56051 38481
rect 55849 38317 56051 38435
rect 55849 38271 55961 38317
rect 56007 38271 56051 38317
rect 55849 38154 56051 38271
rect 55849 38108 55961 38154
rect 56007 38108 56051 38154
rect 55849 37983 56051 38108
rect 33541 37362 33560 37531
rect 35133 37444 35260 37564
rect 36360 37465 36540 37564
rect 36360 37444 36475 37465
rect 35133 37395 35192 37444
rect 33336 37307 33560 37362
rect 33620 37275 33671 37395
rect 34671 37340 35192 37395
rect 36431 37340 36475 37444
rect 34671 37275 35260 37340
rect 35133 37220 35260 37275
rect 36360 37325 36475 37340
rect 36521 37325 36540 37465
rect 36360 37220 36540 37325
rect 36678 37465 36841 37564
rect 36678 37325 36697 37465
rect 36743 37444 36841 37465
rect 37501 37444 37572 37564
rect 37826 37444 37896 37564
rect 38556 37467 38734 37564
rect 43625 37531 43695 37651
rect 44325 37614 44799 37651
rect 44325 37568 44358 37614
rect 44498 37568 44799 37614
rect 44325 37531 44799 37568
rect 45323 37531 45367 37651
rect 51556 37754 51665 37755
rect 51556 37651 51600 37754
rect 38556 37444 38669 37467
rect 36743 37340 36773 37444
rect 38627 37340 38669 37444
rect 36743 37325 36841 37340
rect 36678 37220 36841 37325
rect 37501 37220 37572 37340
rect 37826 37220 37896 37340
rect 38556 37327 38669 37340
rect 38715 37327 38734 37467
rect 48603 37492 48765 37564
rect 38556 37220 38734 37327
rect 38939 37220 39008 37340
rect 39326 37220 39598 37340
rect 39730 37306 39909 37340
rect 43625 37307 43695 37427
rect 44325 37307 44799 37427
rect 45323 37383 45623 37427
rect 45323 37337 45464 37383
rect 45604 37337 45623 37383
rect 45323 37307 45623 37337
rect 48603 37352 48622 37492
rect 48668 37444 48765 37492
rect 49865 37444 49991 37564
rect 50410 37531 50454 37651
rect 51454 37531 51600 37651
rect 48668 37352 48705 37444
rect 48603 37340 48705 37352
rect 49932 37395 49991 37444
rect 49932 37340 50454 37395
rect 39730 37260 39844 37306
rect 39890 37260 39909 37306
rect 39730 37220 39909 37260
rect 48603 37220 48765 37340
rect 49865 37275 50454 37340
rect 51454 37275 51498 37395
rect 51581 37332 51600 37531
rect 51646 37651 51665 37754
rect 51646 37531 51789 37651
rect 53789 37531 53833 37651
rect 51646 37427 51667 37531
rect 51646 37332 51789 37427
rect 51581 37307 51789 37332
rect 53789 37307 53833 37427
rect 49865 37220 49991 37275
rect 29072 36844 29274 36971
rect 29072 36798 29116 36844
rect 29162 36798 29274 36844
rect 29072 36681 29274 36798
rect 29072 36635 29116 36681
rect 29162 36635 29274 36681
rect 29072 36517 29274 36635
rect 29072 36471 29116 36517
rect 29162 36471 29274 36517
rect 29072 36354 29274 36471
rect 29072 36308 29116 36354
rect 29162 36308 29274 36354
rect 29072 36183 29274 36308
rect 30373 36183 30444 36971
rect 54679 37083 54750 37871
rect 55849 37744 56051 37871
rect 55849 37698 55961 37744
rect 56007 37698 56051 37744
rect 55849 37581 56051 37698
rect 55849 37535 55961 37581
rect 56007 37535 56051 37581
rect 55849 37417 56051 37535
rect 55849 37371 55961 37417
rect 56007 37371 56051 37417
rect 55849 37254 56051 37371
rect 55849 37208 55961 37254
rect 56007 37208 56051 37254
rect 55849 37083 56051 37208
rect 35133 36779 35260 36834
rect 31292 36627 31336 36747
rect 33336 36692 33560 36747
rect 33336 36627 33495 36692
rect 33458 36523 33495 36627
rect 31292 36403 31336 36523
rect 33336 36403 33495 36523
rect 33476 36299 33495 36403
rect 31292 36179 31336 36299
rect 33336 36270 33495 36299
rect 33541 36523 33560 36692
rect 33620 36659 33671 36779
rect 34671 36714 35260 36779
rect 36360 36729 36540 36834
rect 36360 36714 36475 36729
rect 34671 36659 35192 36714
rect 35133 36610 35192 36659
rect 36431 36610 36475 36714
rect 33541 36403 33671 36523
rect 34671 36403 34715 36523
rect 35133 36490 35260 36610
rect 36360 36589 36475 36610
rect 36521 36589 36540 36729
rect 36360 36490 36540 36589
rect 36678 36729 36841 36834
rect 36678 36589 36697 36729
rect 36743 36714 36841 36729
rect 37501 36714 37572 36834
rect 37826 36714 37896 36834
rect 38556 36727 38734 36834
rect 38556 36714 38669 36727
rect 36743 36610 36773 36714
rect 38627 36610 38669 36714
rect 36743 36589 36841 36610
rect 36678 36490 36841 36589
rect 37501 36490 37572 36610
rect 37826 36490 37896 36610
rect 38556 36587 38669 36610
rect 38715 36587 38734 36727
rect 38939 36714 39008 36834
rect 39326 36714 39598 36834
rect 39730 36794 39909 36834
rect 39730 36748 39844 36794
rect 39890 36748 39909 36794
rect 39730 36714 39909 36748
rect 43625 36627 43695 36747
rect 44325 36627 44799 36747
rect 45323 36717 45623 36747
rect 45323 36671 45464 36717
rect 45604 36671 45623 36717
rect 45323 36627 45623 36671
rect 48603 36714 48765 36834
rect 49865 36779 49991 36834
rect 49865 36714 50454 36779
rect 48603 36702 48705 36714
rect 38556 36490 38734 36587
rect 48603 36562 48622 36702
rect 48668 36610 48705 36702
rect 49932 36659 50454 36714
rect 51454 36659 51498 36779
rect 51581 36722 51789 36747
rect 49932 36610 49991 36659
rect 48668 36562 48765 36610
rect 33541 36299 33560 36403
rect 43625 36403 43695 36523
rect 44325 36486 44799 36523
rect 44325 36440 44358 36486
rect 44498 36440 44799 36486
rect 44325 36403 44799 36440
rect 45323 36403 45367 36523
rect 48603 36490 48765 36562
rect 49865 36490 49991 36610
rect 51581 36523 51600 36722
rect 40262 36363 40346 36382
rect 40262 36317 40281 36363
rect 40327 36317 40346 36363
rect 40262 36299 40346 36317
rect 50410 36403 50454 36523
rect 51454 36403 51600 36523
rect 33541 36270 33671 36299
rect 33336 36179 33671 36270
rect 34671 36179 34715 36299
rect 39657 36179 39727 36299
rect 40167 36179 40346 36299
rect 43354 36291 43695 36310
rect 43354 36245 43373 36291
rect 43513 36245 43695 36291
rect 43354 36190 43695 36245
rect 44325 36299 44552 36310
rect 44325 36190 44799 36299
rect 44451 36179 44799 36190
rect 45323 36179 45393 36299
rect 51556 36300 51600 36403
rect 51646 36627 51789 36722
rect 53789 36627 53833 36747
rect 51646 36523 51667 36627
rect 51646 36403 51789 36523
rect 53789 36403 53833 36523
rect 51646 36300 51665 36403
rect 51556 36299 51665 36300
rect 50410 36179 50454 36299
rect 51454 36179 51789 36299
rect 53789 36179 53833 36299
rect 54679 36183 54750 36971
rect 55849 36844 56051 36971
rect 55849 36798 55961 36844
rect 56007 36798 56051 36844
rect 55849 36681 56051 36798
rect 55849 36635 55961 36681
rect 56007 36635 56051 36681
rect 55849 36517 56051 36635
rect 55849 36471 55961 36517
rect 56007 36471 56051 36517
rect 55849 36354 56051 36471
rect 55849 36308 55961 36354
rect 56007 36308 56051 36354
rect 55849 36183 56051 36308
<< polycontact >>
rect 29116 65598 29162 65644
rect 29116 65435 29162 65481
rect 29116 65271 29162 65317
rect 29116 65108 29162 65154
rect 42319 65797 42459 65843
rect 44067 65845 44113 65891
rect 38035 65505 38081 65645
rect 40694 65418 40740 65558
rect 44279 65458 44325 65598
rect 46967 65493 47013 65633
rect 29116 64698 29162 64744
rect 29116 64535 29162 64581
rect 29116 64371 29162 64417
rect 29116 64208 29162 64254
rect 33495 64362 33541 64784
rect 43373 64763 43513 64809
rect 40281 64691 40327 64737
rect 55961 65598 56007 65644
rect 55961 65435 56007 65481
rect 55961 65271 56007 65317
rect 55961 65108 56007 65154
rect 36475 64325 36521 64465
rect 36697 64325 36743 64465
rect 44358 64568 44498 64614
rect 38669 64327 38715 64467
rect 45464 64337 45604 64383
rect 48622 64352 48668 64492
rect 39844 64260 39890 64306
rect 51600 64332 51646 64754
rect 29116 63798 29162 63844
rect 29116 63635 29162 63681
rect 29116 63471 29162 63517
rect 29116 63308 29162 63354
rect 55961 64698 56007 64744
rect 55961 64535 56007 64581
rect 55961 64371 56007 64417
rect 55961 64208 56007 64254
rect 29116 62898 29162 62944
rect 29116 62735 29162 62781
rect 29116 62571 29162 62617
rect 29116 62408 29162 62454
rect 33495 63270 33541 63692
rect 36475 63589 36521 63729
rect 36697 63589 36743 63729
rect 38669 63587 38715 63727
rect 39844 63748 39890 63794
rect 45464 63671 45604 63717
rect 48622 63562 48668 63702
rect 44358 63440 44498 63486
rect 40281 63317 40327 63363
rect 33495 62562 33541 62984
rect 43373 63245 43513 63291
rect 51600 63300 51646 63722
rect 43373 62963 43513 63009
rect 40281 62891 40327 62937
rect 55961 63798 56007 63844
rect 55961 63635 56007 63681
rect 55961 63471 56007 63517
rect 55961 63308 56007 63354
rect 36475 62525 36521 62665
rect 36697 62525 36743 62665
rect 44358 62768 44498 62814
rect 38669 62527 38715 62667
rect 45464 62537 45604 62583
rect 48622 62552 48668 62692
rect 39844 62460 39890 62506
rect 51600 62532 51646 62954
rect 29116 61998 29162 62044
rect 29116 61835 29162 61881
rect 29116 61671 29162 61717
rect 29116 61508 29162 61554
rect 55961 62898 56007 62944
rect 55961 62735 56007 62781
rect 55961 62571 56007 62617
rect 55961 62408 56007 62454
rect 29116 61098 29162 61144
rect 29116 60935 29162 60981
rect 29116 60771 29162 60817
rect 29116 60608 29162 60654
rect 33495 61470 33541 61892
rect 36475 61789 36521 61929
rect 36697 61789 36743 61929
rect 38669 61787 38715 61927
rect 39844 61948 39890 61994
rect 45464 61871 45604 61917
rect 48622 61762 48668 61902
rect 44358 61640 44498 61686
rect 40281 61517 40327 61563
rect 33495 60762 33541 61184
rect 43373 61445 43513 61491
rect 51600 61500 51646 61922
rect 43373 61163 43513 61209
rect 40281 61091 40327 61137
rect 55961 61998 56007 62044
rect 55961 61835 56007 61881
rect 55961 61671 56007 61717
rect 55961 61508 56007 61554
rect 36475 60725 36521 60865
rect 36697 60725 36743 60865
rect 44358 60968 44498 61014
rect 38669 60727 38715 60867
rect 45464 60737 45604 60783
rect 48622 60752 48668 60892
rect 39844 60660 39890 60706
rect 51600 60732 51646 61154
rect 29116 60198 29162 60244
rect 29116 60035 29162 60081
rect 29116 59871 29162 59917
rect 29116 59708 29162 59754
rect 55961 61098 56007 61144
rect 55961 60935 56007 60981
rect 55961 60771 56007 60817
rect 55961 60608 56007 60654
rect 29116 59298 29162 59344
rect 29116 59135 29162 59181
rect 29116 58971 29162 59017
rect 29116 58808 29162 58854
rect 33495 59670 33541 60092
rect 36475 59989 36521 60129
rect 36697 59989 36743 60129
rect 38669 59987 38715 60127
rect 39844 60148 39890 60194
rect 45464 60071 45604 60117
rect 48622 59962 48668 60102
rect 44358 59840 44498 59886
rect 40281 59717 40327 59763
rect 33495 58962 33541 59384
rect 43373 59645 43513 59691
rect 51600 59700 51646 60122
rect 43373 59363 43513 59409
rect 40281 59291 40327 59337
rect 55961 60198 56007 60244
rect 55961 60035 56007 60081
rect 55961 59871 56007 59917
rect 55961 59708 56007 59754
rect 36475 58925 36521 59065
rect 36697 58925 36743 59065
rect 44358 59168 44498 59214
rect 38669 58927 38715 59067
rect 45464 58937 45604 58983
rect 48622 58952 48668 59092
rect 39844 58860 39890 58906
rect 51600 58932 51646 59354
rect 29116 58398 29162 58444
rect 29116 58235 29162 58281
rect 29116 58071 29162 58117
rect 29116 57908 29162 57954
rect 55961 59298 56007 59344
rect 55961 59135 56007 59181
rect 55961 58971 56007 59017
rect 55961 58808 56007 58854
rect 29116 57498 29162 57544
rect 29116 57335 29162 57381
rect 29116 57171 29162 57217
rect 29116 57008 29162 57054
rect 33495 57870 33541 58292
rect 36475 58189 36521 58329
rect 36697 58189 36743 58329
rect 38669 58187 38715 58327
rect 39844 58348 39890 58394
rect 45464 58271 45604 58317
rect 48622 58162 48668 58302
rect 44358 58040 44498 58086
rect 40281 57917 40327 57963
rect 33495 57162 33541 57584
rect 43373 57845 43513 57891
rect 51600 57900 51646 58322
rect 43373 57563 43513 57609
rect 40281 57491 40327 57537
rect 55961 58398 56007 58444
rect 55961 58235 56007 58281
rect 55961 58071 56007 58117
rect 55961 57908 56007 57954
rect 36475 57125 36521 57265
rect 36697 57125 36743 57265
rect 44358 57368 44498 57414
rect 38669 57127 38715 57267
rect 45464 57137 45604 57183
rect 48622 57152 48668 57292
rect 39844 57060 39890 57106
rect 51600 57132 51646 57554
rect 29116 56598 29162 56644
rect 29116 56435 29162 56481
rect 29116 56271 29162 56317
rect 29116 56108 29162 56154
rect 55961 57498 56007 57544
rect 55961 57335 56007 57381
rect 55961 57171 56007 57217
rect 55961 57008 56007 57054
rect 29116 55698 29162 55744
rect 29116 55535 29162 55581
rect 29116 55371 29162 55417
rect 29116 55208 29162 55254
rect 33495 56070 33541 56492
rect 36475 56389 36521 56529
rect 36697 56389 36743 56529
rect 38669 56387 38715 56527
rect 39844 56548 39890 56594
rect 45464 56471 45604 56517
rect 48622 56362 48668 56502
rect 44358 56240 44498 56286
rect 40281 56117 40327 56163
rect 33495 55362 33541 55784
rect 43373 56045 43513 56091
rect 51600 56100 51646 56522
rect 43373 55763 43513 55809
rect 40281 55691 40327 55737
rect 55961 56598 56007 56644
rect 55961 56435 56007 56481
rect 55961 56271 56007 56317
rect 55961 56108 56007 56154
rect 36475 55325 36521 55465
rect 36697 55325 36743 55465
rect 44358 55568 44498 55614
rect 38669 55327 38715 55467
rect 45464 55337 45604 55383
rect 48622 55352 48668 55492
rect 39844 55260 39890 55306
rect 51600 55332 51646 55754
rect 29116 54798 29162 54844
rect 29116 54635 29162 54681
rect 29116 54471 29162 54517
rect 29116 54308 29162 54354
rect 55961 55698 56007 55744
rect 55961 55535 56007 55581
rect 55961 55371 56007 55417
rect 55961 55208 56007 55254
rect 29116 53898 29162 53944
rect 29116 53735 29162 53781
rect 29116 53571 29162 53617
rect 29116 53408 29162 53454
rect 33495 54270 33541 54692
rect 36475 54589 36521 54729
rect 36697 54589 36743 54729
rect 38669 54587 38715 54727
rect 39844 54748 39890 54794
rect 45464 54671 45604 54717
rect 48622 54562 48668 54702
rect 44358 54440 44498 54486
rect 40281 54317 40327 54363
rect 33495 53562 33541 53984
rect 43373 54245 43513 54291
rect 51600 54300 51646 54722
rect 43373 53963 43513 54009
rect 40281 53891 40327 53937
rect 55961 54798 56007 54844
rect 55961 54635 56007 54681
rect 55961 54471 56007 54517
rect 55961 54308 56007 54354
rect 36475 53525 36521 53665
rect 36697 53525 36743 53665
rect 44358 53768 44498 53814
rect 38669 53527 38715 53667
rect 45464 53537 45604 53583
rect 48622 53552 48668 53692
rect 39844 53460 39890 53506
rect 51600 53532 51646 53954
rect 29116 52998 29162 53044
rect 29116 52835 29162 52881
rect 29116 52671 29162 52717
rect 29116 52508 29162 52554
rect 55961 53898 56007 53944
rect 55961 53735 56007 53781
rect 55961 53571 56007 53617
rect 55961 53408 56007 53454
rect 29116 52098 29162 52144
rect 29116 51935 29162 51981
rect 29116 51771 29162 51817
rect 29116 51608 29162 51654
rect 33495 52470 33541 52892
rect 36475 52789 36521 52929
rect 36697 52789 36743 52929
rect 38669 52787 38715 52927
rect 39844 52948 39890 52994
rect 45464 52871 45604 52917
rect 48622 52762 48668 52902
rect 44358 52640 44498 52686
rect 40281 52517 40327 52563
rect 33495 51762 33541 52184
rect 43373 52445 43513 52491
rect 51600 52500 51646 52922
rect 43373 52163 43513 52209
rect 40281 52091 40327 52137
rect 55961 52998 56007 53044
rect 55961 52835 56007 52881
rect 55961 52671 56007 52717
rect 55961 52508 56007 52554
rect 36475 51725 36521 51865
rect 36697 51725 36743 51865
rect 44358 51968 44498 52014
rect 38669 51727 38715 51867
rect 45464 51737 45604 51783
rect 48622 51752 48668 51892
rect 39844 51660 39890 51706
rect 51600 51732 51646 52154
rect 29116 51198 29162 51244
rect 29116 51035 29162 51081
rect 29116 50871 29162 50917
rect 29116 50708 29162 50754
rect 55961 52098 56007 52144
rect 55961 51935 56007 51981
rect 55961 51771 56007 51817
rect 55961 51608 56007 51654
rect 29116 50298 29162 50344
rect 29116 50135 29162 50181
rect 29116 49971 29162 50017
rect 29116 49808 29162 49854
rect 33495 50670 33541 51092
rect 36475 50989 36521 51129
rect 36697 50989 36743 51129
rect 38669 50987 38715 51127
rect 39844 51148 39890 51194
rect 45464 51071 45604 51117
rect 48622 50962 48668 51102
rect 44358 50840 44498 50886
rect 40281 50717 40327 50763
rect 33495 49962 33541 50384
rect 43373 50645 43513 50691
rect 51600 50700 51646 51122
rect 43373 50363 43513 50409
rect 40281 50291 40327 50337
rect 55961 51198 56007 51244
rect 55961 51035 56007 51081
rect 55961 50871 56007 50917
rect 55961 50708 56007 50754
rect 36475 49925 36521 50065
rect 36697 49925 36743 50065
rect 44358 50168 44498 50214
rect 38669 49927 38715 50067
rect 45464 49937 45604 49983
rect 48622 49952 48668 50092
rect 39844 49860 39890 49906
rect 51600 49932 51646 50354
rect 29116 49398 29162 49444
rect 29116 49235 29162 49281
rect 29116 49071 29162 49117
rect 29116 48908 29162 48954
rect 55961 50298 56007 50344
rect 55961 50135 56007 50181
rect 55961 49971 56007 50017
rect 55961 49808 56007 49854
rect 29116 48498 29162 48544
rect 29116 48335 29162 48381
rect 29116 48171 29162 48217
rect 29116 48008 29162 48054
rect 33495 48870 33541 49292
rect 36475 49189 36521 49329
rect 36697 49189 36743 49329
rect 38669 49187 38715 49327
rect 39844 49348 39890 49394
rect 45464 49271 45604 49317
rect 48622 49162 48668 49302
rect 44358 49040 44498 49086
rect 40281 48917 40327 48963
rect 33495 48162 33541 48584
rect 43373 48845 43513 48891
rect 51600 48900 51646 49322
rect 43373 48563 43513 48609
rect 40281 48491 40327 48537
rect 55961 49398 56007 49444
rect 55961 49235 56007 49281
rect 55961 49071 56007 49117
rect 55961 48908 56007 48954
rect 36475 48125 36521 48265
rect 36697 48125 36743 48265
rect 44358 48368 44498 48414
rect 38669 48127 38715 48267
rect 45464 48137 45604 48183
rect 48622 48152 48668 48292
rect 39844 48060 39890 48106
rect 51600 48132 51646 48554
rect 29116 47598 29162 47644
rect 29116 47435 29162 47481
rect 29116 47271 29162 47317
rect 29116 47108 29162 47154
rect 55961 48498 56007 48544
rect 55961 48335 56007 48381
rect 55961 48171 56007 48217
rect 55961 48008 56007 48054
rect 29116 46698 29162 46744
rect 29116 46535 29162 46581
rect 29116 46371 29162 46417
rect 29116 46208 29162 46254
rect 33495 47070 33541 47492
rect 36475 47389 36521 47529
rect 36697 47389 36743 47529
rect 38669 47387 38715 47527
rect 39844 47548 39890 47594
rect 45464 47471 45604 47517
rect 48622 47362 48668 47502
rect 44358 47240 44498 47286
rect 40281 47117 40327 47163
rect 33495 46362 33541 46784
rect 43373 47045 43513 47091
rect 51600 47100 51646 47522
rect 43373 46763 43513 46809
rect 40281 46691 40327 46737
rect 55961 47598 56007 47644
rect 55961 47435 56007 47481
rect 55961 47271 56007 47317
rect 55961 47108 56007 47154
rect 36475 46325 36521 46465
rect 36697 46325 36743 46465
rect 44358 46568 44498 46614
rect 38669 46327 38715 46467
rect 45464 46337 45604 46383
rect 48622 46352 48668 46492
rect 39844 46260 39890 46306
rect 51600 46332 51646 46754
rect 29116 45798 29162 45844
rect 29116 45635 29162 45681
rect 29116 45471 29162 45517
rect 29116 45308 29162 45354
rect 55961 46698 56007 46744
rect 55961 46535 56007 46581
rect 55961 46371 56007 46417
rect 55961 46208 56007 46254
rect 29116 44898 29162 44944
rect 29116 44735 29162 44781
rect 29116 44571 29162 44617
rect 29116 44408 29162 44454
rect 33495 45270 33541 45692
rect 36475 45589 36521 45729
rect 36697 45589 36743 45729
rect 38669 45587 38715 45727
rect 39844 45748 39890 45794
rect 45464 45671 45604 45717
rect 48622 45562 48668 45702
rect 44358 45440 44498 45486
rect 40281 45317 40327 45363
rect 33495 44562 33541 44984
rect 43373 45245 43513 45291
rect 51600 45300 51646 45722
rect 43373 44963 43513 45009
rect 40281 44891 40327 44937
rect 55961 45798 56007 45844
rect 55961 45635 56007 45681
rect 55961 45471 56007 45517
rect 55961 45308 56007 45354
rect 36475 44525 36521 44665
rect 36697 44525 36743 44665
rect 44358 44768 44498 44814
rect 38669 44527 38715 44667
rect 45464 44537 45604 44583
rect 48622 44552 48668 44692
rect 39844 44460 39890 44506
rect 51600 44532 51646 44954
rect 29116 43998 29162 44044
rect 29116 43835 29162 43881
rect 29116 43671 29162 43717
rect 29116 43508 29162 43554
rect 55961 44898 56007 44944
rect 55961 44735 56007 44781
rect 55961 44571 56007 44617
rect 55961 44408 56007 44454
rect 29116 43098 29162 43144
rect 29116 42935 29162 42981
rect 29116 42771 29162 42817
rect 29116 42608 29162 42654
rect 33495 43470 33541 43892
rect 36475 43789 36521 43929
rect 36697 43789 36743 43929
rect 38669 43787 38715 43927
rect 39844 43948 39890 43994
rect 45464 43871 45604 43917
rect 48622 43762 48668 43902
rect 44358 43640 44498 43686
rect 40281 43517 40327 43563
rect 33495 42762 33541 43184
rect 43373 43445 43513 43491
rect 51600 43500 51646 43922
rect 43373 43163 43513 43209
rect 40281 43091 40327 43137
rect 55961 43998 56007 44044
rect 55961 43835 56007 43881
rect 55961 43671 56007 43717
rect 55961 43508 56007 43554
rect 36475 42725 36521 42865
rect 36697 42725 36743 42865
rect 44358 42968 44498 43014
rect 38669 42727 38715 42867
rect 45464 42737 45604 42783
rect 48622 42752 48668 42892
rect 39844 42660 39890 42706
rect 51600 42732 51646 43154
rect 29116 42198 29162 42244
rect 29116 42035 29162 42081
rect 29116 41871 29162 41917
rect 29116 41708 29162 41754
rect 55961 43098 56007 43144
rect 55961 42935 56007 42981
rect 55961 42771 56007 42817
rect 55961 42608 56007 42654
rect 29116 41298 29162 41344
rect 29116 41135 29162 41181
rect 29116 40971 29162 41017
rect 29116 40808 29162 40854
rect 33495 41670 33541 42092
rect 36475 41989 36521 42129
rect 36697 41989 36743 42129
rect 38669 41987 38715 42127
rect 39844 42148 39890 42194
rect 45464 42071 45604 42117
rect 48622 41962 48668 42102
rect 44358 41840 44498 41886
rect 40281 41717 40327 41763
rect 33495 40962 33541 41384
rect 43373 41645 43513 41691
rect 51600 41700 51646 42122
rect 43373 41363 43513 41409
rect 40281 41291 40327 41337
rect 55961 42198 56007 42244
rect 55961 42035 56007 42081
rect 55961 41871 56007 41917
rect 55961 41708 56007 41754
rect 36475 40925 36521 41065
rect 36697 40925 36743 41065
rect 44358 41168 44498 41214
rect 38669 40927 38715 41067
rect 45464 40937 45604 40983
rect 48622 40952 48668 41092
rect 39844 40860 39890 40906
rect 51600 40932 51646 41354
rect 29116 40398 29162 40444
rect 29116 40235 29162 40281
rect 29116 40071 29162 40117
rect 29116 39908 29162 39954
rect 55961 41298 56007 41344
rect 55961 41135 56007 41181
rect 55961 40971 56007 41017
rect 55961 40808 56007 40854
rect 29116 39498 29162 39544
rect 29116 39335 29162 39381
rect 29116 39171 29162 39217
rect 29116 39008 29162 39054
rect 33495 39870 33541 40292
rect 36475 40189 36521 40329
rect 36697 40189 36743 40329
rect 38669 40187 38715 40327
rect 39844 40348 39890 40394
rect 45464 40271 45604 40317
rect 48622 40162 48668 40302
rect 44358 40040 44498 40086
rect 40281 39917 40327 39963
rect 33495 39162 33541 39584
rect 43373 39845 43513 39891
rect 51600 39900 51646 40322
rect 43373 39563 43513 39609
rect 40281 39491 40327 39537
rect 55961 40398 56007 40444
rect 55961 40235 56007 40281
rect 55961 40071 56007 40117
rect 55961 39908 56007 39954
rect 36475 39125 36521 39265
rect 36697 39125 36743 39265
rect 44358 39368 44498 39414
rect 38669 39127 38715 39267
rect 45464 39137 45604 39183
rect 48622 39152 48668 39292
rect 39844 39060 39890 39106
rect 51600 39132 51646 39554
rect 29116 38598 29162 38644
rect 29116 38435 29162 38481
rect 29116 38271 29162 38317
rect 29116 38108 29162 38154
rect 55961 39498 56007 39544
rect 55961 39335 56007 39381
rect 55961 39171 56007 39217
rect 55961 39008 56007 39054
rect 29116 37698 29162 37744
rect 29116 37535 29162 37581
rect 29116 37371 29162 37417
rect 29116 37208 29162 37254
rect 33495 38070 33541 38492
rect 36475 38389 36521 38529
rect 36697 38389 36743 38529
rect 38669 38387 38715 38527
rect 39844 38548 39890 38594
rect 45464 38471 45604 38517
rect 48622 38362 48668 38502
rect 44358 38240 44498 38286
rect 40281 38117 40327 38163
rect 33495 37362 33541 37784
rect 43373 38045 43513 38091
rect 51600 38100 51646 38522
rect 43373 37763 43513 37809
rect 40281 37691 40327 37737
rect 55961 38598 56007 38644
rect 55961 38435 56007 38481
rect 55961 38271 56007 38317
rect 55961 38108 56007 38154
rect 36475 37325 36521 37465
rect 36697 37325 36743 37465
rect 44358 37568 44498 37614
rect 38669 37327 38715 37467
rect 45464 37337 45604 37383
rect 48622 37352 48668 37492
rect 39844 37260 39890 37306
rect 51600 37332 51646 37754
rect 29116 36798 29162 36844
rect 29116 36635 29162 36681
rect 29116 36471 29162 36517
rect 29116 36308 29162 36354
rect 55961 37698 56007 37744
rect 55961 37535 56007 37581
rect 55961 37371 56007 37417
rect 55961 37208 56007 37254
rect 33495 36270 33541 36692
rect 36475 36589 36521 36729
rect 36697 36589 36743 36729
rect 38669 36587 38715 36727
rect 39844 36748 39890 36794
rect 45464 36671 45604 36717
rect 48622 36562 48668 36702
rect 44358 36440 44498 36486
rect 40281 36317 40327 36363
rect 43373 36245 43513 36291
rect 51600 36300 51646 36722
rect 55961 36798 56007 36844
rect 55961 36635 56007 36681
rect 55961 36471 56007 36517
rect 55961 36308 56007 36354
<< metal1 >>
rect 282 66894 86090 67894
rect 25313 65914 26039 66894
rect 25313 65862 25380 65914
rect 25432 65862 25504 65914
rect 25556 65862 25628 65914
rect 25680 65862 25752 65914
rect 25804 65862 25876 65914
rect 25928 65862 26039 65914
rect 25313 65790 26039 65862
rect 25313 65738 25380 65790
rect 25432 65738 25504 65790
rect 25556 65738 25628 65790
rect 25680 65738 25752 65790
rect 25804 65738 25876 65790
rect 25928 65738 26039 65790
rect 25313 65678 26039 65738
rect 27387 65853 29196 66894
rect 33544 65966 34341 66894
rect 33001 65909 35013 65966
rect 27387 65801 27790 65853
rect 27842 65801 28001 65853
rect 28053 65801 28212 65853
rect 28264 65801 28423 65853
rect 28475 65801 28634 65853
rect 28686 65801 28845 65853
rect 28897 65801 29056 65853
rect 29108 65801 29196 65853
rect 27387 65722 29196 65801
rect 29283 65853 30365 65894
rect 29283 65850 29582 65853
rect 29283 65804 29317 65850
rect 29363 65804 29478 65850
rect 29524 65804 29582 65850
rect 29283 65801 29582 65804
rect 29634 65850 29793 65853
rect 29845 65850 30005 65853
rect 29634 65804 29638 65850
rect 29684 65804 29793 65850
rect 29845 65804 29959 65850
rect 29634 65801 29793 65804
rect 29845 65801 30005 65804
rect 30057 65850 30216 65853
rect 30057 65804 30121 65850
rect 30167 65804 30216 65850
rect 30057 65801 30216 65804
rect 30268 65850 30365 65853
rect 30268 65804 30284 65850
rect 30330 65804 30365 65850
rect 30268 65801 30365 65804
rect 29283 65761 30365 65801
rect 30583 65853 32694 65894
rect 30583 65801 30807 65853
rect 30859 65836 31018 65853
rect 31070 65836 31229 65853
rect 30583 65790 30854 65801
rect 30900 65790 31012 65836
rect 31070 65801 31170 65836
rect 31058 65790 31170 65801
rect 31216 65801 31229 65836
rect 31281 65836 31440 65853
rect 31492 65836 31651 65853
rect 31703 65836 31861 65853
rect 31281 65801 31328 65836
rect 31216 65790 31328 65801
rect 31374 65801 31440 65836
rect 31374 65790 31487 65801
rect 31533 65790 31645 65836
rect 31703 65801 31803 65836
rect 31691 65790 31803 65801
rect 31849 65801 31861 65836
rect 31913 65836 32072 65853
rect 32124 65836 32283 65853
rect 32335 65836 32494 65853
rect 31913 65801 31961 65836
rect 31849 65790 31961 65801
rect 32007 65801 32072 65836
rect 32007 65790 32119 65801
rect 32165 65790 32277 65836
rect 32335 65801 32435 65836
rect 32323 65790 32435 65801
rect 32481 65801 32494 65836
rect 32546 65836 32694 65853
rect 32546 65801 32593 65836
rect 32481 65790 32593 65801
rect 32639 65790 32694 65836
rect 29544 65760 30306 65761
rect 27387 65676 28810 65722
rect 28856 65676 29196 65722
rect 27387 65644 29196 65676
rect 27387 65598 29116 65644
rect 29162 65598 29196 65644
rect 27387 65558 29196 65598
rect 27387 65512 28810 65558
rect 28856 65512 29196 65558
rect 27387 65481 29196 65512
rect 27387 65435 29116 65481
rect 29162 65435 29196 65481
rect 27387 65395 29196 65435
rect 27387 65349 28810 65395
rect 28856 65349 29196 65395
rect 27387 65317 29196 65349
rect 27387 65271 29116 65317
rect 29162 65271 29196 65317
rect 27387 65232 29196 65271
rect 27387 65186 28810 65232
rect 28856 65186 29196 65232
rect 27387 65154 29196 65186
rect 27387 65108 29116 65154
rect 29162 65108 29196 65154
rect 27387 65068 29196 65108
rect 27387 65022 28810 65068
rect 28856 65022 29196 65068
rect 27387 64866 29196 65022
rect 30583 65722 32694 65790
rect 30583 65676 30637 65722
rect 30683 65676 32694 65722
rect 30583 65673 32694 65676
rect 30583 65635 30854 65673
rect 30583 65583 30807 65635
rect 30900 65627 31012 65673
rect 31058 65635 31170 65673
rect 31070 65627 31170 65635
rect 31216 65635 31328 65673
rect 31216 65627 31229 65635
rect 30859 65583 31018 65627
rect 31070 65583 31229 65627
rect 31281 65627 31328 65635
rect 31374 65635 31487 65673
rect 31374 65627 31440 65635
rect 31533 65627 31645 65673
rect 31691 65635 31803 65673
rect 31703 65627 31803 65635
rect 31849 65635 31961 65673
rect 31849 65627 31861 65635
rect 31281 65583 31440 65627
rect 31492 65583 31651 65627
rect 31703 65583 31861 65627
rect 31913 65627 31961 65635
rect 32007 65635 32119 65673
rect 32007 65627 32072 65635
rect 32165 65627 32277 65673
rect 32323 65635 32435 65673
rect 32335 65627 32435 65635
rect 32481 65635 32593 65673
rect 32481 65627 32494 65635
rect 31913 65583 32072 65627
rect 32124 65583 32283 65627
rect 32335 65583 32494 65627
rect 32546 65627 32593 65635
rect 32639 65627 32694 65673
rect 32546 65583 32694 65627
rect 30583 65558 32694 65583
rect 30583 65512 30637 65558
rect 30683 65512 32694 65558
rect 33001 65863 33044 65909
rect 33090 65863 33202 65909
rect 33248 65863 33360 65909
rect 33406 65863 33518 65909
rect 33564 65863 33677 65909
rect 33723 65863 33835 65909
rect 33881 65863 33993 65909
rect 34039 65863 34151 65909
rect 34197 65863 34309 65909
rect 34355 65863 34467 65909
rect 34513 65863 34625 65909
rect 34671 65863 34783 65909
rect 34829 65863 35013 65909
rect 40062 65946 40923 66894
rect 43738 65946 44599 66894
rect 50001 65946 50913 66894
rect 40062 65909 41937 65946
rect 33001 65853 35013 65863
rect 33001 65801 34290 65853
rect 34342 65801 34501 65853
rect 34553 65801 34712 65853
rect 34764 65801 34923 65853
rect 34975 65801 35013 65853
rect 35405 65833 36377 65873
rect 35405 65818 35443 65833
rect 35495 65818 35654 65833
rect 35706 65818 35865 65833
rect 35917 65818 36076 65833
rect 36128 65818 36287 65833
rect 36339 65818 36377 65833
rect 40062 65863 40117 65909
rect 40163 65863 40275 65909
rect 40321 65863 40433 65909
rect 40479 65863 40591 65909
rect 40637 65863 40750 65909
rect 40796 65863 40908 65909
rect 40954 65863 41066 65909
rect 41112 65863 41224 65909
rect 41270 65863 41382 65909
rect 41428 65863 41540 65909
rect 41586 65863 41698 65909
rect 41744 65863 41856 65909
rect 41902 65863 41937 65909
rect 40062 65858 41937 65863
rect 33001 65635 35013 65801
rect 35396 65772 35409 65818
rect 37291 65772 37348 65818
rect 37394 65772 37451 65818
rect 37497 65772 37554 65818
rect 37600 65772 37657 65818
rect 37703 65772 37760 65818
rect 37806 65772 37863 65818
rect 37909 65772 37922 65818
rect 40062 65806 40252 65858
rect 40304 65806 40432 65858
rect 40484 65826 41937 65858
rect 42208 65909 43589 65946
rect 42208 65905 42717 65909
rect 42208 65853 42710 65905
rect 42763 65863 42875 65909
rect 42921 65905 43033 65909
rect 42762 65853 42921 65863
rect 42973 65863 43033 65905
rect 43079 65905 43191 65909
rect 43079 65863 43132 65905
rect 42973 65853 43132 65863
rect 43184 65863 43191 65905
rect 43237 65863 43350 65909
rect 43396 65863 43508 65909
rect 43554 65863 43589 65909
rect 43184 65853 43589 65863
rect 42208 65844 43589 65853
rect 40484 65806 40590 65826
rect 35405 65741 36377 65772
rect 38000 65645 38116 65712
rect 33001 65594 34290 65635
rect 33001 65548 33014 65594
rect 33774 65548 33831 65594
rect 33877 65548 33934 65594
rect 33980 65548 34037 65594
rect 34083 65548 34140 65594
rect 34186 65548 34243 65594
rect 34289 65583 34290 65594
rect 34342 65594 34501 65635
rect 34553 65594 34712 65635
rect 34764 65594 34923 65635
rect 34975 65594 35013 65635
rect 35159 65594 35444 65635
rect 34342 65583 34346 65594
rect 34289 65548 34346 65583
rect 34392 65548 34449 65594
rect 34495 65583 34501 65594
rect 34495 65548 34552 65583
rect 34598 65548 34655 65594
rect 34701 65583 34712 65594
rect 34701 65548 34758 65583
rect 34804 65548 34861 65594
rect 34907 65583 34923 65594
rect 34907 65548 34964 65583
rect 35010 65548 35023 65594
rect 35159 65548 35409 65594
rect 37291 65548 37348 65594
rect 37394 65548 37451 65594
rect 37497 65548 37554 65594
rect 37600 65548 37657 65594
rect 37703 65548 37760 65594
rect 37806 65548 37863 65594
rect 37909 65548 37922 65594
rect 34251 65543 35013 65548
rect 30583 65509 32694 65512
rect 30583 65463 30854 65509
rect 30900 65463 31012 65509
rect 31058 65463 31170 65509
rect 31216 65463 31328 65509
rect 31374 65463 31487 65509
rect 31533 65463 31645 65509
rect 31691 65463 31803 65509
rect 31849 65463 31961 65509
rect 32007 65463 32119 65509
rect 32165 65463 32277 65509
rect 32323 65463 32435 65509
rect 32481 65463 32593 65509
rect 32639 65463 32694 65509
rect 30583 65418 32694 65463
rect 30583 65395 30807 65418
rect 30583 65349 30637 65395
rect 30683 65366 30807 65395
rect 30859 65366 31018 65418
rect 31070 65366 31229 65418
rect 31281 65366 31440 65418
rect 31492 65366 31651 65418
rect 31703 65366 31861 65418
rect 31913 65366 32072 65418
rect 32124 65366 32283 65418
rect 32335 65366 32494 65418
rect 32546 65366 32694 65418
rect 35159 65515 35444 65548
rect 33012 65372 33984 65412
rect 35159 65404 35275 65515
rect 38000 65505 38035 65645
rect 38081 65505 38116 65645
rect 39015 65635 39565 65642
rect 39014 65601 39565 65635
rect 39014 65594 39053 65601
rect 39105 65594 39264 65601
rect 39316 65594 39475 65601
rect 39527 65594 39565 65601
rect 40062 65640 40590 65806
rect 42208 65792 42246 65844
rect 42298 65843 42458 65844
rect 42298 65797 42319 65843
rect 42510 65826 43589 65844
rect 43738 65909 44960 65946
rect 43738 65905 44514 65909
rect 43738 65853 43777 65905
rect 43829 65853 43988 65905
rect 44040 65891 44199 65905
rect 44040 65853 44067 65891
rect 43738 65845 44067 65853
rect 44113 65853 44199 65891
rect 44251 65853 44410 65905
rect 44462 65863 44514 65905
rect 44560 65863 44672 65909
rect 44718 65863 44830 65909
rect 44876 65863 44960 65909
rect 50001 65909 52023 65946
rect 48789 65867 49551 65873
rect 44462 65853 44960 65863
rect 44113 65845 44960 65853
rect 42510 65813 43222 65826
rect 42510 65812 42717 65813
rect 43738 65812 44960 65845
rect 42298 65792 42458 65797
rect 42510 65792 42548 65812
rect 42208 65751 42548 65792
rect 40062 65594 40252 65640
rect 40304 65594 40432 65640
rect 40484 65594 40590 65640
rect 44268 65598 44336 65609
rect 38363 65548 38376 65594
rect 38422 65548 38479 65594
rect 38525 65548 38582 65594
rect 38628 65548 38686 65594
rect 38732 65548 38790 65594
rect 38836 65548 38894 65594
rect 38940 65548 38998 65594
rect 39044 65549 39053 65594
rect 39044 65548 39102 65549
rect 39148 65548 39206 65594
rect 39252 65549 39264 65594
rect 39252 65548 39310 65549
rect 39356 65548 39414 65594
rect 39460 65549 39475 65594
rect 39460 65548 39518 65549
rect 39564 65548 39622 65594
rect 39668 65548 39681 65594
rect 40062 65548 40075 65594
rect 40121 65548 40189 65594
rect 40235 65588 40252 65594
rect 40235 65548 40303 65588
rect 40349 65548 40417 65594
rect 40484 65588 40531 65594
rect 40463 65548 40531 65588
rect 40577 65548 40590 65594
rect 40683 65558 40976 65595
rect 39014 65515 39565 65548
rect 39015 65509 39565 65515
rect 33012 65370 33050 65372
rect 33102 65370 33261 65372
rect 33313 65370 33472 65372
rect 33524 65370 33683 65372
rect 33735 65370 33894 65372
rect 33946 65370 33984 65372
rect 34917 65370 35275 65404
rect 35405 65370 36377 65410
rect 38000 65404 38116 65505
rect 40683 65418 40694 65558
rect 40740 65549 40976 65558
rect 41022 65549 41079 65595
rect 41125 65549 41182 65595
rect 41228 65549 41286 65595
rect 41332 65549 41390 65595
rect 41436 65549 41494 65595
rect 41540 65549 41598 65595
rect 41644 65549 41702 65595
rect 41748 65549 41806 65595
rect 41852 65549 41910 65595
rect 41956 65549 42014 65595
rect 42060 65549 42118 65595
rect 42164 65549 42222 65595
rect 42268 65594 42851 65595
rect 44268 65594 44279 65598
rect 42268 65549 42676 65594
rect 40740 65418 40751 65549
rect 42663 65548 42676 65549
rect 42722 65548 42779 65594
rect 42825 65548 42882 65594
rect 42928 65548 42986 65594
rect 43032 65548 43090 65594
rect 43136 65548 43194 65594
rect 43240 65548 43298 65594
rect 43344 65548 43402 65594
rect 43448 65548 43506 65594
rect 43552 65548 43610 65594
rect 43656 65548 43714 65594
rect 43760 65548 43818 65594
rect 43864 65548 43922 65594
rect 43968 65548 44279 65594
rect 44268 65458 44279 65548
rect 44325 65458 44336 65598
rect 44432 65594 44960 65812
rect 44432 65548 44445 65594
rect 44491 65548 44559 65594
rect 44605 65548 44673 65594
rect 44719 65548 44787 65594
rect 44833 65548 44901 65594
rect 44947 65548 44960 65594
rect 45333 65833 49619 65867
rect 45333 65818 48828 65833
rect 48880 65818 49039 65833
rect 49091 65818 49250 65833
rect 49302 65818 49461 65833
rect 49513 65818 49619 65833
rect 50001 65863 50129 65909
rect 50175 65863 50287 65909
rect 50333 65863 50445 65909
rect 50491 65863 50603 65909
rect 50649 65863 50762 65909
rect 50808 65863 50920 65909
rect 50966 65863 51078 65909
rect 51124 65863 51236 65909
rect 51282 65863 51394 65909
rect 51440 65863 51552 65909
rect 51598 65863 51710 65909
rect 51756 65863 51868 65909
rect 51914 65863 52023 65909
rect 50001 65853 52023 65863
rect 45333 65772 47114 65818
rect 48996 65781 49039 65818
rect 48996 65772 49053 65781
rect 49099 65772 49156 65818
rect 49202 65781 49250 65818
rect 49202 65772 49259 65781
rect 49305 65772 49362 65818
rect 49408 65781 49461 65818
rect 49513 65781 49568 65818
rect 49408 65772 49465 65781
rect 49511 65772 49568 65781
rect 49614 65772 49627 65818
rect 50001 65801 50137 65853
rect 50189 65801 50348 65853
rect 50400 65801 50559 65853
rect 50611 65801 50770 65853
rect 50822 65801 52023 65853
rect 45333 65747 49619 65772
rect 45333 65594 46651 65747
rect 48789 65740 49551 65747
rect 45333 65548 45346 65594
rect 45392 65548 45449 65594
rect 45495 65548 45552 65594
rect 45598 65548 45656 65594
rect 45702 65548 45760 65594
rect 45806 65548 45864 65594
rect 45910 65548 45968 65594
rect 46014 65548 46072 65594
rect 46118 65548 46176 65594
rect 46222 65548 46280 65594
rect 46326 65548 46384 65594
rect 46430 65548 46488 65594
rect 46534 65548 46592 65594
rect 46638 65548 46651 65594
rect 46956 65633 47024 65644
rect 44432 65515 44960 65548
rect 44268 65447 44336 65458
rect 46956 65493 46967 65633
rect 47013 65493 47024 65633
rect 50001 65635 52023 65801
rect 50001 65594 50137 65635
rect 50189 65594 50348 65635
rect 50400 65594 50559 65635
rect 50611 65594 50770 65635
rect 50822 65594 52023 65635
rect 47101 65548 47114 65594
rect 48996 65548 49053 65594
rect 49099 65548 49156 65594
rect 49202 65548 49259 65594
rect 49305 65548 49362 65594
rect 49408 65548 49465 65594
rect 49511 65548 49568 65594
rect 49614 65548 49861 65594
rect 46956 65482 47024 65493
rect 40683 65407 40751 65418
rect 38000 65370 40590 65404
rect 40971 65371 42155 65411
rect 46956 65404 47023 65482
rect 30683 65349 32694 65366
rect 30583 65346 32694 65349
rect 30583 65300 30854 65346
rect 30900 65300 31012 65346
rect 31058 65300 31170 65346
rect 31216 65300 31328 65346
rect 31374 65300 31487 65346
rect 31533 65300 31645 65346
rect 31691 65300 31803 65346
rect 31849 65300 31961 65346
rect 32007 65300 32119 65346
rect 32165 65300 32277 65346
rect 32323 65300 32435 65346
rect 32481 65300 32593 65346
rect 32639 65300 32694 65346
rect 33001 65324 33014 65370
rect 33774 65324 33831 65370
rect 33877 65324 33894 65370
rect 33980 65324 34037 65370
rect 34083 65324 34140 65370
rect 34186 65324 34243 65370
rect 34289 65324 34346 65370
rect 34392 65324 34449 65370
rect 34495 65324 34552 65370
rect 34598 65324 34655 65370
rect 34701 65324 34758 65370
rect 34804 65324 34861 65370
rect 34907 65324 34964 65370
rect 35010 65324 35275 65370
rect 35396 65324 35409 65370
rect 37291 65324 37348 65370
rect 37394 65324 37451 65370
rect 37497 65324 37554 65370
rect 37600 65324 37657 65370
rect 37703 65324 37760 65370
rect 37806 65324 37863 65370
rect 37909 65324 37922 65370
rect 38000 65324 38376 65370
rect 38422 65324 38479 65370
rect 38525 65324 38582 65370
rect 38628 65324 38686 65370
rect 38732 65324 38790 65370
rect 38836 65324 38894 65370
rect 38940 65324 38998 65370
rect 39044 65324 39102 65370
rect 39148 65324 39206 65370
rect 39252 65324 39310 65370
rect 39356 65324 39414 65370
rect 39460 65324 39518 65370
rect 39564 65324 39622 65370
rect 39668 65324 40075 65370
rect 40121 65324 40189 65370
rect 40235 65324 40303 65370
rect 40349 65324 40417 65370
rect 40463 65324 40531 65370
rect 40577 65324 40590 65370
rect 40963 65325 40976 65371
rect 41022 65370 41079 65371
rect 41062 65325 41079 65370
rect 41125 65325 41182 65371
rect 41228 65370 41286 65371
rect 41273 65325 41286 65370
rect 41332 65325 41390 65371
rect 41436 65370 41494 65371
rect 41484 65325 41494 65370
rect 41540 65325 41598 65371
rect 41644 65370 41702 65371
rect 41695 65325 41702 65370
rect 41748 65325 41806 65371
rect 41852 65370 41910 65371
rect 41852 65325 41854 65370
rect 30583 65243 32694 65300
rect 33012 65320 33050 65324
rect 33102 65320 33261 65324
rect 33313 65320 33472 65324
rect 33524 65320 33683 65324
rect 33735 65320 33894 65324
rect 33946 65320 33984 65324
rect 33012 65280 33984 65320
rect 34917 65284 35275 65324
rect 35405 65318 35443 65324
rect 35495 65318 35654 65324
rect 35706 65318 35865 65324
rect 35917 65318 36076 65324
rect 36128 65318 36287 65324
rect 36339 65318 36377 65324
rect 35405 65278 36377 65318
rect 38000 65284 40590 65324
rect 40971 65318 41010 65325
rect 41062 65318 41221 65325
rect 41273 65318 41432 65325
rect 41484 65318 41643 65325
rect 41695 65318 41854 65325
rect 41906 65325 41910 65370
rect 41956 65325 42014 65371
rect 42060 65370 42118 65371
rect 42060 65325 42064 65370
rect 41906 65318 42064 65325
rect 42116 65325 42118 65370
rect 42164 65325 42222 65371
rect 42268 65370 42851 65371
rect 44432 65370 47023 65404
rect 48789 65370 49551 65410
rect 49744 65370 49861 65548
rect 50001 65548 50014 65594
rect 50822 65583 50831 65594
rect 50774 65548 50831 65583
rect 50877 65548 50934 65594
rect 50980 65548 51037 65594
rect 51083 65548 51140 65594
rect 51186 65548 51243 65594
rect 51289 65548 51346 65594
rect 51392 65548 51449 65594
rect 51495 65548 51552 65594
rect 51598 65548 51655 65594
rect 51701 65548 51758 65594
rect 51804 65548 51861 65594
rect 51907 65548 51964 65594
rect 52010 65548 52023 65594
rect 50001 65529 52023 65548
rect 52428 65853 54540 65894
rect 52428 65836 52576 65853
rect 52428 65790 52483 65836
rect 52529 65801 52576 65836
rect 52628 65836 52787 65853
rect 52839 65836 52998 65853
rect 53050 65836 53209 65853
rect 52628 65801 52641 65836
rect 52529 65790 52641 65801
rect 52687 65801 52787 65836
rect 52687 65790 52799 65801
rect 52845 65790 52957 65836
rect 53050 65801 53115 65836
rect 53003 65790 53115 65801
rect 53161 65801 53209 65836
rect 53261 65836 53419 65853
rect 53471 65836 53630 65853
rect 53682 65836 53841 65853
rect 53261 65801 53273 65836
rect 53161 65790 53273 65801
rect 53319 65801 53419 65836
rect 53319 65790 53431 65801
rect 53477 65790 53589 65836
rect 53682 65801 53748 65836
rect 53635 65790 53748 65801
rect 53794 65801 53841 65836
rect 53893 65836 54052 65853
rect 54104 65836 54263 65853
rect 53893 65801 53906 65836
rect 53794 65790 53906 65801
rect 53952 65801 54052 65836
rect 53952 65790 54064 65801
rect 54110 65790 54222 65836
rect 54315 65801 54540 65853
rect 54268 65790 54540 65801
rect 52428 65722 54540 65790
rect 54758 65853 55840 65894
rect 54758 65850 54855 65853
rect 54758 65804 54793 65850
rect 54839 65804 54855 65850
rect 54758 65801 54855 65804
rect 54907 65850 55066 65853
rect 54907 65804 54956 65850
rect 55002 65804 55066 65850
rect 54907 65801 55066 65804
rect 55118 65850 55278 65853
rect 55330 65850 55489 65853
rect 55164 65804 55278 65850
rect 55330 65804 55439 65850
rect 55485 65804 55489 65850
rect 55118 65801 55278 65804
rect 55330 65801 55489 65804
rect 55541 65850 55840 65853
rect 55541 65804 55599 65850
rect 55645 65804 55760 65850
rect 55806 65804 55840 65850
rect 55541 65801 55840 65804
rect 54758 65761 55840 65801
rect 55927 65853 57736 66894
rect 55927 65801 56015 65853
rect 56067 65801 56226 65853
rect 56278 65801 56437 65853
rect 56489 65801 56648 65853
rect 56700 65801 56859 65853
rect 56911 65801 57070 65853
rect 57122 65801 57281 65853
rect 57333 65801 57736 65853
rect 54817 65760 55579 65761
rect 52428 65676 54440 65722
rect 54486 65676 54540 65722
rect 52428 65673 54540 65676
rect 52428 65627 52483 65673
rect 52529 65635 52641 65673
rect 52529 65627 52576 65635
rect 52428 65583 52576 65627
rect 52628 65627 52641 65635
rect 52687 65635 52799 65673
rect 52687 65627 52787 65635
rect 52845 65627 52957 65673
rect 53003 65635 53115 65673
rect 53050 65627 53115 65635
rect 53161 65635 53273 65673
rect 53161 65627 53209 65635
rect 52628 65583 52787 65627
rect 52839 65583 52998 65627
rect 53050 65583 53209 65627
rect 53261 65627 53273 65635
rect 53319 65635 53431 65673
rect 53319 65627 53419 65635
rect 53477 65627 53589 65673
rect 53635 65635 53748 65673
rect 53682 65627 53748 65635
rect 53794 65635 53906 65673
rect 53794 65627 53841 65635
rect 53261 65583 53419 65627
rect 53471 65583 53630 65627
rect 53682 65583 53841 65627
rect 53893 65627 53906 65635
rect 53952 65635 54064 65673
rect 53952 65627 54052 65635
rect 54110 65627 54222 65673
rect 54268 65635 54540 65673
rect 53893 65583 54052 65627
rect 54104 65583 54263 65627
rect 54315 65583 54540 65635
rect 52428 65558 54540 65583
rect 52428 65512 54440 65558
rect 54486 65512 54540 65558
rect 52428 65509 54540 65512
rect 52428 65463 52483 65509
rect 52529 65463 52641 65509
rect 52687 65463 52799 65509
rect 52845 65463 52957 65509
rect 53003 65463 53115 65509
rect 53161 65463 53273 65509
rect 53319 65463 53431 65509
rect 53477 65463 53589 65509
rect 53635 65463 53748 65509
rect 53794 65463 53906 65509
rect 53952 65463 54064 65509
rect 54110 65463 54222 65509
rect 54268 65463 54540 65509
rect 52428 65418 54540 65463
rect 51043 65370 52015 65410
rect 42268 65325 42676 65370
rect 42116 65318 42155 65325
rect 42663 65324 42676 65325
rect 42722 65324 42779 65370
rect 42825 65324 42882 65370
rect 42928 65324 42986 65370
rect 43032 65324 43090 65370
rect 43136 65324 43194 65370
rect 43240 65324 43298 65370
rect 43344 65324 43402 65370
rect 43448 65324 43506 65370
rect 43552 65324 43610 65370
rect 43656 65324 43714 65370
rect 43760 65324 43818 65370
rect 43864 65324 43922 65370
rect 43968 65324 43981 65370
rect 44432 65324 44445 65370
rect 44491 65324 44559 65370
rect 44605 65324 44673 65370
rect 44719 65324 44787 65370
rect 44833 65324 44901 65370
rect 44947 65324 45346 65370
rect 45392 65324 45449 65370
rect 45495 65324 45552 65370
rect 45598 65324 45656 65370
rect 45702 65324 45760 65370
rect 45806 65324 45864 65370
rect 45910 65324 45968 65370
rect 46014 65324 46072 65370
rect 46118 65324 46176 65370
rect 46222 65324 46280 65370
rect 46326 65324 46384 65370
rect 46430 65324 46488 65370
rect 46534 65324 46592 65370
rect 46638 65324 47023 65370
rect 47101 65324 47114 65370
rect 48996 65324 49039 65370
rect 49099 65324 49156 65370
rect 49202 65324 49250 65370
rect 49305 65324 49362 65370
rect 49408 65324 49461 65370
rect 49513 65324 49568 65370
rect 49614 65324 49627 65370
rect 49744 65324 50014 65370
rect 50774 65324 50831 65370
rect 50877 65324 50934 65370
rect 50980 65324 51037 65370
rect 51133 65324 51140 65370
rect 51186 65324 51243 65370
rect 51289 65324 51292 65370
rect 40971 65277 42155 65318
rect 44432 65284 47023 65324
rect 48789 65318 48828 65324
rect 48880 65318 49039 65324
rect 49091 65318 49250 65324
rect 49302 65318 49461 65324
rect 49513 65318 49551 65324
rect 48789 65277 49551 65318
rect 51043 65318 51081 65324
rect 51133 65318 51292 65324
rect 51344 65324 51346 65370
rect 51392 65324 51449 65370
rect 51495 65324 51503 65370
rect 51598 65324 51655 65370
rect 51701 65324 51714 65370
rect 51804 65324 51861 65370
rect 51907 65324 51925 65370
rect 52010 65324 52023 65370
rect 52428 65366 52576 65418
rect 52628 65366 52787 65418
rect 52839 65366 52998 65418
rect 53050 65366 53209 65418
rect 53261 65366 53419 65418
rect 53471 65366 53630 65418
rect 53682 65366 53841 65418
rect 53893 65366 54052 65418
rect 54104 65366 54263 65418
rect 54315 65395 54540 65418
rect 54315 65366 54440 65395
rect 52428 65349 54440 65366
rect 54486 65349 54540 65395
rect 52428 65346 54540 65349
rect 51344 65318 51503 65324
rect 51555 65318 51714 65324
rect 51766 65318 51925 65324
rect 51977 65318 52015 65324
rect 51043 65278 52015 65318
rect 52428 65300 52483 65346
rect 52529 65300 52641 65346
rect 52687 65300 52799 65346
rect 52845 65300 52957 65346
rect 53003 65300 53115 65346
rect 53161 65300 53273 65346
rect 53319 65300 53431 65346
rect 53477 65300 53589 65346
rect 53635 65300 53748 65346
rect 53794 65300 53906 65346
rect 53952 65300 54064 65346
rect 54110 65300 54222 65346
rect 54268 65300 54540 65346
rect 52428 65243 54540 65300
rect 30583 65232 30955 65243
rect 30583 65186 30637 65232
rect 30683 65186 30955 65232
rect 30583 65068 30955 65186
rect 30583 65022 30637 65068
rect 30683 65022 30955 65068
rect 30583 64994 30955 65022
rect 54167 65232 54540 65243
rect 54167 65186 54440 65232
rect 54486 65186 54540 65232
rect 54167 65068 54540 65186
rect 54167 65022 54440 65068
rect 54486 65022 54540 65068
rect 27387 64820 28810 64866
rect 28856 64820 29196 64866
rect 29283 64953 30365 64994
rect 29283 64950 29582 64953
rect 29283 64904 29317 64950
rect 29363 64904 29478 64950
rect 29524 64904 29582 64950
rect 29283 64901 29582 64904
rect 29634 64950 29793 64953
rect 29845 64950 30005 64953
rect 29634 64904 29638 64950
rect 29684 64904 29793 64950
rect 29845 64904 29959 64950
rect 29634 64901 29793 64904
rect 29845 64901 30005 64904
rect 30057 64950 30216 64953
rect 30057 64904 30121 64950
rect 30167 64904 30216 64950
rect 30057 64901 30216 64904
rect 30268 64950 30365 64953
rect 30268 64904 30284 64950
rect 30330 64904 30365 64950
rect 30268 64901 30365 64904
rect 29283 64861 30365 64901
rect 30583 64953 32842 64994
rect 34247 64987 35008 64993
rect 30583 64901 30854 64953
rect 30906 64901 31065 64953
rect 31117 64901 31276 64953
rect 31328 64950 31486 64953
rect 31538 64950 31697 64953
rect 31749 64950 31909 64953
rect 31961 64950 32120 64953
rect 32172 64950 32330 64953
rect 32382 64950 32541 64953
rect 32593 64950 32752 64953
rect 32804 64950 32842 64953
rect 34246 64953 35008 64987
rect 34246 64950 34284 64953
rect 34336 64950 34495 64953
rect 34547 64950 34707 64953
rect 31328 64904 31349 64950
rect 33323 64904 33336 64950
rect 33671 64904 33684 64950
rect 33730 64904 33787 64950
rect 33833 64904 33890 64950
rect 33936 64904 33993 64950
rect 34039 64904 34096 64950
rect 34142 64904 34199 64950
rect 34245 64904 34284 64950
rect 34348 64904 34405 64950
rect 34451 64904 34495 64950
rect 34554 64904 34612 64950
rect 34658 64904 34707 64950
rect 31328 64901 31486 64904
rect 31538 64901 31697 64904
rect 31749 64901 31909 64904
rect 31961 64901 32120 64904
rect 32172 64901 32330 64904
rect 32382 64901 32541 64904
rect 32593 64901 32752 64904
rect 32804 64901 32842 64904
rect 30583 64866 32842 64901
rect 34246 64901 34284 64904
rect 34336 64901 34495 64904
rect 34547 64901 34707 64904
rect 34759 64901 34918 64953
rect 34970 64901 35008 64953
rect 34246 64867 35008 64901
rect 29544 64860 30306 64861
rect 27387 64744 29196 64820
rect 27387 64703 29116 64744
rect 27387 64657 28810 64703
rect 28856 64698 29116 64703
rect 29162 64698 29196 64744
rect 28856 64657 29196 64698
rect 27387 64581 29196 64657
rect 27387 64540 29116 64581
rect 27387 64494 28810 64540
rect 28856 64535 29116 64540
rect 29162 64535 29196 64581
rect 28856 64494 29196 64535
rect 27387 64417 29196 64494
rect 27387 64377 29116 64417
rect 27387 64331 28810 64377
rect 28856 64371 29116 64377
rect 29162 64371 29196 64417
rect 28856 64331 29196 64371
rect 27387 64254 29196 64331
rect 27387 64213 29116 64254
rect 27387 64167 28810 64213
rect 28856 64208 29116 64213
rect 29162 64208 29196 64254
rect 28856 64167 29196 64208
rect 27387 64053 29196 64167
rect 30583 64820 30637 64866
rect 30683 64860 32842 64866
rect 34247 64860 35008 64867
rect 35182 64987 36364 64994
rect 37946 64993 38324 64994
rect 35182 64953 36958 64987
rect 35182 64901 35220 64953
rect 35272 64901 35430 64953
rect 35482 64901 35641 64953
rect 35693 64901 35853 64953
rect 35905 64901 36064 64953
rect 36116 64901 36274 64953
rect 36326 64950 36958 64953
rect 36326 64904 36489 64950
rect 36723 64904 36958 64950
rect 36326 64901 36958 64904
rect 35182 64867 36958 64901
rect 37946 64953 38842 64993
rect 37946 64950 38330 64953
rect 38382 64950 38541 64953
rect 37946 64904 37957 64950
rect 38473 64904 38541 64950
rect 37946 64901 38330 64904
rect 38382 64901 38541 64904
rect 38593 64901 38752 64953
rect 38804 64901 38842 64953
rect 35182 64860 36364 64867
rect 37946 64860 38842 64901
rect 39014 64987 39322 64994
rect 40215 64987 40523 64994
rect 40788 64987 42986 65001
rect 54167 64994 54540 65022
rect 55927 65722 57736 65801
rect 55927 65676 56267 65722
rect 56313 65676 57736 65722
rect 58791 65914 59517 66894
rect 58791 65862 58858 65914
rect 58910 65862 58982 65914
rect 59034 65862 59106 65914
rect 59158 65862 59230 65914
rect 59282 65862 59354 65914
rect 59406 65862 59517 65914
rect 58791 65790 59517 65862
rect 58791 65738 58858 65790
rect 58910 65738 58982 65790
rect 59034 65738 59106 65790
rect 59158 65738 59230 65790
rect 59282 65738 59354 65790
rect 59406 65738 59517 65790
rect 58791 65678 59517 65738
rect 55927 65644 57736 65676
rect 55927 65598 55961 65644
rect 56007 65598 57736 65644
rect 55927 65558 57736 65598
rect 55927 65512 56267 65558
rect 56313 65512 57736 65558
rect 55927 65481 57736 65512
rect 55927 65435 55961 65481
rect 56007 65435 57736 65481
rect 55927 65395 57736 65435
rect 55927 65349 56267 65395
rect 56313 65349 57736 65395
rect 55927 65317 57736 65349
rect 55927 65271 55961 65317
rect 56007 65271 57736 65317
rect 55927 65232 57736 65271
rect 55927 65186 56267 65232
rect 56313 65186 57736 65232
rect 55927 65154 57736 65186
rect 55927 65108 55961 65154
rect 56007 65108 57736 65154
rect 55927 65068 57736 65108
rect 55927 65022 56267 65068
rect 56313 65022 57736 65068
rect 43753 64987 44514 64993
rect 39014 64953 39323 64987
rect 39014 64901 39052 64953
rect 39104 64950 39232 64953
rect 39108 64904 39220 64950
rect 39104 64901 39232 64904
rect 39284 64901 39323 64953
rect 30683 64826 31040 64860
rect 30683 64820 30855 64826
rect 30583 64780 30855 64820
rect 30901 64780 31040 64826
rect 30583 64703 31040 64780
rect 33484 64784 33552 64795
rect 33019 64729 33327 64770
rect 33019 64726 33057 64729
rect 33109 64726 33237 64729
rect 33289 64726 33327 64729
rect 30583 64657 30637 64703
rect 30683 64662 31040 64703
rect 31336 64680 31349 64726
rect 33323 64680 33336 64726
rect 30683 64657 30855 64662
rect 30583 64616 30855 64657
rect 30901 64616 31040 64662
rect 33019 64677 33057 64680
rect 33109 64677 33237 64680
rect 33289 64677 33327 64680
rect 33019 64637 33327 64677
rect 30583 64540 31040 64616
rect 30583 64494 30637 64540
rect 30683 64524 31040 64540
rect 30683 64502 31493 64524
rect 30683 64499 31349 64502
rect 30683 64494 30855 64499
rect 30583 64453 30855 64494
rect 30901 64456 31349 64499
rect 33323 64456 33336 64502
rect 30901 64453 31493 64456
rect 30583 64405 31493 64453
rect 30583 64377 31040 64405
rect 30583 64331 30637 64377
rect 30683 64336 31040 64377
rect 30683 64331 30855 64336
rect 30583 64290 30855 64331
rect 30901 64290 31040 64336
rect 33484 64362 33495 64784
rect 33541 64362 33552 64784
rect 33781 64737 34089 64778
rect 33781 64726 33819 64737
rect 33871 64726 33999 64737
rect 34051 64726 34089 64737
rect 33671 64680 33684 64726
rect 33730 64680 33787 64726
rect 33871 64685 33890 64726
rect 33833 64680 33890 64685
rect 33936 64680 33993 64726
rect 34051 64685 34096 64726
rect 34039 64680 34096 64685
rect 34142 64680 34199 64726
rect 34245 64680 34302 64726
rect 34348 64680 34405 64726
rect 34451 64680 34508 64726
rect 34554 64680 34612 64726
rect 34658 64680 34671 64726
rect 33781 64645 34089 64680
rect 35294 64651 36266 64691
rect 37853 64688 38161 64704
rect 35294 64639 35332 64651
rect 35384 64639 35543 64651
rect 35595 64639 35754 64651
rect 35806 64639 35965 64651
rect 36017 64639 36176 64651
rect 36228 64639 36266 64651
rect 36438 64639 36953 64688
rect 37439 64663 38161 64688
rect 37439 64639 37891 64663
rect 37943 64639 38071 64663
rect 38123 64639 38161 64663
rect 35260 64593 35273 64639
rect 35523 64599 35543 64639
rect 35523 64593 35580 64599
rect 35626 64593 35683 64639
rect 35729 64599 35754 64639
rect 35729 64593 35786 64599
rect 35832 64593 35889 64639
rect 35935 64599 35965 64639
rect 35935 64593 35992 64599
rect 36038 64593 36095 64639
rect 36141 64599 36176 64639
rect 36141 64593 36198 64599
rect 36244 64593 36301 64639
rect 36347 64593 36360 64639
rect 36438 64593 36854 64639
rect 36900 64593 36971 64639
rect 37017 64593 37088 64639
rect 37134 64593 37206 64639
rect 37252 64593 37324 64639
rect 37370 64593 37442 64639
rect 37488 64611 37891 64639
rect 37488 64593 37909 64611
rect 37955 64593 38026 64639
rect 38123 64611 38143 64639
rect 38072 64593 38143 64611
rect 38189 64593 38261 64639
rect 38307 64593 38379 64639
rect 38425 64593 38497 64639
rect 38543 64593 38556 64639
rect 35294 64559 36266 64593
rect 36438 64568 36953 64593
rect 37439 64571 38161 64593
rect 37439 64568 37931 64571
rect 34228 64502 34718 64531
rect 33671 64456 33684 64502
rect 33730 64456 33787 64502
rect 33833 64456 33890 64502
rect 33936 64456 33993 64502
rect 34039 64456 34096 64502
rect 34142 64456 34199 64502
rect 34245 64491 34302 64502
rect 34245 64456 34267 64491
rect 34348 64456 34405 64502
rect 34451 64491 34508 64502
rect 34499 64456 34508 64491
rect 34554 64456 34612 64502
rect 34658 64491 34718 64502
rect 34228 64439 34267 64456
rect 34319 64439 34447 64456
rect 34499 64439 34627 64456
rect 34679 64439 34718 64491
rect 36438 64465 36554 64568
rect 34228 64398 34718 64439
rect 34964 64415 36360 64459
rect 30583 64213 31040 64290
rect 33019 64281 33327 64322
rect 33019 64278 33057 64281
rect 33109 64278 33237 64281
rect 33289 64278 33327 64281
rect 33484 64280 33552 64362
rect 34964 64369 35273 64415
rect 35523 64369 35580 64415
rect 35626 64369 35683 64415
rect 35729 64369 35786 64415
rect 35832 64369 35889 64415
rect 35935 64369 35992 64415
rect 36038 64369 36095 64415
rect 36141 64369 36198 64415
rect 36244 64369 36301 64415
rect 36347 64369 36360 64415
rect 34964 64337 36360 64369
rect 34964 64280 35082 64337
rect 31336 64232 31349 64278
rect 33323 64232 33336 64278
rect 33484 64243 35082 64280
rect 30583 64167 30637 64213
rect 30683 64173 31040 64213
rect 33019 64229 33057 64232
rect 33109 64229 33237 64232
rect 33289 64229 33327 64232
rect 33019 64189 33327 64229
rect 33484 64197 33816 64243
rect 33862 64197 34002 64243
rect 34048 64197 34189 64243
rect 34235 64197 34376 64243
rect 34422 64197 34562 64243
rect 34608 64197 35082 64243
rect 36438 64325 36475 64465
rect 36521 64325 36554 64465
rect 33484 64189 35082 64197
rect 35294 64191 36266 64231
rect 36438 64225 36554 64325
rect 36640 64465 36773 64488
rect 36640 64416 36697 64465
rect 36640 64364 36678 64416
rect 36640 64325 36697 64364
rect 36743 64325 36773 64465
rect 38658 64467 38726 64478
rect 36924 64457 37685 64463
rect 36923 64456 37685 64457
rect 36923 64423 37931 64456
rect 36923 64415 36961 64423
rect 37013 64415 37172 64423
rect 37224 64415 37384 64423
rect 36841 64369 36854 64415
rect 36900 64371 36961 64415
rect 36900 64369 36971 64371
rect 37017 64369 37088 64415
rect 37134 64371 37172 64415
rect 37134 64369 37206 64371
rect 37252 64369 37324 64415
rect 37370 64371 37384 64415
rect 37436 64415 37595 64423
rect 37436 64371 37442 64415
rect 37370 64369 37442 64371
rect 37488 64371 37595 64415
rect 37647 64415 37931 64423
rect 37647 64371 37909 64415
rect 37488 64369 37909 64371
rect 37955 64369 38026 64415
rect 38072 64369 38143 64415
rect 38189 64369 38261 64415
rect 38307 64369 38379 64415
rect 38425 64369 38497 64415
rect 38543 64369 38556 64415
rect 36923 64337 37931 64369
rect 36924 64330 37685 64337
rect 36640 64305 36773 64325
rect 38658 64327 38669 64467
rect 38715 64327 38726 64467
rect 39014 64415 39323 64901
rect 39492 64964 42986 64987
rect 43704 64964 44514 64987
rect 39492 64953 44514 64964
rect 39492 64950 40253 64953
rect 39492 64904 39740 64950
rect 39786 64904 39862 64950
rect 39908 64904 39985 64950
rect 40031 64904 40108 64950
rect 40154 64904 40253 64950
rect 39492 64901 40253 64904
rect 40305 64901 40433 64953
rect 40485 64950 43790 64953
rect 40485 64904 40836 64950
rect 40882 64904 40994 64950
rect 41040 64904 41152 64950
rect 41198 64904 41310 64950
rect 41356 64904 41469 64950
rect 41515 64904 41627 64950
rect 41673 64904 41785 64950
rect 41831 64904 41943 64950
rect 41989 64904 42101 64950
rect 42147 64904 42259 64950
rect 42305 64904 42418 64950
rect 42464 64904 42576 64950
rect 42622 64904 42734 64950
rect 42780 64904 42892 64950
rect 42938 64904 43739 64950
rect 43785 64904 43790 64950
rect 40485 64901 43790 64904
rect 43842 64950 44001 64953
rect 43842 64904 43906 64950
rect 43952 64904 44001 64950
rect 43842 64901 44001 64904
rect 44053 64950 44213 64953
rect 44265 64950 44424 64953
rect 44053 64904 44071 64950
rect 44117 64904 44213 64950
rect 44282 64904 44424 64950
rect 44053 64901 44213 64904
rect 44265 64901 44424 64904
rect 44476 64901 44514 64953
rect 39492 64890 44514 64901
rect 39492 64867 42986 64890
rect 43704 64867 44514 64890
rect 39492 64415 39608 64867
rect 40215 64861 40523 64867
rect 40788 64853 42986 64867
rect 43753 64860 44514 64867
rect 44796 64987 45346 64993
rect 48800 64987 49982 64994
rect 50308 64987 50859 64994
rect 44796 64953 49982 64987
rect 44796 64950 44834 64953
rect 44886 64950 45045 64953
rect 45097 64950 45256 64953
rect 45308 64950 48838 64953
rect 44796 64904 44812 64950
rect 44886 64904 44925 64950
rect 44971 64904 45038 64950
rect 45097 64904 45151 64950
rect 45197 64904 45256 64950
rect 45310 64904 45619 64950
rect 45665 64904 45777 64950
rect 45823 64904 45935 64950
rect 45981 64904 46093 64950
rect 46139 64904 46251 64950
rect 46297 64904 46409 64950
rect 46455 64904 46568 64950
rect 46614 64904 46726 64950
rect 46772 64904 46884 64950
rect 46930 64904 47042 64950
rect 47088 64904 47200 64950
rect 47246 64904 47358 64950
rect 47404 64904 47516 64950
rect 47562 64904 47675 64950
rect 47721 64904 47833 64950
rect 47879 64904 47991 64950
rect 48037 64904 48149 64950
rect 48195 64904 48307 64950
rect 48353 64904 48465 64950
rect 48511 64904 48838 64950
rect 44796 64901 44834 64904
rect 44886 64901 45045 64904
rect 45097 64901 45256 64904
rect 45308 64901 48838 64904
rect 48890 64901 49048 64953
rect 49100 64901 49259 64953
rect 49311 64901 49471 64953
rect 49523 64901 49682 64953
rect 49734 64901 49892 64953
rect 49944 64901 49982 64953
rect 44796 64867 49982 64901
rect 50307 64953 50859 64987
rect 50307 64901 50346 64953
rect 50398 64950 50557 64953
rect 50609 64950 50768 64953
rect 50820 64950 50859 64953
rect 52278 64953 54540 64994
rect 52278 64950 52316 64953
rect 52368 64950 52527 64953
rect 52579 64950 52738 64953
rect 52790 64950 52948 64953
rect 53000 64950 53159 64953
rect 53211 64950 53371 64953
rect 53423 64950 53582 64953
rect 53634 64950 53792 64953
rect 50398 64904 50467 64950
rect 50513 64904 50557 64950
rect 50617 64904 50674 64950
rect 50720 64904 50768 64950
rect 50823 64904 50880 64950
rect 50926 64904 50983 64950
rect 51029 64904 51086 64950
rect 51132 64904 51189 64950
rect 51235 64904 51292 64950
rect 51338 64904 51395 64950
rect 51441 64904 51454 64950
rect 51789 64904 51802 64950
rect 53776 64904 53792 64950
rect 50398 64901 50557 64904
rect 50609 64901 50768 64904
rect 50820 64901 50859 64904
rect 50307 64867 50859 64901
rect 44796 64860 45346 64867
rect 43362 64809 43524 64820
rect 39737 64726 39866 64755
rect 40246 64737 40362 64774
rect 43362 64763 43373 64809
rect 43513 64763 43524 64809
rect 43362 64756 43524 64763
rect 39727 64680 39740 64726
rect 39786 64715 39862 64726
rect 39827 64680 39862 64715
rect 39908 64680 39985 64726
rect 40031 64680 40108 64726
rect 40154 64680 40167 64726
rect 40246 64691 40281 64737
rect 40327 64691 40362 64737
rect 39737 64663 39775 64680
rect 39827 64663 39866 64680
rect 39737 64636 39866 64663
rect 39737 64623 39865 64636
rect 39923 64500 40085 64540
rect 39923 64448 39994 64500
rect 40046 64448 40085 64500
rect 39008 64369 39021 64415
rect 39067 64369 39144 64415
rect 39190 64369 39267 64415
rect 39313 64369 39326 64415
rect 39492 64369 39641 64415
rect 39687 64369 39730 64415
rect 39014 64337 39323 64369
rect 39492 64337 39608 64369
rect 37853 64225 38161 64230
rect 36438 64191 36953 64225
rect 37439 64191 38161 64225
rect 38658 64205 38726 64327
rect 39923 64317 40085 64448
rect 39809 64314 40085 64317
rect 39809 64306 39994 64314
rect 39809 64260 39844 64306
rect 39890 64262 39994 64306
rect 40046 64293 40085 64314
rect 40246 64293 40362 64691
rect 40718 64715 43524 64756
rect 45584 64786 48546 64867
rect 48800 64860 49982 64867
rect 50308 64860 50859 64867
rect 52278 64901 52316 64904
rect 52368 64901 52527 64904
rect 52579 64901 52738 64904
rect 52790 64901 52948 64904
rect 53000 64901 53159 64904
rect 53211 64901 53371 64904
rect 53423 64901 53582 64904
rect 53634 64901 53792 64904
rect 53844 64901 54003 64953
rect 54055 64901 54214 64953
rect 54266 64901 54540 64953
rect 52278 64866 54540 64901
rect 52278 64860 54440 64866
rect 45584 64740 45619 64786
rect 45665 64740 45777 64786
rect 45823 64740 45935 64786
rect 45981 64740 46093 64786
rect 46139 64740 46251 64786
rect 46297 64740 46409 64786
rect 46455 64740 46568 64786
rect 46614 64740 46726 64786
rect 46772 64740 46884 64786
rect 46930 64740 47042 64786
rect 47088 64740 47200 64786
rect 47246 64740 47358 64786
rect 47404 64740 47516 64786
rect 47562 64740 47675 64786
rect 47721 64740 47833 64786
rect 47879 64740 47991 64786
rect 48037 64740 48149 64786
rect 48195 64740 48307 64786
rect 48353 64740 48465 64786
rect 48511 64740 48546 64786
rect 54085 64826 54440 64860
rect 54085 64780 54223 64826
rect 54269 64820 54440 64826
rect 54486 64820 54540 64866
rect 54758 64953 55840 64994
rect 54758 64950 54855 64953
rect 54758 64904 54793 64950
rect 54839 64904 54855 64950
rect 54758 64901 54855 64904
rect 54907 64950 55066 64953
rect 54907 64904 54956 64950
rect 55002 64904 55066 64950
rect 54907 64901 55066 64904
rect 55118 64950 55278 64953
rect 55330 64950 55489 64953
rect 55164 64904 55278 64950
rect 55330 64904 55439 64950
rect 55485 64904 55489 64950
rect 55118 64901 55278 64904
rect 55330 64901 55489 64904
rect 55541 64950 55840 64953
rect 55541 64904 55599 64950
rect 55645 64904 55760 64950
rect 55806 64904 55840 64950
rect 55541 64901 55840 64904
rect 54758 64861 55840 64901
rect 55927 64866 57736 65022
rect 54817 64860 55579 64861
rect 54269 64780 54540 64820
rect 40718 64663 41935 64715
rect 41987 64663 43524 64715
rect 40718 64622 43524 64663
rect 44605 64680 44812 64726
rect 44858 64680 44925 64726
rect 44971 64680 45038 64726
rect 45084 64680 45151 64726
rect 45197 64680 45264 64726
rect 45310 64680 45323 64726
rect 45584 64704 48546 64740
rect 51035 64729 51343 64770
rect 51035 64726 51073 64729
rect 51125 64726 51253 64729
rect 51305 64726 51343 64729
rect 51589 64754 51657 64765
rect 44341 64614 44509 64625
rect 44341 64568 44358 64614
rect 44498 64568 44509 64614
rect 44341 64524 44509 64568
rect 42229 64484 44509 64524
rect 42229 64432 42312 64484
rect 42364 64432 44509 64484
rect 42229 64391 44509 64432
rect 44605 64293 44721 64680
rect 48905 64654 49877 64694
rect 50454 64680 50467 64726
rect 50513 64680 50571 64726
rect 50617 64680 50674 64726
rect 50720 64680 50777 64726
rect 50823 64680 50880 64726
rect 50926 64680 50983 64726
rect 51029 64680 51073 64726
rect 51132 64680 51189 64726
rect 51235 64680 51253 64726
rect 51338 64680 51395 64726
rect 51441 64680 51454 64726
rect 48905 64639 48943 64654
rect 48995 64639 49154 64654
rect 49206 64639 49365 64654
rect 49417 64639 49576 64654
rect 49628 64639 49787 64654
rect 49839 64639 49877 64654
rect 48765 64593 48778 64639
rect 48824 64593 48881 64639
rect 48927 64602 48943 64639
rect 48927 64593 48984 64602
rect 49030 64593 49087 64639
rect 49133 64602 49154 64639
rect 49133 64593 49190 64602
rect 49236 64593 49293 64639
rect 49339 64602 49365 64639
rect 49339 64593 49396 64602
rect 49442 64593 49499 64639
rect 49545 64602 49576 64639
rect 49545 64593 49602 64602
rect 49852 64593 49877 64639
rect 51035 64677 51073 64680
rect 51125 64677 51253 64680
rect 51305 64677 51343 64680
rect 51035 64637 51343 64677
rect 48557 64547 48687 64588
rect 48905 64562 49877 64593
rect 44901 64502 45241 64531
rect 44799 64456 44812 64502
rect 44858 64456 44925 64502
rect 44971 64491 45038 64502
rect 44991 64456 45038 64491
rect 45084 64456 45151 64502
rect 45197 64491 45264 64502
rect 45203 64456 45264 64491
rect 45310 64456 45323 64502
rect 48557 64495 48596 64547
rect 48648 64495 48687 64547
rect 48557 64492 48687 64495
rect 44901 64439 44939 64456
rect 44991 64439 45151 64456
rect 45203 64439 45241 64456
rect 44901 64398 45241 64439
rect 45400 64383 48379 64416
rect 45400 64337 45464 64383
rect 45604 64375 48379 64383
rect 45400 64323 45597 64337
rect 45649 64323 48379 64375
rect 40046 64278 44918 64293
rect 45400 64282 48379 64323
rect 48557 64352 48622 64492
rect 48668 64352 48687 64492
rect 50262 64502 50812 64531
rect 50262 64491 50467 64502
rect 50513 64491 50571 64502
rect 49820 64415 50160 64456
rect 48765 64369 48778 64415
rect 48824 64369 48881 64415
rect 48927 64369 48984 64415
rect 49030 64369 49087 64415
rect 49133 64369 49190 64415
rect 49236 64369 49293 64415
rect 49339 64369 49396 64415
rect 49442 64369 49499 64415
rect 49545 64369 49602 64415
rect 49852 64369 50160 64415
rect 50262 64439 50300 64491
rect 50352 64456 50467 64491
rect 50563 64456 50571 64491
rect 50617 64456 50674 64502
rect 50720 64491 50777 64502
rect 50720 64456 50722 64491
rect 50352 64439 50511 64456
rect 50563 64439 50722 64456
rect 50774 64456 50777 64491
rect 50823 64456 50880 64502
rect 50926 64456 50983 64502
rect 51029 64456 51086 64502
rect 51132 64456 51189 64502
rect 51235 64456 51292 64502
rect 51338 64456 51395 64502
rect 51441 64456 51454 64502
rect 50774 64439 50812 64456
rect 50262 64398 50812 64439
rect 48557 64329 48687 64352
rect 49820 64337 50160 64369
rect 40046 64262 44812 64278
rect 39890 64260 44812 64262
rect 39809 64257 44812 64260
rect 39809 64211 43739 64257
rect 43785 64211 43906 64257
rect 43952 64211 44071 64257
rect 44117 64211 44236 64257
rect 44282 64232 44812 64257
rect 44858 64232 44925 64278
rect 44971 64232 45038 64278
rect 45084 64232 45151 64278
rect 45197 64232 45264 64278
rect 45310 64232 45323 64278
rect 48557 64277 48596 64329
rect 48648 64277 48687 64329
rect 48557 64237 48687 64277
rect 50044 64280 50160 64337
rect 51589 64332 51600 64754
rect 51646 64332 51657 64754
rect 51797 64726 52105 64763
rect 51789 64680 51802 64726
rect 53776 64680 53789 64726
rect 54085 64703 54540 64780
rect 51797 64670 51835 64680
rect 51887 64670 52015 64680
rect 52067 64670 52105 64680
rect 51797 64630 52105 64670
rect 54085 64662 54440 64703
rect 54085 64616 54223 64662
rect 54269 64657 54440 64662
rect 54486 64657 54540 64703
rect 54269 64616 54540 64657
rect 54085 64540 54540 64616
rect 54085 64524 54440 64540
rect 53585 64502 54440 64524
rect 51789 64456 51802 64502
rect 53776 64494 54440 64502
rect 54486 64494 54540 64540
rect 53776 64456 54540 64494
rect 53585 64405 54540 64456
rect 51589 64280 51657 64332
rect 54085 64377 54540 64405
rect 54085 64331 54440 64377
rect 54486 64331 54540 64377
rect 50044 64243 51657 64280
rect 51797 64278 52105 64300
rect 44282 64211 44918 64232
rect 38658 64191 39723 64205
rect 30683 64167 30855 64173
rect 30583 64127 30855 64167
rect 30901 64127 31040 64173
rect 33484 64160 34643 64189
rect 35260 64145 35273 64191
rect 35523 64145 35543 64191
rect 35626 64145 35683 64191
rect 35729 64145 35754 64191
rect 35832 64145 35889 64191
rect 35935 64145 35965 64191
rect 36038 64145 36095 64191
rect 36141 64145 36176 64191
rect 36244 64145 36301 64191
rect 36347 64145 36360 64191
rect 36438 64145 36854 64191
rect 36900 64145 36971 64191
rect 37017 64145 37088 64191
rect 37134 64145 37206 64191
rect 37252 64145 37324 64191
rect 37370 64145 37442 64191
rect 37488 64189 37909 64191
rect 37488 64145 37891 64189
rect 37955 64145 38026 64191
rect 38072 64189 38143 64191
rect 38123 64145 38143 64189
rect 38189 64145 38261 64191
rect 38307 64145 38379 64191
rect 38425 64145 38497 64191
rect 38543 64145 38556 64191
rect 38658 64145 39021 64191
rect 39067 64145 39144 64191
rect 39190 64145 39267 64191
rect 39313 64145 39641 64191
rect 39687 64145 39730 64191
rect 39809 64173 44918 64211
rect 48905 64191 49877 64231
rect 48765 64145 48778 64191
rect 48824 64145 48881 64191
rect 48927 64145 48943 64191
rect 49030 64145 49087 64191
rect 49133 64145 49154 64191
rect 49236 64145 49293 64191
rect 49339 64145 49365 64191
rect 49442 64145 49499 64191
rect 49545 64145 49576 64191
rect 49852 64145 49877 64191
rect 50044 64197 50516 64243
rect 50562 64197 50703 64243
rect 50749 64197 50890 64243
rect 50936 64197 51076 64243
rect 51122 64197 51263 64243
rect 51309 64197 51657 64243
rect 51789 64232 51802 64278
rect 53776 64232 53789 64278
rect 50044 64187 51657 64197
rect 50481 64160 51657 64187
rect 51797 64207 51835 64232
rect 51887 64207 52015 64232
rect 52067 64207 52105 64232
rect 51797 64167 52105 64207
rect 54085 64213 54540 64331
rect 54085 64173 54440 64213
rect 30583 64094 31040 64127
rect 35294 64139 35332 64145
rect 35384 64139 35543 64145
rect 35595 64139 35754 64145
rect 35806 64139 35965 64145
rect 36017 64139 36176 64145
rect 36228 64139 36266 64145
rect 34870 64094 35025 64101
rect 35294 64099 36266 64139
rect 36438 64105 36953 64145
rect 37439 64137 37891 64145
rect 37943 64137 38071 64145
rect 38123 64137 38161 64145
rect 37439 64105 38161 64137
rect 37853 64097 38161 64105
rect 27387 64001 27790 64053
rect 27842 64001 28001 64053
rect 28053 64001 28212 64053
rect 28264 64001 28423 64053
rect 28475 64001 28634 64053
rect 28686 64050 28845 64053
rect 28686 64004 28810 64050
rect 28686 64001 28845 64004
rect 28897 64001 29056 64053
rect 29108 64001 29196 64053
rect 27387 63887 29196 64001
rect 29283 64053 30365 64094
rect 29283 64050 29582 64053
rect 29283 64004 29317 64050
rect 29363 64004 29478 64050
rect 29524 64004 29582 64050
rect 29283 64001 29582 64004
rect 29634 64050 29793 64053
rect 29845 64050 30005 64053
rect 29634 64004 29638 64050
rect 29684 64004 29793 64050
rect 29845 64004 29959 64050
rect 29634 64001 29793 64004
rect 29845 64001 30005 64004
rect 30057 64050 30216 64053
rect 30057 64004 30121 64050
rect 30167 64004 30216 64050
rect 30057 64001 30216 64004
rect 30268 64050 30365 64053
rect 30268 64004 30284 64050
rect 30330 64004 30365 64050
rect 30268 64001 30365 64004
rect 29283 63961 30365 64001
rect 30583 64053 32842 64094
rect 30583 64050 30854 64053
rect 30583 64004 30637 64050
rect 30683 64004 30854 64050
rect 30583 64001 30854 64004
rect 30906 64001 31065 64053
rect 31117 64001 31276 64053
rect 31328 64001 31486 64053
rect 31538 64001 31697 64053
rect 31749 64001 31909 64053
rect 31961 64001 32120 64053
rect 32172 64001 32330 64053
rect 32382 64001 32541 64053
rect 32593 64001 32752 64053
rect 32804 64001 32842 64053
rect 29544 63960 30306 63961
rect 30583 63960 32842 64001
rect 34717 64053 35025 64094
rect 38658 64085 39723 64145
rect 48905 64139 48943 64145
rect 48995 64139 49154 64145
rect 49206 64139 49365 64145
rect 49417 64139 49576 64145
rect 49628 64139 49787 64145
rect 49839 64139 49877 64145
rect 48905 64099 49877 64139
rect 54085 64127 54223 64173
rect 54269 64167 54440 64173
rect 54486 64167 54540 64213
rect 54269 64127 54540 64167
rect 50099 64094 50255 64101
rect 54085 64094 54540 64127
rect 55927 64820 56267 64866
rect 56313 64820 57736 64866
rect 55927 64744 57736 64820
rect 55927 64698 55961 64744
rect 56007 64703 57736 64744
rect 56007 64698 56267 64703
rect 55927 64657 56267 64698
rect 56313 64657 57736 64703
rect 55927 64581 57736 64657
rect 55927 64535 55961 64581
rect 56007 64540 57736 64581
rect 56007 64535 56267 64540
rect 55927 64494 56267 64535
rect 56313 64494 57736 64540
rect 55927 64417 57736 64494
rect 55927 64371 55961 64417
rect 56007 64377 57736 64417
rect 56007 64371 56267 64377
rect 55927 64331 56267 64371
rect 56313 64331 57736 64377
rect 55927 64254 57736 64331
rect 55927 64208 55961 64254
rect 56007 64213 57736 64254
rect 56007 64208 56267 64213
rect 55927 64167 56267 64208
rect 56313 64167 57736 64213
rect 34717 64001 34755 64053
rect 34807 64050 34935 64053
rect 34807 64004 34916 64050
rect 34807 64001 34935 64004
rect 34987 64001 35025 64053
rect 34717 63960 35025 64001
rect 50099 64053 50408 64094
rect 50099 64001 50138 64053
rect 50190 64050 50318 64053
rect 50206 64004 50318 64050
rect 50190 64001 50318 64004
rect 50370 64001 50408 64053
rect 27387 63841 28810 63887
rect 28856 63844 29196 63887
rect 28856 63841 29116 63844
rect 27387 63798 29116 63841
rect 29162 63798 29196 63844
rect 27387 63723 29196 63798
rect 27387 63677 28810 63723
rect 28856 63681 29196 63723
rect 28856 63677 29116 63681
rect 27387 63635 29116 63677
rect 29162 63635 29196 63681
rect 27387 63560 29196 63635
rect 27387 63514 28810 63560
rect 28856 63517 29196 63560
rect 28856 63514 29116 63517
rect 27387 63471 29116 63514
rect 29162 63471 29196 63517
rect 27387 63397 29196 63471
rect 27387 63351 28810 63397
rect 28856 63354 29196 63397
rect 28856 63351 29116 63354
rect 27387 63308 29116 63351
rect 29162 63308 29196 63354
rect 27387 63234 29196 63308
rect 27387 63188 28810 63234
rect 28856 63188 29196 63234
rect 30583 63927 31040 63960
rect 34870 63953 35025 63960
rect 30583 63887 30855 63927
rect 30583 63841 30637 63887
rect 30683 63881 30855 63887
rect 30901 63881 31040 63927
rect 35294 63915 36266 63955
rect 37853 63949 38161 63957
rect 35294 63909 35332 63915
rect 35384 63909 35543 63915
rect 35595 63909 35754 63915
rect 35806 63909 35965 63915
rect 36017 63909 36176 63915
rect 36228 63909 36266 63915
rect 36438 63909 36953 63949
rect 37439 63917 38161 63949
rect 37439 63909 37891 63917
rect 37943 63909 38071 63917
rect 38123 63909 38161 63917
rect 38658 63909 39723 63969
rect 50099 63960 50408 64001
rect 52278 64053 54540 64094
rect 52278 64001 52316 64053
rect 52368 64001 52527 64053
rect 52579 64001 52738 64053
rect 52790 64001 52948 64053
rect 53000 64001 53159 64053
rect 53211 64001 53371 64053
rect 53423 64001 53582 64053
rect 53634 64001 53792 64053
rect 53844 64001 54003 64053
rect 54055 64001 54214 64053
rect 54266 64050 54540 64053
rect 54266 64004 54440 64050
rect 54486 64004 54540 64050
rect 54266 64001 54540 64004
rect 52278 63960 54540 64001
rect 54758 64053 55840 64094
rect 54758 64050 54855 64053
rect 54758 64004 54793 64050
rect 54839 64004 54855 64050
rect 54758 64001 54855 64004
rect 54907 64050 55066 64053
rect 54907 64004 54956 64050
rect 55002 64004 55066 64050
rect 54907 64001 55066 64004
rect 55118 64050 55278 64053
rect 55330 64050 55489 64053
rect 55164 64004 55278 64050
rect 55330 64004 55439 64050
rect 55485 64004 55489 64050
rect 55118 64001 55278 64004
rect 55330 64001 55489 64004
rect 55541 64050 55840 64053
rect 55541 64004 55599 64050
rect 55645 64004 55760 64050
rect 55806 64004 55840 64050
rect 55541 64001 55840 64004
rect 54758 63961 55840 64001
rect 55927 64053 57736 64167
rect 55927 64001 56015 64053
rect 56067 64001 56226 64053
rect 56278 64050 56437 64053
rect 56313 64004 56437 64050
rect 56278 64001 56437 64004
rect 56489 64001 56648 64053
rect 56700 64001 56859 64053
rect 56911 64001 57070 64053
rect 57122 64001 57281 64053
rect 57333 64001 57736 64053
rect 54817 63960 55579 63961
rect 48905 63915 49877 63955
rect 50099 63953 50255 63960
rect 48905 63909 48943 63915
rect 48995 63909 49154 63915
rect 49206 63909 49365 63915
rect 49417 63909 49576 63915
rect 49628 63909 49787 63915
rect 49839 63909 49877 63915
rect 30683 63841 31040 63881
rect 33484 63865 34643 63894
rect 30583 63764 31040 63841
rect 33019 63825 33327 63865
rect 33019 63822 33057 63825
rect 33109 63822 33237 63825
rect 33289 63822 33327 63825
rect 33484 63857 35082 63865
rect 35260 63863 35273 63909
rect 35523 63863 35543 63909
rect 35626 63863 35683 63909
rect 35729 63863 35754 63909
rect 35832 63863 35889 63909
rect 35935 63863 35965 63909
rect 36038 63863 36095 63909
rect 36141 63863 36176 63909
rect 36244 63863 36301 63909
rect 36347 63863 36360 63909
rect 36438 63863 36854 63909
rect 36900 63863 36971 63909
rect 37017 63863 37088 63909
rect 37134 63863 37206 63909
rect 37252 63863 37324 63909
rect 37370 63863 37442 63909
rect 37488 63865 37891 63909
rect 37488 63863 37909 63865
rect 37955 63863 38026 63909
rect 38123 63865 38143 63909
rect 38072 63863 38143 63865
rect 38189 63863 38261 63909
rect 38307 63863 38379 63909
rect 38425 63863 38497 63909
rect 38543 63863 38556 63909
rect 38658 63863 39021 63909
rect 39067 63863 39144 63909
rect 39190 63863 39267 63909
rect 39313 63863 39641 63909
rect 39687 63863 39730 63909
rect 31336 63776 31349 63822
rect 33323 63776 33336 63822
rect 33484 63811 33816 63857
rect 33862 63811 34002 63857
rect 34048 63811 34189 63857
rect 34235 63811 34376 63857
rect 34422 63811 34562 63857
rect 34608 63811 35082 63857
rect 35294 63823 36266 63863
rect 36438 63829 36953 63863
rect 37439 63829 38161 63863
rect 30583 63723 30855 63764
rect 30583 63677 30637 63723
rect 30683 63718 30855 63723
rect 30901 63718 31040 63764
rect 33019 63773 33057 63776
rect 33109 63773 33237 63776
rect 33289 63773 33327 63776
rect 33019 63732 33327 63773
rect 33484 63774 35082 63811
rect 30683 63677 31040 63718
rect 30583 63649 31040 63677
rect 33484 63692 33552 63774
rect 30583 63601 31493 63649
rect 30583 63560 30855 63601
rect 30583 63514 30637 63560
rect 30683 63555 30855 63560
rect 30901 63598 31493 63601
rect 30901 63555 31349 63598
rect 30683 63552 31349 63555
rect 33323 63552 33336 63598
rect 30683 63530 31493 63552
rect 30683 63514 31040 63530
rect 30583 63438 31040 63514
rect 30583 63397 30855 63438
rect 30583 63351 30637 63397
rect 30683 63392 30855 63397
rect 30901 63392 31040 63438
rect 30683 63351 31040 63392
rect 33019 63377 33327 63417
rect 33019 63374 33057 63377
rect 33109 63374 33237 63377
rect 33289 63374 33327 63377
rect 30583 63274 31040 63351
rect 31336 63328 31349 63374
rect 33323 63328 33336 63374
rect 33019 63325 33057 63328
rect 33109 63325 33237 63328
rect 33289 63325 33327 63328
rect 33019 63284 33327 63325
rect 30583 63234 30855 63274
rect 27387 63066 29196 63188
rect 27387 63020 28810 63066
rect 28856 63020 29196 63066
rect 29283 63153 30365 63194
rect 29283 63150 29582 63153
rect 29283 63104 29317 63150
rect 29363 63104 29478 63150
rect 29524 63104 29582 63150
rect 29283 63101 29582 63104
rect 29634 63150 29793 63153
rect 29845 63150 30005 63153
rect 29634 63104 29638 63150
rect 29684 63104 29793 63150
rect 29845 63104 29959 63150
rect 29634 63101 29793 63104
rect 29845 63101 30005 63104
rect 30057 63150 30216 63153
rect 30057 63104 30121 63150
rect 30167 63104 30216 63150
rect 30057 63101 30216 63104
rect 30268 63150 30365 63153
rect 30268 63104 30284 63150
rect 30330 63104 30365 63150
rect 30268 63101 30365 63104
rect 29283 63061 30365 63101
rect 30583 63188 30637 63234
rect 30683 63228 30855 63234
rect 30901 63228 31040 63274
rect 33484 63270 33495 63692
rect 33541 63270 33552 63692
rect 34964 63717 35082 63774
rect 36438 63729 36554 63829
rect 37853 63824 38161 63829
rect 38658 63849 39723 63863
rect 34964 63685 36360 63717
rect 34228 63615 34718 63656
rect 34228 63598 34267 63615
rect 34319 63598 34447 63615
rect 34499 63598 34627 63615
rect 33671 63552 33684 63598
rect 33730 63552 33787 63598
rect 33833 63552 33890 63598
rect 33936 63552 33993 63598
rect 34039 63552 34096 63598
rect 34142 63552 34199 63598
rect 34245 63563 34267 63598
rect 34245 63552 34302 63563
rect 34348 63552 34405 63598
rect 34499 63563 34508 63598
rect 34451 63552 34508 63563
rect 34554 63552 34612 63598
rect 34679 63563 34718 63615
rect 34964 63639 35273 63685
rect 35523 63639 35580 63685
rect 35626 63639 35683 63685
rect 35729 63639 35786 63685
rect 35832 63639 35889 63685
rect 35935 63639 35992 63685
rect 36038 63639 36095 63685
rect 36141 63639 36198 63685
rect 36244 63639 36301 63685
rect 36347 63639 36360 63685
rect 34964 63595 36360 63639
rect 34658 63552 34718 63563
rect 34228 63523 34718 63552
rect 36438 63589 36475 63729
rect 36521 63589 36554 63729
rect 35294 63461 36266 63495
rect 36438 63486 36554 63589
rect 36640 63729 36773 63749
rect 36640 63690 36697 63729
rect 36640 63638 36678 63690
rect 36640 63589 36697 63638
rect 36743 63589 36773 63729
rect 38658 63727 38726 63849
rect 39809 63843 44918 63881
rect 48765 63863 48778 63909
rect 48824 63863 48881 63909
rect 48927 63863 48943 63909
rect 49030 63863 49087 63909
rect 49133 63863 49154 63909
rect 49236 63863 49293 63909
rect 49339 63863 49365 63909
rect 49442 63863 49499 63909
rect 49545 63863 49576 63909
rect 49852 63863 49877 63909
rect 54085 63927 54540 63960
rect 50481 63867 51657 63894
rect 39809 63797 43739 63843
rect 43785 63797 43906 63843
rect 43952 63797 44071 63843
rect 44117 63797 44236 63843
rect 44282 63822 44918 63843
rect 48905 63823 49877 63863
rect 50044 63857 51657 63867
rect 44282 63797 44812 63822
rect 39809 63794 44812 63797
rect 39809 63748 39844 63794
rect 39890 63792 44812 63794
rect 39890 63748 39994 63792
rect 39809 63740 39994 63748
rect 40046 63776 44812 63792
rect 44858 63776 44925 63822
rect 44971 63776 45038 63822
rect 45084 63776 45151 63822
rect 45197 63776 45264 63822
rect 45310 63776 45323 63822
rect 48557 63777 48687 63817
rect 40046 63761 44918 63776
rect 40046 63740 40085 63761
rect 39809 63737 40085 63740
rect 36924 63717 37685 63724
rect 36923 63685 37931 63717
rect 36841 63639 36854 63685
rect 36900 63683 36971 63685
rect 36900 63639 36961 63683
rect 37017 63639 37088 63685
rect 37134 63683 37206 63685
rect 37134 63639 37172 63683
rect 37252 63639 37324 63685
rect 37370 63683 37442 63685
rect 37370 63639 37384 63683
rect 36923 63631 36961 63639
rect 37013 63631 37172 63639
rect 37224 63631 37384 63639
rect 37436 63639 37442 63683
rect 37488 63683 37909 63685
rect 37488 63639 37595 63683
rect 37436 63631 37595 63639
rect 37647 63639 37909 63683
rect 37955 63639 38026 63685
rect 38072 63639 38143 63685
rect 38189 63639 38261 63685
rect 38307 63639 38379 63685
rect 38425 63639 38497 63685
rect 38543 63639 38556 63685
rect 37647 63631 37931 63639
rect 36923 63598 37931 63631
rect 36923 63597 37685 63598
rect 36924 63591 37685 63597
rect 36640 63566 36773 63589
rect 38658 63587 38669 63727
rect 38715 63587 38726 63727
rect 39014 63685 39323 63717
rect 39492 63685 39608 63717
rect 39008 63639 39021 63685
rect 39067 63639 39144 63685
rect 39190 63639 39267 63685
rect 39313 63639 39326 63685
rect 39492 63639 39641 63685
rect 39687 63639 39730 63685
rect 38658 63576 38726 63587
rect 36438 63461 36953 63486
rect 37439 63483 37931 63486
rect 37439 63461 38161 63483
rect 35260 63415 35273 63461
rect 35523 63455 35580 63461
rect 35523 63415 35543 63455
rect 35626 63415 35683 63461
rect 35729 63455 35786 63461
rect 35729 63415 35754 63455
rect 35832 63415 35889 63461
rect 35935 63455 35992 63461
rect 35935 63415 35965 63455
rect 36038 63415 36095 63461
rect 36141 63455 36198 63461
rect 36141 63415 36176 63455
rect 36244 63415 36301 63461
rect 36347 63415 36360 63461
rect 36438 63415 36854 63461
rect 36900 63415 36971 63461
rect 37017 63415 37088 63461
rect 37134 63415 37206 63461
rect 37252 63415 37324 63461
rect 37370 63415 37442 63461
rect 37488 63443 37909 63461
rect 37488 63415 37891 63443
rect 37955 63415 38026 63461
rect 38072 63443 38143 63461
rect 38123 63415 38143 63443
rect 38189 63415 38261 63461
rect 38307 63415 38379 63461
rect 38425 63415 38497 63461
rect 38543 63415 38556 63461
rect 33781 63374 34089 63409
rect 35294 63403 35332 63415
rect 35384 63403 35543 63415
rect 35595 63403 35754 63415
rect 35806 63403 35965 63415
rect 36017 63403 36176 63415
rect 36228 63403 36266 63415
rect 33671 63328 33684 63374
rect 33730 63328 33787 63374
rect 33833 63369 33890 63374
rect 33871 63328 33890 63369
rect 33936 63328 33993 63374
rect 34039 63369 34096 63374
rect 34051 63328 34096 63369
rect 34142 63328 34199 63374
rect 34245 63328 34302 63374
rect 34348 63328 34405 63374
rect 34451 63328 34508 63374
rect 34554 63328 34612 63374
rect 34658 63328 34671 63374
rect 35294 63363 36266 63403
rect 36438 63366 36953 63415
rect 37439 63391 37891 63415
rect 37943 63391 38071 63415
rect 38123 63391 38161 63415
rect 37439 63366 38161 63391
rect 37853 63350 38161 63366
rect 33781 63317 33819 63328
rect 33871 63317 33999 63328
rect 34051 63317 34089 63328
rect 33781 63276 34089 63317
rect 33484 63259 33552 63270
rect 30683 63194 31040 63228
rect 30683 63188 32842 63194
rect 30583 63153 32842 63188
rect 34247 63187 35008 63194
rect 30583 63101 30854 63153
rect 30906 63101 31065 63153
rect 31117 63101 31276 63153
rect 31328 63150 31486 63153
rect 31538 63150 31697 63153
rect 31749 63150 31909 63153
rect 31961 63150 32120 63153
rect 32172 63150 32330 63153
rect 32382 63150 32541 63153
rect 32593 63150 32752 63153
rect 32804 63150 32842 63153
rect 34246 63153 35008 63187
rect 34246 63150 34284 63153
rect 34336 63150 34495 63153
rect 34547 63150 34707 63153
rect 31328 63104 31349 63150
rect 33323 63104 33336 63150
rect 33671 63104 33684 63150
rect 33730 63104 33787 63150
rect 33833 63104 33890 63150
rect 33936 63104 33993 63150
rect 34039 63104 34096 63150
rect 34142 63104 34199 63150
rect 34245 63104 34284 63150
rect 34348 63104 34405 63150
rect 34451 63104 34495 63150
rect 34554 63104 34612 63150
rect 34658 63104 34707 63150
rect 31328 63101 31486 63104
rect 31538 63101 31697 63104
rect 31749 63101 31909 63104
rect 31961 63101 32120 63104
rect 32172 63101 32330 63104
rect 32382 63101 32541 63104
rect 32593 63101 32752 63104
rect 32804 63101 32842 63104
rect 30583 63066 32842 63101
rect 34246 63101 34284 63104
rect 34336 63101 34495 63104
rect 34547 63101 34707 63104
rect 34759 63101 34918 63153
rect 34970 63101 35008 63153
rect 34246 63067 35008 63101
rect 29544 63060 30306 63061
rect 27387 62944 29196 63020
rect 27387 62903 29116 62944
rect 27387 62857 28810 62903
rect 28856 62898 29116 62903
rect 29162 62898 29196 62944
rect 28856 62857 29196 62898
rect 27387 62781 29196 62857
rect 27387 62740 29116 62781
rect 27387 62694 28810 62740
rect 28856 62735 29116 62740
rect 29162 62735 29196 62781
rect 28856 62694 29196 62735
rect 27387 62617 29196 62694
rect 27387 62577 29116 62617
rect 27387 62531 28810 62577
rect 28856 62571 29116 62577
rect 29162 62571 29196 62617
rect 28856 62531 29196 62571
rect 27387 62454 29196 62531
rect 27387 62413 29116 62454
rect 27387 62367 28810 62413
rect 28856 62408 29116 62413
rect 29162 62408 29196 62454
rect 28856 62367 29196 62408
rect 27387 62253 29196 62367
rect 30583 63020 30637 63066
rect 30683 63060 32842 63066
rect 34247 63060 35008 63067
rect 35182 63187 36364 63194
rect 35182 63153 36958 63187
rect 35182 63101 35220 63153
rect 35272 63101 35430 63153
rect 35482 63101 35641 63153
rect 35693 63101 35853 63153
rect 35905 63101 36064 63153
rect 36116 63101 36274 63153
rect 36326 63150 36958 63153
rect 36326 63104 36489 63150
rect 36723 63104 36958 63150
rect 36326 63101 36958 63104
rect 35182 63067 36958 63101
rect 37946 63153 38842 63194
rect 37946 63150 38330 63153
rect 38382 63150 38541 63153
rect 37946 63104 37957 63150
rect 38473 63104 38541 63150
rect 37946 63101 38330 63104
rect 38382 63101 38541 63104
rect 38593 63101 38752 63153
rect 38804 63101 38842 63153
rect 35182 63060 36364 63067
rect 37946 63060 38842 63101
rect 39014 63153 39323 63639
rect 39014 63101 39052 63153
rect 39104 63150 39232 63153
rect 39108 63104 39220 63150
rect 39104 63101 39232 63104
rect 39284 63101 39323 63153
rect 30683 63026 31040 63060
rect 30683 63020 30855 63026
rect 30583 62980 30855 63020
rect 30901 62980 31040 63026
rect 30583 62903 31040 62980
rect 33484 62984 33552 62995
rect 33019 62929 33327 62970
rect 33019 62926 33057 62929
rect 33109 62926 33237 62929
rect 33289 62926 33327 62929
rect 30583 62857 30637 62903
rect 30683 62862 31040 62903
rect 31336 62880 31349 62926
rect 33323 62880 33336 62926
rect 30683 62857 30855 62862
rect 30583 62816 30855 62857
rect 30901 62816 31040 62862
rect 33019 62877 33057 62880
rect 33109 62877 33237 62880
rect 33289 62877 33327 62880
rect 33019 62837 33327 62877
rect 30583 62740 31040 62816
rect 30583 62694 30637 62740
rect 30683 62724 31040 62740
rect 30683 62702 31493 62724
rect 30683 62699 31349 62702
rect 30683 62694 30855 62699
rect 30583 62653 30855 62694
rect 30901 62656 31349 62699
rect 33323 62656 33336 62702
rect 30901 62653 31493 62656
rect 30583 62605 31493 62653
rect 30583 62577 31040 62605
rect 30583 62531 30637 62577
rect 30683 62536 31040 62577
rect 30683 62531 30855 62536
rect 30583 62490 30855 62531
rect 30901 62490 31040 62536
rect 33484 62562 33495 62984
rect 33541 62562 33552 62984
rect 33781 62937 34089 62978
rect 33781 62926 33819 62937
rect 33871 62926 33999 62937
rect 34051 62926 34089 62937
rect 33671 62880 33684 62926
rect 33730 62880 33787 62926
rect 33871 62885 33890 62926
rect 33833 62880 33890 62885
rect 33936 62880 33993 62926
rect 34051 62885 34096 62926
rect 34039 62880 34096 62885
rect 34142 62880 34199 62926
rect 34245 62880 34302 62926
rect 34348 62880 34405 62926
rect 34451 62880 34508 62926
rect 34554 62880 34612 62926
rect 34658 62880 34671 62926
rect 33781 62845 34089 62880
rect 35294 62851 36266 62891
rect 37853 62888 38161 62904
rect 35294 62839 35332 62851
rect 35384 62839 35543 62851
rect 35595 62839 35754 62851
rect 35806 62839 35965 62851
rect 36017 62839 36176 62851
rect 36228 62839 36266 62851
rect 36438 62839 36953 62888
rect 37439 62863 38161 62888
rect 37439 62839 37891 62863
rect 37943 62839 38071 62863
rect 38123 62839 38161 62863
rect 35260 62793 35273 62839
rect 35523 62799 35543 62839
rect 35523 62793 35580 62799
rect 35626 62793 35683 62839
rect 35729 62799 35754 62839
rect 35729 62793 35786 62799
rect 35832 62793 35889 62839
rect 35935 62799 35965 62839
rect 35935 62793 35992 62799
rect 36038 62793 36095 62839
rect 36141 62799 36176 62839
rect 36141 62793 36198 62799
rect 36244 62793 36301 62839
rect 36347 62793 36360 62839
rect 36438 62793 36854 62839
rect 36900 62793 36971 62839
rect 37017 62793 37088 62839
rect 37134 62793 37206 62839
rect 37252 62793 37324 62839
rect 37370 62793 37442 62839
rect 37488 62811 37891 62839
rect 37488 62793 37909 62811
rect 37955 62793 38026 62839
rect 38123 62811 38143 62839
rect 38072 62793 38143 62811
rect 38189 62793 38261 62839
rect 38307 62793 38379 62839
rect 38425 62793 38497 62839
rect 38543 62793 38556 62839
rect 35294 62759 36266 62793
rect 36438 62768 36953 62793
rect 37439 62771 38161 62793
rect 37439 62768 37931 62771
rect 34228 62702 34718 62731
rect 33671 62656 33684 62702
rect 33730 62656 33787 62702
rect 33833 62656 33890 62702
rect 33936 62656 33993 62702
rect 34039 62656 34096 62702
rect 34142 62656 34199 62702
rect 34245 62691 34302 62702
rect 34245 62656 34267 62691
rect 34348 62656 34405 62702
rect 34451 62691 34508 62702
rect 34499 62656 34508 62691
rect 34554 62656 34612 62702
rect 34658 62691 34718 62702
rect 34228 62639 34267 62656
rect 34319 62639 34447 62656
rect 34499 62639 34627 62656
rect 34679 62639 34718 62691
rect 36438 62665 36554 62768
rect 34228 62598 34718 62639
rect 34964 62615 36360 62659
rect 30583 62413 31040 62490
rect 33019 62481 33327 62522
rect 33019 62478 33057 62481
rect 33109 62478 33237 62481
rect 33289 62478 33327 62481
rect 33484 62480 33552 62562
rect 34964 62569 35273 62615
rect 35523 62569 35580 62615
rect 35626 62569 35683 62615
rect 35729 62569 35786 62615
rect 35832 62569 35889 62615
rect 35935 62569 35992 62615
rect 36038 62569 36095 62615
rect 36141 62569 36198 62615
rect 36244 62569 36301 62615
rect 36347 62569 36360 62615
rect 34964 62537 36360 62569
rect 34964 62480 35082 62537
rect 31336 62432 31349 62478
rect 33323 62432 33336 62478
rect 33484 62443 35082 62480
rect 30583 62367 30637 62413
rect 30683 62373 31040 62413
rect 33019 62429 33057 62432
rect 33109 62429 33237 62432
rect 33289 62429 33327 62432
rect 33019 62389 33327 62429
rect 33484 62397 33816 62443
rect 33862 62397 34002 62443
rect 34048 62397 34189 62443
rect 34235 62397 34376 62443
rect 34422 62397 34562 62443
rect 34608 62397 35082 62443
rect 36438 62525 36475 62665
rect 36521 62525 36554 62665
rect 33484 62389 35082 62397
rect 35294 62391 36266 62431
rect 36438 62425 36554 62525
rect 36640 62665 36773 62688
rect 36640 62616 36697 62665
rect 36640 62564 36678 62616
rect 36640 62525 36697 62564
rect 36743 62525 36773 62665
rect 38658 62667 38726 62678
rect 36924 62657 37685 62663
rect 36923 62656 37685 62657
rect 36923 62623 37931 62656
rect 36923 62615 36961 62623
rect 37013 62615 37172 62623
rect 37224 62615 37384 62623
rect 36841 62569 36854 62615
rect 36900 62571 36961 62615
rect 36900 62569 36971 62571
rect 37017 62569 37088 62615
rect 37134 62571 37172 62615
rect 37134 62569 37206 62571
rect 37252 62569 37324 62615
rect 37370 62571 37384 62615
rect 37436 62615 37595 62623
rect 37436 62571 37442 62615
rect 37370 62569 37442 62571
rect 37488 62571 37595 62615
rect 37647 62615 37931 62623
rect 37647 62571 37909 62615
rect 37488 62569 37909 62571
rect 37955 62569 38026 62615
rect 38072 62569 38143 62615
rect 38189 62569 38261 62615
rect 38307 62569 38379 62615
rect 38425 62569 38497 62615
rect 38543 62569 38556 62615
rect 36923 62537 37931 62569
rect 36924 62530 37685 62537
rect 36640 62505 36773 62525
rect 38658 62527 38669 62667
rect 38715 62527 38726 62667
rect 39014 62615 39323 63101
rect 39492 63187 39608 63639
rect 39923 63606 40085 63737
rect 39923 63554 39994 63606
rect 40046 63554 40085 63606
rect 39923 63514 40085 63554
rect 39737 63418 39865 63431
rect 39737 63391 39866 63418
rect 39737 63374 39775 63391
rect 39827 63374 39866 63391
rect 39727 63328 39740 63374
rect 39827 63339 39862 63374
rect 39786 63328 39862 63339
rect 39908 63328 39985 63374
rect 40031 63328 40108 63374
rect 40154 63328 40167 63374
rect 40246 63363 40362 63761
rect 42229 63622 44509 63663
rect 42229 63570 42312 63622
rect 42364 63570 44509 63622
rect 42229 63530 44509 63570
rect 44341 63486 44509 63530
rect 44341 63440 44358 63486
rect 44498 63440 44509 63486
rect 39737 63299 39866 63328
rect 40246 63317 40281 63363
rect 40327 63317 40362 63363
rect 40246 63280 40362 63317
rect 40718 63391 43524 63432
rect 44341 63429 44509 63440
rect 40718 63339 41935 63391
rect 41987 63339 43524 63391
rect 40718 63298 43524 63339
rect 44605 63374 44721 63761
rect 45400 63731 48379 63772
rect 45400 63717 45975 63731
rect 45400 63671 45464 63717
rect 45604 63679 45975 63717
rect 46027 63679 48379 63731
rect 45604 63671 48379 63679
rect 44901 63615 45241 63656
rect 45400 63638 48379 63671
rect 48557 63725 48596 63777
rect 48648 63725 48687 63777
rect 48557 63702 48687 63725
rect 50044 63811 50516 63857
rect 50562 63811 50703 63857
rect 50749 63811 50890 63857
rect 50936 63811 51076 63857
rect 51122 63811 51263 63857
rect 51309 63811 51657 63857
rect 51797 63847 52105 63887
rect 51797 63822 51835 63847
rect 51887 63822 52015 63847
rect 52067 63822 52105 63847
rect 54085 63881 54223 63927
rect 54269 63887 54540 63927
rect 54269 63881 54440 63887
rect 54085 63841 54440 63881
rect 54486 63841 54540 63887
rect 50044 63774 51657 63811
rect 51789 63776 51802 63822
rect 53776 63776 53789 63822
rect 50044 63717 50160 63774
rect 44901 63598 44939 63615
rect 44991 63598 45151 63615
rect 45203 63598 45241 63615
rect 44799 63552 44812 63598
rect 44858 63552 44925 63598
rect 44991 63563 45038 63598
rect 44971 63552 45038 63563
rect 45084 63552 45151 63598
rect 45203 63563 45264 63598
rect 45197 63552 45264 63563
rect 45310 63552 45323 63598
rect 48557 63562 48622 63702
rect 48668 63562 48687 63702
rect 49820 63685 50160 63717
rect 48765 63639 48778 63685
rect 48824 63639 48881 63685
rect 48927 63639 48984 63685
rect 49030 63639 49087 63685
rect 49133 63639 49190 63685
rect 49236 63639 49293 63685
rect 49339 63639 49396 63685
rect 49442 63639 49499 63685
rect 49545 63639 49602 63685
rect 49852 63639 50160 63685
rect 51589 63722 51657 63774
rect 51797 63754 52105 63776
rect 49820 63598 50160 63639
rect 50262 63615 50812 63656
rect 48557 63559 48687 63562
rect 44901 63523 45241 63552
rect 48557 63507 48596 63559
rect 48648 63507 48687 63559
rect 50262 63563 50300 63615
rect 50352 63598 50511 63615
rect 50563 63598 50722 63615
rect 50352 63563 50467 63598
rect 50563 63563 50571 63598
rect 50262 63552 50467 63563
rect 50513 63552 50571 63563
rect 50617 63552 50674 63598
rect 50720 63563 50722 63598
rect 50774 63598 50812 63615
rect 50774 63563 50777 63598
rect 50720 63552 50777 63563
rect 50823 63552 50880 63598
rect 50926 63552 50983 63598
rect 51029 63552 51086 63598
rect 51132 63552 51189 63598
rect 51235 63552 51292 63598
rect 51338 63552 51395 63598
rect 51441 63552 51454 63598
rect 50262 63523 50812 63552
rect 48557 63466 48687 63507
rect 48905 63461 49877 63492
rect 48765 63415 48778 63461
rect 48824 63415 48881 63461
rect 48927 63452 48984 63461
rect 48927 63415 48943 63452
rect 49030 63415 49087 63461
rect 49133 63452 49190 63461
rect 49133 63415 49154 63452
rect 49236 63415 49293 63461
rect 49339 63452 49396 63461
rect 49339 63415 49365 63452
rect 49442 63415 49499 63461
rect 49545 63452 49602 63461
rect 49545 63415 49576 63452
rect 49852 63415 49877 63461
rect 48905 63400 48943 63415
rect 48995 63400 49154 63415
rect 49206 63400 49365 63415
rect 49417 63400 49576 63415
rect 49628 63400 49787 63415
rect 49839 63400 49877 63415
rect 44605 63328 44812 63374
rect 44858 63328 44925 63374
rect 44971 63328 45038 63374
rect 45084 63328 45151 63374
rect 45197 63328 45264 63374
rect 45310 63328 45323 63374
rect 48905 63360 49877 63400
rect 51035 63377 51343 63417
rect 51035 63374 51073 63377
rect 51125 63374 51253 63377
rect 51305 63374 51343 63377
rect 43362 63291 43524 63298
rect 43362 63245 43373 63291
rect 43513 63245 43524 63291
rect 43362 63234 43524 63245
rect 45584 63314 48546 63350
rect 50454 63328 50467 63374
rect 50513 63328 50571 63374
rect 50617 63328 50674 63374
rect 50720 63328 50777 63374
rect 50823 63328 50880 63374
rect 50926 63328 50983 63374
rect 51029 63328 51073 63374
rect 51132 63328 51189 63374
rect 51235 63328 51253 63374
rect 51338 63328 51395 63374
rect 51441 63328 51454 63374
rect 45584 63268 45619 63314
rect 45665 63268 45777 63314
rect 45823 63268 45935 63314
rect 45981 63268 46093 63314
rect 46139 63268 46251 63314
rect 46297 63268 46409 63314
rect 46455 63268 46568 63314
rect 46614 63268 46726 63314
rect 46772 63268 46884 63314
rect 46930 63268 47042 63314
rect 47088 63268 47200 63314
rect 47246 63268 47358 63314
rect 47404 63268 47516 63314
rect 47562 63268 47675 63314
rect 47721 63268 47833 63314
rect 47879 63268 47991 63314
rect 48037 63268 48149 63314
rect 48195 63268 48307 63314
rect 48353 63268 48465 63314
rect 48511 63268 48546 63314
rect 51035 63325 51073 63328
rect 51125 63325 51253 63328
rect 51305 63325 51343 63328
rect 51035 63284 51343 63325
rect 51589 63300 51600 63722
rect 51646 63300 51657 63722
rect 54085 63723 54540 63841
rect 54085 63677 54440 63723
rect 54486 63677 54540 63723
rect 54085 63649 54540 63677
rect 53585 63598 54540 63649
rect 51789 63552 51802 63598
rect 53776 63560 54540 63598
rect 53776 63552 54440 63560
rect 53585 63530 54440 63552
rect 54085 63514 54440 63530
rect 54486 63514 54540 63560
rect 54085 63438 54540 63514
rect 51797 63384 52105 63424
rect 51797 63374 51835 63384
rect 51887 63374 52015 63384
rect 52067 63374 52105 63384
rect 54085 63392 54223 63438
rect 54269 63397 54540 63438
rect 54269 63392 54440 63397
rect 51789 63328 51802 63374
rect 53776 63328 53789 63374
rect 54085 63351 54440 63392
rect 54486 63351 54540 63397
rect 51589 63289 51657 63300
rect 51797 63291 52105 63328
rect 40215 63187 40523 63194
rect 40788 63187 42986 63201
rect 43753 63187 44514 63194
rect 39492 63164 42986 63187
rect 43704 63164 44514 63187
rect 39492 63153 44514 63164
rect 39492 63150 40253 63153
rect 39492 63104 39740 63150
rect 39786 63104 39862 63150
rect 39908 63104 39985 63150
rect 40031 63104 40108 63150
rect 40154 63104 40253 63150
rect 39492 63101 40253 63104
rect 40305 63101 40433 63153
rect 40485 63150 43790 63153
rect 40485 63104 40836 63150
rect 40882 63104 40994 63150
rect 41040 63104 41152 63150
rect 41198 63104 41310 63150
rect 41356 63104 41469 63150
rect 41515 63104 41627 63150
rect 41673 63104 41785 63150
rect 41831 63104 41943 63150
rect 41989 63104 42101 63150
rect 42147 63104 42259 63150
rect 42305 63104 42418 63150
rect 42464 63104 42576 63150
rect 42622 63104 42734 63150
rect 42780 63104 42892 63150
rect 42938 63104 43739 63150
rect 43785 63104 43790 63150
rect 40485 63101 43790 63104
rect 43842 63150 44001 63153
rect 43842 63104 43906 63150
rect 43952 63104 44001 63150
rect 43842 63101 44001 63104
rect 44053 63150 44213 63153
rect 44265 63150 44424 63153
rect 44053 63104 44071 63150
rect 44117 63104 44213 63150
rect 44282 63104 44424 63150
rect 44053 63101 44213 63104
rect 44265 63101 44424 63104
rect 44476 63101 44514 63153
rect 39492 63090 44514 63101
rect 39492 63067 42986 63090
rect 43704 63067 44514 63090
rect 39492 62615 39608 63067
rect 40215 63060 40523 63067
rect 40788 63053 42986 63067
rect 43753 63060 44514 63067
rect 44796 63187 45346 63194
rect 45584 63187 48546 63268
rect 54085 63274 54540 63351
rect 54085 63228 54223 63274
rect 54269 63234 54540 63274
rect 54269 63228 54440 63234
rect 54085 63194 54440 63228
rect 48800 63187 49982 63194
rect 50308 63187 50859 63194
rect 44796 63153 49982 63187
rect 44796 63150 44834 63153
rect 44886 63150 45045 63153
rect 45097 63150 45256 63153
rect 45308 63150 48838 63153
rect 44796 63104 44812 63150
rect 44886 63104 44925 63150
rect 44971 63104 45038 63150
rect 45097 63104 45151 63150
rect 45197 63104 45256 63150
rect 45310 63104 45619 63150
rect 45665 63104 45777 63150
rect 45823 63104 45935 63150
rect 45981 63104 46093 63150
rect 46139 63104 46251 63150
rect 46297 63104 46409 63150
rect 46455 63104 46568 63150
rect 46614 63104 46726 63150
rect 46772 63104 46884 63150
rect 46930 63104 47042 63150
rect 47088 63104 47200 63150
rect 47246 63104 47358 63150
rect 47404 63104 47516 63150
rect 47562 63104 47675 63150
rect 47721 63104 47833 63150
rect 47879 63104 47991 63150
rect 48037 63104 48149 63150
rect 48195 63104 48307 63150
rect 48353 63104 48465 63150
rect 48511 63104 48838 63150
rect 44796 63101 44834 63104
rect 44886 63101 45045 63104
rect 45097 63101 45256 63104
rect 45308 63101 48838 63104
rect 48890 63101 49048 63153
rect 49100 63101 49259 63153
rect 49311 63101 49471 63153
rect 49523 63101 49682 63153
rect 49734 63101 49892 63153
rect 49944 63101 49982 63153
rect 44796 63067 49982 63101
rect 50307 63153 50859 63187
rect 50307 63101 50346 63153
rect 50398 63150 50557 63153
rect 50609 63150 50768 63153
rect 50820 63150 50859 63153
rect 52278 63188 54440 63194
rect 54486 63188 54540 63234
rect 55927 63887 57736 64001
rect 55927 63844 56267 63887
rect 55927 63798 55961 63844
rect 56007 63841 56267 63844
rect 56313 63841 57736 63887
rect 56007 63798 57736 63841
rect 55927 63723 57736 63798
rect 55927 63681 56267 63723
rect 55927 63635 55961 63681
rect 56007 63677 56267 63681
rect 56313 63677 57736 63723
rect 56007 63635 57736 63677
rect 55927 63560 57736 63635
rect 55927 63517 56267 63560
rect 55927 63471 55961 63517
rect 56007 63514 56267 63517
rect 56313 63514 57736 63560
rect 56007 63471 57736 63514
rect 55927 63397 57736 63471
rect 55927 63354 56267 63397
rect 55927 63308 55961 63354
rect 56007 63351 56267 63354
rect 56313 63351 57736 63397
rect 56007 63308 57736 63351
rect 55927 63234 57736 63308
rect 52278 63153 54540 63188
rect 52278 63150 52316 63153
rect 52368 63150 52527 63153
rect 52579 63150 52738 63153
rect 52790 63150 52948 63153
rect 53000 63150 53159 63153
rect 53211 63150 53371 63153
rect 53423 63150 53582 63153
rect 53634 63150 53792 63153
rect 50398 63104 50467 63150
rect 50513 63104 50557 63150
rect 50617 63104 50674 63150
rect 50720 63104 50768 63150
rect 50823 63104 50880 63150
rect 50926 63104 50983 63150
rect 51029 63104 51086 63150
rect 51132 63104 51189 63150
rect 51235 63104 51292 63150
rect 51338 63104 51395 63150
rect 51441 63104 51454 63150
rect 51789 63104 51802 63150
rect 53776 63104 53792 63150
rect 50398 63101 50557 63104
rect 50609 63101 50768 63104
rect 50820 63101 50859 63104
rect 50307 63067 50859 63101
rect 44796 63060 45346 63067
rect 43362 63009 43524 63020
rect 39737 62926 39866 62955
rect 40246 62937 40362 62974
rect 43362 62963 43373 63009
rect 43513 62963 43524 63009
rect 43362 62956 43524 62963
rect 39727 62880 39740 62926
rect 39786 62915 39862 62926
rect 39827 62880 39862 62915
rect 39908 62880 39985 62926
rect 40031 62880 40108 62926
rect 40154 62880 40167 62926
rect 40246 62891 40281 62937
rect 40327 62891 40362 62937
rect 39737 62863 39775 62880
rect 39827 62863 39866 62880
rect 39737 62836 39866 62863
rect 39737 62823 39865 62836
rect 39923 62700 40085 62740
rect 39923 62648 39994 62700
rect 40046 62648 40085 62700
rect 39008 62569 39021 62615
rect 39067 62569 39144 62615
rect 39190 62569 39267 62615
rect 39313 62569 39326 62615
rect 39492 62569 39641 62615
rect 39687 62569 39730 62615
rect 39014 62537 39323 62569
rect 39492 62537 39608 62569
rect 37853 62425 38161 62430
rect 36438 62391 36953 62425
rect 37439 62391 38161 62425
rect 38658 62405 38726 62527
rect 39923 62517 40085 62648
rect 39809 62514 40085 62517
rect 39809 62506 39994 62514
rect 39809 62460 39844 62506
rect 39890 62462 39994 62506
rect 40046 62493 40085 62514
rect 40246 62493 40362 62891
rect 40718 62915 43524 62956
rect 45584 62986 48546 63067
rect 48800 63060 49982 63067
rect 50308 63060 50859 63067
rect 52278 63101 52316 63104
rect 52368 63101 52527 63104
rect 52579 63101 52738 63104
rect 52790 63101 52948 63104
rect 53000 63101 53159 63104
rect 53211 63101 53371 63104
rect 53423 63101 53582 63104
rect 53634 63101 53792 63104
rect 53844 63101 54003 63153
rect 54055 63101 54214 63153
rect 54266 63101 54540 63153
rect 52278 63066 54540 63101
rect 52278 63060 54440 63066
rect 45584 62940 45619 62986
rect 45665 62940 45777 62986
rect 45823 62940 45935 62986
rect 45981 62940 46093 62986
rect 46139 62940 46251 62986
rect 46297 62940 46409 62986
rect 46455 62940 46568 62986
rect 46614 62940 46726 62986
rect 46772 62940 46884 62986
rect 46930 62940 47042 62986
rect 47088 62940 47200 62986
rect 47246 62940 47358 62986
rect 47404 62940 47516 62986
rect 47562 62940 47675 62986
rect 47721 62940 47833 62986
rect 47879 62940 47991 62986
rect 48037 62940 48149 62986
rect 48195 62940 48307 62986
rect 48353 62940 48465 62986
rect 48511 62940 48546 62986
rect 54085 63026 54440 63060
rect 54085 62980 54223 63026
rect 54269 63020 54440 63026
rect 54486 63020 54540 63066
rect 54758 63153 55840 63194
rect 54758 63150 54855 63153
rect 54758 63104 54793 63150
rect 54839 63104 54855 63150
rect 54758 63101 54855 63104
rect 54907 63150 55066 63153
rect 54907 63104 54956 63150
rect 55002 63104 55066 63150
rect 54907 63101 55066 63104
rect 55118 63150 55278 63153
rect 55330 63150 55489 63153
rect 55164 63104 55278 63150
rect 55330 63104 55439 63150
rect 55485 63104 55489 63150
rect 55118 63101 55278 63104
rect 55330 63101 55489 63104
rect 55541 63150 55840 63153
rect 55541 63104 55599 63150
rect 55645 63104 55760 63150
rect 55806 63104 55840 63150
rect 55541 63101 55840 63104
rect 54758 63061 55840 63101
rect 55927 63188 56267 63234
rect 56313 63188 57736 63234
rect 55927 63066 57736 63188
rect 54817 63060 55579 63061
rect 54269 62980 54540 63020
rect 40718 62863 41935 62915
rect 41987 62863 43524 62915
rect 40718 62822 43524 62863
rect 44605 62880 44812 62926
rect 44858 62880 44925 62926
rect 44971 62880 45038 62926
rect 45084 62880 45151 62926
rect 45197 62880 45264 62926
rect 45310 62880 45323 62926
rect 45584 62904 48546 62940
rect 51035 62929 51343 62970
rect 51035 62926 51073 62929
rect 51125 62926 51253 62929
rect 51305 62926 51343 62929
rect 51589 62954 51657 62965
rect 44341 62814 44509 62825
rect 44341 62768 44358 62814
rect 44498 62768 44509 62814
rect 44341 62724 44509 62768
rect 42229 62684 44509 62724
rect 42229 62632 42312 62684
rect 42364 62632 44509 62684
rect 42229 62591 44509 62632
rect 44605 62493 44721 62880
rect 48905 62854 49877 62894
rect 50454 62880 50467 62926
rect 50513 62880 50571 62926
rect 50617 62880 50674 62926
rect 50720 62880 50777 62926
rect 50823 62880 50880 62926
rect 50926 62880 50983 62926
rect 51029 62880 51073 62926
rect 51132 62880 51189 62926
rect 51235 62880 51253 62926
rect 51338 62880 51395 62926
rect 51441 62880 51454 62926
rect 48905 62839 48943 62854
rect 48995 62839 49154 62854
rect 49206 62839 49365 62854
rect 49417 62839 49576 62854
rect 49628 62839 49787 62854
rect 49839 62839 49877 62854
rect 48765 62793 48778 62839
rect 48824 62793 48881 62839
rect 48927 62802 48943 62839
rect 48927 62793 48984 62802
rect 49030 62793 49087 62839
rect 49133 62802 49154 62839
rect 49133 62793 49190 62802
rect 49236 62793 49293 62839
rect 49339 62802 49365 62839
rect 49339 62793 49396 62802
rect 49442 62793 49499 62839
rect 49545 62802 49576 62839
rect 49545 62793 49602 62802
rect 49852 62793 49877 62839
rect 51035 62877 51073 62880
rect 51125 62877 51253 62880
rect 51305 62877 51343 62880
rect 51035 62837 51343 62877
rect 48557 62747 48687 62788
rect 48905 62762 49877 62793
rect 44901 62702 45241 62731
rect 44799 62656 44812 62702
rect 44858 62656 44925 62702
rect 44971 62691 45038 62702
rect 44991 62656 45038 62691
rect 45084 62656 45151 62702
rect 45197 62691 45264 62702
rect 45203 62656 45264 62691
rect 45310 62656 45323 62702
rect 48557 62695 48596 62747
rect 48648 62695 48687 62747
rect 48557 62692 48687 62695
rect 44901 62639 44939 62656
rect 44991 62639 45151 62656
rect 45203 62639 45241 62656
rect 44901 62598 45241 62639
rect 45400 62583 48379 62616
rect 45400 62537 45464 62583
rect 45604 62575 48379 62583
rect 45604 62537 46353 62575
rect 45400 62523 46353 62537
rect 46405 62523 48379 62575
rect 40046 62478 44918 62493
rect 45400 62482 48379 62523
rect 48557 62552 48622 62692
rect 48668 62552 48687 62692
rect 50262 62702 50812 62731
rect 50262 62691 50467 62702
rect 50513 62691 50571 62702
rect 49820 62615 50160 62656
rect 48765 62569 48778 62615
rect 48824 62569 48881 62615
rect 48927 62569 48984 62615
rect 49030 62569 49087 62615
rect 49133 62569 49190 62615
rect 49236 62569 49293 62615
rect 49339 62569 49396 62615
rect 49442 62569 49499 62615
rect 49545 62569 49602 62615
rect 49852 62569 50160 62615
rect 50262 62639 50300 62691
rect 50352 62656 50467 62691
rect 50563 62656 50571 62691
rect 50617 62656 50674 62702
rect 50720 62691 50777 62702
rect 50720 62656 50722 62691
rect 50352 62639 50511 62656
rect 50563 62639 50722 62656
rect 50774 62656 50777 62691
rect 50823 62656 50880 62702
rect 50926 62656 50983 62702
rect 51029 62656 51086 62702
rect 51132 62656 51189 62702
rect 51235 62656 51292 62702
rect 51338 62656 51395 62702
rect 51441 62656 51454 62702
rect 50774 62639 50812 62656
rect 50262 62598 50812 62639
rect 48557 62529 48687 62552
rect 49820 62537 50160 62569
rect 40046 62462 44812 62478
rect 39890 62460 44812 62462
rect 39809 62457 44812 62460
rect 39809 62411 43739 62457
rect 43785 62411 43906 62457
rect 43952 62411 44071 62457
rect 44117 62411 44236 62457
rect 44282 62432 44812 62457
rect 44858 62432 44925 62478
rect 44971 62432 45038 62478
rect 45084 62432 45151 62478
rect 45197 62432 45264 62478
rect 45310 62432 45323 62478
rect 48557 62477 48596 62529
rect 48648 62477 48687 62529
rect 48557 62437 48687 62477
rect 50044 62480 50160 62537
rect 51589 62532 51600 62954
rect 51646 62532 51657 62954
rect 51797 62926 52105 62963
rect 51789 62880 51802 62926
rect 53776 62880 53789 62926
rect 54085 62903 54540 62980
rect 51797 62870 51835 62880
rect 51887 62870 52015 62880
rect 52067 62870 52105 62880
rect 51797 62830 52105 62870
rect 54085 62862 54440 62903
rect 54085 62816 54223 62862
rect 54269 62857 54440 62862
rect 54486 62857 54540 62903
rect 54269 62816 54540 62857
rect 54085 62740 54540 62816
rect 54085 62724 54440 62740
rect 53585 62702 54440 62724
rect 51789 62656 51802 62702
rect 53776 62694 54440 62702
rect 54486 62694 54540 62740
rect 53776 62656 54540 62694
rect 53585 62605 54540 62656
rect 51589 62480 51657 62532
rect 54085 62577 54540 62605
rect 54085 62531 54440 62577
rect 54486 62531 54540 62577
rect 50044 62443 51657 62480
rect 51797 62478 52105 62500
rect 44282 62411 44918 62432
rect 38658 62391 39723 62405
rect 30683 62367 30855 62373
rect 30583 62327 30855 62367
rect 30901 62327 31040 62373
rect 33484 62360 34643 62389
rect 35260 62345 35273 62391
rect 35523 62345 35543 62391
rect 35626 62345 35683 62391
rect 35729 62345 35754 62391
rect 35832 62345 35889 62391
rect 35935 62345 35965 62391
rect 36038 62345 36095 62391
rect 36141 62345 36176 62391
rect 36244 62345 36301 62391
rect 36347 62345 36360 62391
rect 36438 62345 36854 62391
rect 36900 62345 36971 62391
rect 37017 62345 37088 62391
rect 37134 62345 37206 62391
rect 37252 62345 37324 62391
rect 37370 62345 37442 62391
rect 37488 62389 37909 62391
rect 37488 62345 37891 62389
rect 37955 62345 38026 62391
rect 38072 62389 38143 62391
rect 38123 62345 38143 62389
rect 38189 62345 38261 62391
rect 38307 62345 38379 62391
rect 38425 62345 38497 62391
rect 38543 62345 38556 62391
rect 38658 62345 39021 62391
rect 39067 62345 39144 62391
rect 39190 62345 39267 62391
rect 39313 62345 39641 62391
rect 39687 62345 39730 62391
rect 39809 62373 44918 62411
rect 48905 62391 49877 62431
rect 48765 62345 48778 62391
rect 48824 62345 48881 62391
rect 48927 62345 48943 62391
rect 49030 62345 49087 62391
rect 49133 62345 49154 62391
rect 49236 62345 49293 62391
rect 49339 62345 49365 62391
rect 49442 62345 49499 62391
rect 49545 62345 49576 62391
rect 49852 62345 49877 62391
rect 50044 62397 50516 62443
rect 50562 62397 50703 62443
rect 50749 62397 50890 62443
rect 50936 62397 51076 62443
rect 51122 62397 51263 62443
rect 51309 62397 51657 62443
rect 51789 62432 51802 62478
rect 53776 62432 53789 62478
rect 50044 62387 51657 62397
rect 50481 62360 51657 62387
rect 51797 62407 51835 62432
rect 51887 62407 52015 62432
rect 52067 62407 52105 62432
rect 51797 62367 52105 62407
rect 54085 62413 54540 62531
rect 54085 62373 54440 62413
rect 30583 62294 31040 62327
rect 35294 62339 35332 62345
rect 35384 62339 35543 62345
rect 35595 62339 35754 62345
rect 35806 62339 35965 62345
rect 36017 62339 36176 62345
rect 36228 62339 36266 62345
rect 34870 62294 35025 62301
rect 35294 62299 36266 62339
rect 36438 62305 36953 62345
rect 37439 62337 37891 62345
rect 37943 62337 38071 62345
rect 38123 62337 38161 62345
rect 37439 62305 38161 62337
rect 37853 62297 38161 62305
rect 27387 62201 27790 62253
rect 27842 62201 28001 62253
rect 28053 62201 28212 62253
rect 28264 62201 28423 62253
rect 28475 62201 28634 62253
rect 28686 62250 28845 62253
rect 28686 62204 28810 62250
rect 28686 62201 28845 62204
rect 28897 62201 29056 62253
rect 29108 62201 29196 62253
rect 27387 62087 29196 62201
rect 29283 62253 30365 62294
rect 29283 62250 29582 62253
rect 29283 62204 29317 62250
rect 29363 62204 29478 62250
rect 29524 62204 29582 62250
rect 29283 62201 29582 62204
rect 29634 62250 29793 62253
rect 29845 62250 30005 62253
rect 29634 62204 29638 62250
rect 29684 62204 29793 62250
rect 29845 62204 29959 62250
rect 29634 62201 29793 62204
rect 29845 62201 30005 62204
rect 30057 62250 30216 62253
rect 30057 62204 30121 62250
rect 30167 62204 30216 62250
rect 30057 62201 30216 62204
rect 30268 62250 30365 62253
rect 30268 62204 30284 62250
rect 30330 62204 30365 62250
rect 30268 62201 30365 62204
rect 29283 62161 30365 62201
rect 30583 62253 32842 62294
rect 30583 62250 30854 62253
rect 30583 62204 30637 62250
rect 30683 62204 30854 62250
rect 30583 62201 30854 62204
rect 30906 62201 31065 62253
rect 31117 62201 31276 62253
rect 31328 62201 31486 62253
rect 31538 62201 31697 62253
rect 31749 62201 31909 62253
rect 31961 62201 32120 62253
rect 32172 62201 32330 62253
rect 32382 62201 32541 62253
rect 32593 62201 32752 62253
rect 32804 62201 32842 62253
rect 29544 62160 30306 62161
rect 30583 62160 32842 62201
rect 34717 62253 35025 62294
rect 38658 62285 39723 62345
rect 48905 62339 48943 62345
rect 48995 62339 49154 62345
rect 49206 62339 49365 62345
rect 49417 62339 49576 62345
rect 49628 62339 49787 62345
rect 49839 62339 49877 62345
rect 48905 62299 49877 62339
rect 54085 62327 54223 62373
rect 54269 62367 54440 62373
rect 54486 62367 54540 62413
rect 54269 62327 54540 62367
rect 50099 62294 50255 62301
rect 54085 62294 54540 62327
rect 55927 63020 56267 63066
rect 56313 63020 57736 63066
rect 55927 62944 57736 63020
rect 55927 62898 55961 62944
rect 56007 62903 57736 62944
rect 56007 62898 56267 62903
rect 55927 62857 56267 62898
rect 56313 62857 57736 62903
rect 55927 62781 57736 62857
rect 55927 62735 55961 62781
rect 56007 62740 57736 62781
rect 56007 62735 56267 62740
rect 55927 62694 56267 62735
rect 56313 62694 57736 62740
rect 55927 62617 57736 62694
rect 55927 62571 55961 62617
rect 56007 62577 57736 62617
rect 56007 62571 56267 62577
rect 55927 62531 56267 62571
rect 56313 62531 57736 62577
rect 55927 62454 57736 62531
rect 55927 62408 55961 62454
rect 56007 62413 57736 62454
rect 56007 62408 56267 62413
rect 55927 62367 56267 62408
rect 56313 62367 57736 62413
rect 34717 62201 34755 62253
rect 34807 62250 34935 62253
rect 34807 62204 34916 62250
rect 34807 62201 34935 62204
rect 34987 62201 35025 62253
rect 34717 62160 35025 62201
rect 50099 62253 50408 62294
rect 50099 62201 50138 62253
rect 50190 62250 50318 62253
rect 50206 62204 50318 62250
rect 50190 62201 50318 62204
rect 50370 62201 50408 62253
rect 27387 62041 28810 62087
rect 28856 62044 29196 62087
rect 28856 62041 29116 62044
rect 27387 61998 29116 62041
rect 29162 61998 29196 62044
rect 27387 61923 29196 61998
rect 27387 61877 28810 61923
rect 28856 61881 29196 61923
rect 28856 61877 29116 61881
rect 27387 61835 29116 61877
rect 29162 61835 29196 61881
rect 27387 61760 29196 61835
rect 27387 61714 28810 61760
rect 28856 61717 29196 61760
rect 28856 61714 29116 61717
rect 27387 61671 29116 61714
rect 29162 61671 29196 61717
rect 27387 61597 29196 61671
rect 27387 61551 28810 61597
rect 28856 61554 29196 61597
rect 28856 61551 29116 61554
rect 27387 61508 29116 61551
rect 29162 61508 29196 61554
rect 27387 61434 29196 61508
rect 27387 61388 28810 61434
rect 28856 61388 29196 61434
rect 30583 62127 31040 62160
rect 34870 62153 35025 62160
rect 30583 62087 30855 62127
rect 30583 62041 30637 62087
rect 30683 62081 30855 62087
rect 30901 62081 31040 62127
rect 35294 62115 36266 62155
rect 37853 62149 38161 62157
rect 35294 62109 35332 62115
rect 35384 62109 35543 62115
rect 35595 62109 35754 62115
rect 35806 62109 35965 62115
rect 36017 62109 36176 62115
rect 36228 62109 36266 62115
rect 36438 62109 36953 62149
rect 37439 62117 38161 62149
rect 37439 62109 37891 62117
rect 37943 62109 38071 62117
rect 38123 62109 38161 62117
rect 38658 62109 39723 62169
rect 50099 62160 50408 62201
rect 52278 62253 54540 62294
rect 52278 62201 52316 62253
rect 52368 62201 52527 62253
rect 52579 62201 52738 62253
rect 52790 62201 52948 62253
rect 53000 62201 53159 62253
rect 53211 62201 53371 62253
rect 53423 62201 53582 62253
rect 53634 62201 53792 62253
rect 53844 62201 54003 62253
rect 54055 62201 54214 62253
rect 54266 62250 54540 62253
rect 54266 62204 54440 62250
rect 54486 62204 54540 62250
rect 54266 62201 54540 62204
rect 52278 62160 54540 62201
rect 54758 62253 55840 62294
rect 54758 62250 54855 62253
rect 54758 62204 54793 62250
rect 54839 62204 54855 62250
rect 54758 62201 54855 62204
rect 54907 62250 55066 62253
rect 54907 62204 54956 62250
rect 55002 62204 55066 62250
rect 54907 62201 55066 62204
rect 55118 62250 55278 62253
rect 55330 62250 55489 62253
rect 55164 62204 55278 62250
rect 55330 62204 55439 62250
rect 55485 62204 55489 62250
rect 55118 62201 55278 62204
rect 55330 62201 55489 62204
rect 55541 62250 55840 62253
rect 55541 62204 55599 62250
rect 55645 62204 55760 62250
rect 55806 62204 55840 62250
rect 55541 62201 55840 62204
rect 54758 62161 55840 62201
rect 55927 62253 57736 62367
rect 55927 62201 56015 62253
rect 56067 62201 56226 62253
rect 56278 62250 56437 62253
rect 56313 62204 56437 62250
rect 56278 62201 56437 62204
rect 56489 62201 56648 62253
rect 56700 62201 56859 62253
rect 56911 62201 57070 62253
rect 57122 62201 57281 62253
rect 57333 62201 57736 62253
rect 54817 62160 55579 62161
rect 48905 62115 49877 62155
rect 50099 62153 50255 62160
rect 48905 62109 48943 62115
rect 48995 62109 49154 62115
rect 49206 62109 49365 62115
rect 49417 62109 49576 62115
rect 49628 62109 49787 62115
rect 49839 62109 49877 62115
rect 30683 62041 31040 62081
rect 33484 62065 34643 62094
rect 30583 61964 31040 62041
rect 33019 62025 33327 62065
rect 33019 62022 33057 62025
rect 33109 62022 33237 62025
rect 33289 62022 33327 62025
rect 33484 62057 35082 62065
rect 35260 62063 35273 62109
rect 35523 62063 35543 62109
rect 35626 62063 35683 62109
rect 35729 62063 35754 62109
rect 35832 62063 35889 62109
rect 35935 62063 35965 62109
rect 36038 62063 36095 62109
rect 36141 62063 36176 62109
rect 36244 62063 36301 62109
rect 36347 62063 36360 62109
rect 36438 62063 36854 62109
rect 36900 62063 36971 62109
rect 37017 62063 37088 62109
rect 37134 62063 37206 62109
rect 37252 62063 37324 62109
rect 37370 62063 37442 62109
rect 37488 62065 37891 62109
rect 37488 62063 37909 62065
rect 37955 62063 38026 62109
rect 38123 62065 38143 62109
rect 38072 62063 38143 62065
rect 38189 62063 38261 62109
rect 38307 62063 38379 62109
rect 38425 62063 38497 62109
rect 38543 62063 38556 62109
rect 38658 62063 39021 62109
rect 39067 62063 39144 62109
rect 39190 62063 39267 62109
rect 39313 62063 39641 62109
rect 39687 62063 39730 62109
rect 31336 61976 31349 62022
rect 33323 61976 33336 62022
rect 33484 62011 33816 62057
rect 33862 62011 34002 62057
rect 34048 62011 34189 62057
rect 34235 62011 34376 62057
rect 34422 62011 34562 62057
rect 34608 62011 35082 62057
rect 35294 62023 36266 62063
rect 36438 62029 36953 62063
rect 37439 62029 38161 62063
rect 30583 61923 30855 61964
rect 30583 61877 30637 61923
rect 30683 61918 30855 61923
rect 30901 61918 31040 61964
rect 33019 61973 33057 61976
rect 33109 61973 33237 61976
rect 33289 61973 33327 61976
rect 33019 61932 33327 61973
rect 33484 61974 35082 62011
rect 30683 61877 31040 61918
rect 30583 61849 31040 61877
rect 33484 61892 33552 61974
rect 30583 61801 31493 61849
rect 30583 61760 30855 61801
rect 30583 61714 30637 61760
rect 30683 61755 30855 61760
rect 30901 61798 31493 61801
rect 30901 61755 31349 61798
rect 30683 61752 31349 61755
rect 33323 61752 33336 61798
rect 30683 61730 31493 61752
rect 30683 61714 31040 61730
rect 30583 61638 31040 61714
rect 30583 61597 30855 61638
rect 30583 61551 30637 61597
rect 30683 61592 30855 61597
rect 30901 61592 31040 61638
rect 30683 61551 31040 61592
rect 33019 61577 33327 61617
rect 33019 61574 33057 61577
rect 33109 61574 33237 61577
rect 33289 61574 33327 61577
rect 30583 61474 31040 61551
rect 31336 61528 31349 61574
rect 33323 61528 33336 61574
rect 33019 61525 33057 61528
rect 33109 61525 33237 61528
rect 33289 61525 33327 61528
rect 33019 61484 33327 61525
rect 30583 61434 30855 61474
rect 27387 61266 29196 61388
rect 27387 61220 28810 61266
rect 28856 61220 29196 61266
rect 29283 61353 30365 61394
rect 29283 61350 29582 61353
rect 29283 61304 29317 61350
rect 29363 61304 29478 61350
rect 29524 61304 29582 61350
rect 29283 61301 29582 61304
rect 29634 61350 29793 61353
rect 29845 61350 30005 61353
rect 29634 61304 29638 61350
rect 29684 61304 29793 61350
rect 29845 61304 29959 61350
rect 29634 61301 29793 61304
rect 29845 61301 30005 61304
rect 30057 61350 30216 61353
rect 30057 61304 30121 61350
rect 30167 61304 30216 61350
rect 30057 61301 30216 61304
rect 30268 61350 30365 61353
rect 30268 61304 30284 61350
rect 30330 61304 30365 61350
rect 30268 61301 30365 61304
rect 29283 61261 30365 61301
rect 30583 61388 30637 61434
rect 30683 61428 30855 61434
rect 30901 61428 31040 61474
rect 33484 61470 33495 61892
rect 33541 61470 33552 61892
rect 34964 61917 35082 61974
rect 36438 61929 36554 62029
rect 37853 62024 38161 62029
rect 38658 62049 39723 62063
rect 34964 61885 36360 61917
rect 34228 61815 34718 61856
rect 34228 61798 34267 61815
rect 34319 61798 34447 61815
rect 34499 61798 34627 61815
rect 33671 61752 33684 61798
rect 33730 61752 33787 61798
rect 33833 61752 33890 61798
rect 33936 61752 33993 61798
rect 34039 61752 34096 61798
rect 34142 61752 34199 61798
rect 34245 61763 34267 61798
rect 34245 61752 34302 61763
rect 34348 61752 34405 61798
rect 34499 61763 34508 61798
rect 34451 61752 34508 61763
rect 34554 61752 34612 61798
rect 34679 61763 34718 61815
rect 34964 61839 35273 61885
rect 35523 61839 35580 61885
rect 35626 61839 35683 61885
rect 35729 61839 35786 61885
rect 35832 61839 35889 61885
rect 35935 61839 35992 61885
rect 36038 61839 36095 61885
rect 36141 61839 36198 61885
rect 36244 61839 36301 61885
rect 36347 61839 36360 61885
rect 34964 61795 36360 61839
rect 34658 61752 34718 61763
rect 34228 61723 34718 61752
rect 36438 61789 36475 61929
rect 36521 61789 36554 61929
rect 35294 61661 36266 61695
rect 36438 61686 36554 61789
rect 36640 61929 36773 61949
rect 36640 61890 36697 61929
rect 36640 61838 36678 61890
rect 36640 61789 36697 61838
rect 36743 61789 36773 61929
rect 38658 61927 38726 62049
rect 39809 62043 44918 62081
rect 48765 62063 48778 62109
rect 48824 62063 48881 62109
rect 48927 62063 48943 62109
rect 49030 62063 49087 62109
rect 49133 62063 49154 62109
rect 49236 62063 49293 62109
rect 49339 62063 49365 62109
rect 49442 62063 49499 62109
rect 49545 62063 49576 62109
rect 49852 62063 49877 62109
rect 54085 62127 54540 62160
rect 50481 62067 51657 62094
rect 39809 61997 43739 62043
rect 43785 61997 43906 62043
rect 43952 61997 44071 62043
rect 44117 61997 44236 62043
rect 44282 62022 44918 62043
rect 48905 62023 49877 62063
rect 50044 62057 51657 62067
rect 44282 61997 44812 62022
rect 39809 61994 44812 61997
rect 39809 61948 39844 61994
rect 39890 61992 44812 61994
rect 39890 61948 39994 61992
rect 39809 61940 39994 61948
rect 40046 61976 44812 61992
rect 44858 61976 44925 62022
rect 44971 61976 45038 62022
rect 45084 61976 45151 62022
rect 45197 61976 45264 62022
rect 45310 61976 45323 62022
rect 48557 61977 48687 62017
rect 40046 61961 44918 61976
rect 40046 61940 40085 61961
rect 39809 61937 40085 61940
rect 36924 61917 37685 61924
rect 36923 61885 37931 61917
rect 36841 61839 36854 61885
rect 36900 61883 36971 61885
rect 36900 61839 36961 61883
rect 37017 61839 37088 61885
rect 37134 61883 37206 61885
rect 37134 61839 37172 61883
rect 37252 61839 37324 61885
rect 37370 61883 37442 61885
rect 37370 61839 37384 61883
rect 36923 61831 36961 61839
rect 37013 61831 37172 61839
rect 37224 61831 37384 61839
rect 37436 61839 37442 61883
rect 37488 61883 37909 61885
rect 37488 61839 37595 61883
rect 37436 61831 37595 61839
rect 37647 61839 37909 61883
rect 37955 61839 38026 61885
rect 38072 61839 38143 61885
rect 38189 61839 38261 61885
rect 38307 61839 38379 61885
rect 38425 61839 38497 61885
rect 38543 61839 38556 61885
rect 37647 61831 37931 61839
rect 36923 61798 37931 61831
rect 36923 61797 37685 61798
rect 36924 61791 37685 61797
rect 36640 61766 36773 61789
rect 38658 61787 38669 61927
rect 38715 61787 38726 61927
rect 39014 61885 39323 61917
rect 39492 61885 39608 61917
rect 39008 61839 39021 61885
rect 39067 61839 39144 61885
rect 39190 61839 39267 61885
rect 39313 61839 39326 61885
rect 39492 61839 39641 61885
rect 39687 61839 39730 61885
rect 38658 61776 38726 61787
rect 36438 61661 36953 61686
rect 37439 61683 37931 61686
rect 37439 61661 38161 61683
rect 35260 61615 35273 61661
rect 35523 61655 35580 61661
rect 35523 61615 35543 61655
rect 35626 61615 35683 61661
rect 35729 61655 35786 61661
rect 35729 61615 35754 61655
rect 35832 61615 35889 61661
rect 35935 61655 35992 61661
rect 35935 61615 35965 61655
rect 36038 61615 36095 61661
rect 36141 61655 36198 61661
rect 36141 61615 36176 61655
rect 36244 61615 36301 61661
rect 36347 61615 36360 61661
rect 36438 61615 36854 61661
rect 36900 61615 36971 61661
rect 37017 61615 37088 61661
rect 37134 61615 37206 61661
rect 37252 61615 37324 61661
rect 37370 61615 37442 61661
rect 37488 61643 37909 61661
rect 37488 61615 37891 61643
rect 37955 61615 38026 61661
rect 38072 61643 38143 61661
rect 38123 61615 38143 61643
rect 38189 61615 38261 61661
rect 38307 61615 38379 61661
rect 38425 61615 38497 61661
rect 38543 61615 38556 61661
rect 33781 61574 34089 61609
rect 35294 61603 35332 61615
rect 35384 61603 35543 61615
rect 35595 61603 35754 61615
rect 35806 61603 35965 61615
rect 36017 61603 36176 61615
rect 36228 61603 36266 61615
rect 33671 61528 33684 61574
rect 33730 61528 33787 61574
rect 33833 61569 33890 61574
rect 33871 61528 33890 61569
rect 33936 61528 33993 61574
rect 34039 61569 34096 61574
rect 34051 61528 34096 61569
rect 34142 61528 34199 61574
rect 34245 61528 34302 61574
rect 34348 61528 34405 61574
rect 34451 61528 34508 61574
rect 34554 61528 34612 61574
rect 34658 61528 34671 61574
rect 35294 61563 36266 61603
rect 36438 61566 36953 61615
rect 37439 61591 37891 61615
rect 37943 61591 38071 61615
rect 38123 61591 38161 61615
rect 37439 61566 38161 61591
rect 37853 61550 38161 61566
rect 33781 61517 33819 61528
rect 33871 61517 33999 61528
rect 34051 61517 34089 61528
rect 33781 61476 34089 61517
rect 33484 61459 33552 61470
rect 30683 61394 31040 61428
rect 30683 61388 32842 61394
rect 30583 61353 32842 61388
rect 34247 61387 35008 61394
rect 30583 61301 30854 61353
rect 30906 61301 31065 61353
rect 31117 61301 31276 61353
rect 31328 61350 31486 61353
rect 31538 61350 31697 61353
rect 31749 61350 31909 61353
rect 31961 61350 32120 61353
rect 32172 61350 32330 61353
rect 32382 61350 32541 61353
rect 32593 61350 32752 61353
rect 32804 61350 32842 61353
rect 34246 61353 35008 61387
rect 34246 61350 34284 61353
rect 34336 61350 34495 61353
rect 34547 61350 34707 61353
rect 31328 61304 31349 61350
rect 33323 61304 33336 61350
rect 33671 61304 33684 61350
rect 33730 61304 33787 61350
rect 33833 61304 33890 61350
rect 33936 61304 33993 61350
rect 34039 61304 34096 61350
rect 34142 61304 34199 61350
rect 34245 61304 34284 61350
rect 34348 61304 34405 61350
rect 34451 61304 34495 61350
rect 34554 61304 34612 61350
rect 34658 61304 34707 61350
rect 31328 61301 31486 61304
rect 31538 61301 31697 61304
rect 31749 61301 31909 61304
rect 31961 61301 32120 61304
rect 32172 61301 32330 61304
rect 32382 61301 32541 61304
rect 32593 61301 32752 61304
rect 32804 61301 32842 61304
rect 30583 61266 32842 61301
rect 34246 61301 34284 61304
rect 34336 61301 34495 61304
rect 34547 61301 34707 61304
rect 34759 61301 34918 61353
rect 34970 61301 35008 61353
rect 34246 61267 35008 61301
rect 29544 61260 30306 61261
rect 27387 61144 29196 61220
rect 27387 61103 29116 61144
rect 27387 61057 28810 61103
rect 28856 61098 29116 61103
rect 29162 61098 29196 61144
rect 28856 61057 29196 61098
rect 27387 60981 29196 61057
rect 27387 60940 29116 60981
rect 27387 60894 28810 60940
rect 28856 60935 29116 60940
rect 29162 60935 29196 60981
rect 28856 60894 29196 60935
rect 27387 60817 29196 60894
rect 27387 60777 29116 60817
rect 27387 60731 28810 60777
rect 28856 60771 29116 60777
rect 29162 60771 29196 60817
rect 28856 60731 29196 60771
rect 27387 60654 29196 60731
rect 27387 60613 29116 60654
rect 27387 60567 28810 60613
rect 28856 60608 29116 60613
rect 29162 60608 29196 60654
rect 28856 60567 29196 60608
rect 27387 60453 29196 60567
rect 30583 61220 30637 61266
rect 30683 61260 32842 61266
rect 34247 61260 35008 61267
rect 35182 61387 36364 61394
rect 35182 61353 36958 61387
rect 35182 61301 35220 61353
rect 35272 61301 35430 61353
rect 35482 61301 35641 61353
rect 35693 61301 35853 61353
rect 35905 61301 36064 61353
rect 36116 61301 36274 61353
rect 36326 61350 36958 61353
rect 36326 61304 36489 61350
rect 36723 61304 36958 61350
rect 36326 61301 36958 61304
rect 35182 61267 36958 61301
rect 37946 61353 38842 61394
rect 37946 61350 38330 61353
rect 38382 61350 38541 61353
rect 37946 61304 37957 61350
rect 38473 61304 38541 61350
rect 37946 61301 38330 61304
rect 38382 61301 38541 61304
rect 38593 61301 38752 61353
rect 38804 61301 38842 61353
rect 35182 61260 36364 61267
rect 37946 61260 38842 61301
rect 39014 61353 39323 61839
rect 39014 61301 39052 61353
rect 39104 61350 39232 61353
rect 39108 61304 39220 61350
rect 39104 61301 39232 61304
rect 39284 61301 39323 61353
rect 30683 61226 31040 61260
rect 30683 61220 30855 61226
rect 30583 61180 30855 61220
rect 30901 61180 31040 61226
rect 30583 61103 31040 61180
rect 33484 61184 33552 61195
rect 33019 61129 33327 61170
rect 33019 61126 33057 61129
rect 33109 61126 33237 61129
rect 33289 61126 33327 61129
rect 30583 61057 30637 61103
rect 30683 61062 31040 61103
rect 31336 61080 31349 61126
rect 33323 61080 33336 61126
rect 30683 61057 30855 61062
rect 30583 61016 30855 61057
rect 30901 61016 31040 61062
rect 33019 61077 33057 61080
rect 33109 61077 33237 61080
rect 33289 61077 33327 61080
rect 33019 61037 33327 61077
rect 30583 60940 31040 61016
rect 30583 60894 30637 60940
rect 30683 60924 31040 60940
rect 30683 60902 31493 60924
rect 30683 60899 31349 60902
rect 30683 60894 30855 60899
rect 30583 60853 30855 60894
rect 30901 60856 31349 60899
rect 33323 60856 33336 60902
rect 30901 60853 31493 60856
rect 30583 60805 31493 60853
rect 30583 60777 31040 60805
rect 30583 60731 30637 60777
rect 30683 60736 31040 60777
rect 30683 60731 30855 60736
rect 30583 60690 30855 60731
rect 30901 60690 31040 60736
rect 33484 60762 33495 61184
rect 33541 60762 33552 61184
rect 33781 61137 34089 61178
rect 33781 61126 33819 61137
rect 33871 61126 33999 61137
rect 34051 61126 34089 61137
rect 33671 61080 33684 61126
rect 33730 61080 33787 61126
rect 33871 61085 33890 61126
rect 33833 61080 33890 61085
rect 33936 61080 33993 61126
rect 34051 61085 34096 61126
rect 34039 61080 34096 61085
rect 34142 61080 34199 61126
rect 34245 61080 34302 61126
rect 34348 61080 34405 61126
rect 34451 61080 34508 61126
rect 34554 61080 34612 61126
rect 34658 61080 34671 61126
rect 33781 61045 34089 61080
rect 35294 61051 36266 61091
rect 37853 61088 38161 61104
rect 35294 61039 35332 61051
rect 35384 61039 35543 61051
rect 35595 61039 35754 61051
rect 35806 61039 35965 61051
rect 36017 61039 36176 61051
rect 36228 61039 36266 61051
rect 36438 61039 36953 61088
rect 37439 61063 38161 61088
rect 37439 61039 37891 61063
rect 37943 61039 38071 61063
rect 38123 61039 38161 61063
rect 35260 60993 35273 61039
rect 35523 60999 35543 61039
rect 35523 60993 35580 60999
rect 35626 60993 35683 61039
rect 35729 60999 35754 61039
rect 35729 60993 35786 60999
rect 35832 60993 35889 61039
rect 35935 60999 35965 61039
rect 35935 60993 35992 60999
rect 36038 60993 36095 61039
rect 36141 60999 36176 61039
rect 36141 60993 36198 60999
rect 36244 60993 36301 61039
rect 36347 60993 36360 61039
rect 36438 60993 36854 61039
rect 36900 60993 36971 61039
rect 37017 60993 37088 61039
rect 37134 60993 37206 61039
rect 37252 60993 37324 61039
rect 37370 60993 37442 61039
rect 37488 61011 37891 61039
rect 37488 60993 37909 61011
rect 37955 60993 38026 61039
rect 38123 61011 38143 61039
rect 38072 60993 38143 61011
rect 38189 60993 38261 61039
rect 38307 60993 38379 61039
rect 38425 60993 38497 61039
rect 38543 60993 38556 61039
rect 35294 60959 36266 60993
rect 36438 60968 36953 60993
rect 37439 60971 38161 60993
rect 37439 60968 37931 60971
rect 34228 60902 34718 60931
rect 33671 60856 33684 60902
rect 33730 60856 33787 60902
rect 33833 60856 33890 60902
rect 33936 60856 33993 60902
rect 34039 60856 34096 60902
rect 34142 60856 34199 60902
rect 34245 60891 34302 60902
rect 34245 60856 34267 60891
rect 34348 60856 34405 60902
rect 34451 60891 34508 60902
rect 34499 60856 34508 60891
rect 34554 60856 34612 60902
rect 34658 60891 34718 60902
rect 34228 60839 34267 60856
rect 34319 60839 34447 60856
rect 34499 60839 34627 60856
rect 34679 60839 34718 60891
rect 36438 60865 36554 60968
rect 34228 60798 34718 60839
rect 34964 60815 36360 60859
rect 30583 60613 31040 60690
rect 33019 60681 33327 60722
rect 33019 60678 33057 60681
rect 33109 60678 33237 60681
rect 33289 60678 33327 60681
rect 33484 60680 33552 60762
rect 34964 60769 35273 60815
rect 35523 60769 35580 60815
rect 35626 60769 35683 60815
rect 35729 60769 35786 60815
rect 35832 60769 35889 60815
rect 35935 60769 35992 60815
rect 36038 60769 36095 60815
rect 36141 60769 36198 60815
rect 36244 60769 36301 60815
rect 36347 60769 36360 60815
rect 34964 60737 36360 60769
rect 34964 60680 35082 60737
rect 31336 60632 31349 60678
rect 33323 60632 33336 60678
rect 33484 60643 35082 60680
rect 30583 60567 30637 60613
rect 30683 60573 31040 60613
rect 33019 60629 33057 60632
rect 33109 60629 33237 60632
rect 33289 60629 33327 60632
rect 33019 60589 33327 60629
rect 33484 60597 33816 60643
rect 33862 60597 34002 60643
rect 34048 60597 34189 60643
rect 34235 60597 34376 60643
rect 34422 60597 34562 60643
rect 34608 60597 35082 60643
rect 36438 60725 36475 60865
rect 36521 60725 36554 60865
rect 33484 60589 35082 60597
rect 35294 60591 36266 60631
rect 36438 60625 36554 60725
rect 36640 60865 36773 60888
rect 36640 60816 36697 60865
rect 36640 60764 36678 60816
rect 36640 60725 36697 60764
rect 36743 60725 36773 60865
rect 38658 60867 38726 60878
rect 36924 60857 37685 60863
rect 36923 60856 37685 60857
rect 36923 60823 37931 60856
rect 36923 60815 36961 60823
rect 37013 60815 37172 60823
rect 37224 60815 37384 60823
rect 36841 60769 36854 60815
rect 36900 60771 36961 60815
rect 36900 60769 36971 60771
rect 37017 60769 37088 60815
rect 37134 60771 37172 60815
rect 37134 60769 37206 60771
rect 37252 60769 37324 60815
rect 37370 60771 37384 60815
rect 37436 60815 37595 60823
rect 37436 60771 37442 60815
rect 37370 60769 37442 60771
rect 37488 60771 37595 60815
rect 37647 60815 37931 60823
rect 37647 60771 37909 60815
rect 37488 60769 37909 60771
rect 37955 60769 38026 60815
rect 38072 60769 38143 60815
rect 38189 60769 38261 60815
rect 38307 60769 38379 60815
rect 38425 60769 38497 60815
rect 38543 60769 38556 60815
rect 36923 60737 37931 60769
rect 36924 60730 37685 60737
rect 36640 60705 36773 60725
rect 38658 60727 38669 60867
rect 38715 60727 38726 60867
rect 39014 60815 39323 61301
rect 39492 61387 39608 61839
rect 39923 61806 40085 61937
rect 39923 61754 39994 61806
rect 40046 61754 40085 61806
rect 39923 61714 40085 61754
rect 39737 61618 39865 61631
rect 39737 61591 39866 61618
rect 39737 61574 39775 61591
rect 39827 61574 39866 61591
rect 39727 61528 39740 61574
rect 39827 61539 39862 61574
rect 39786 61528 39862 61539
rect 39908 61528 39985 61574
rect 40031 61528 40108 61574
rect 40154 61528 40167 61574
rect 40246 61563 40362 61961
rect 42229 61822 44509 61863
rect 42229 61770 42312 61822
rect 42364 61770 44509 61822
rect 42229 61730 44509 61770
rect 44341 61686 44509 61730
rect 44341 61640 44358 61686
rect 44498 61640 44509 61686
rect 39737 61499 39866 61528
rect 40246 61517 40281 61563
rect 40327 61517 40362 61563
rect 40246 61480 40362 61517
rect 40718 61591 43524 61632
rect 44341 61629 44509 61640
rect 40718 61539 41935 61591
rect 41987 61539 43524 61591
rect 40718 61498 43524 61539
rect 44605 61574 44721 61961
rect 45400 61931 48379 61972
rect 45400 61917 46731 61931
rect 45400 61871 45464 61917
rect 45604 61879 46731 61917
rect 46783 61879 48379 61931
rect 45604 61871 48379 61879
rect 44901 61815 45241 61856
rect 45400 61838 48379 61871
rect 48557 61925 48596 61977
rect 48648 61925 48687 61977
rect 48557 61902 48687 61925
rect 50044 62011 50516 62057
rect 50562 62011 50703 62057
rect 50749 62011 50890 62057
rect 50936 62011 51076 62057
rect 51122 62011 51263 62057
rect 51309 62011 51657 62057
rect 51797 62047 52105 62087
rect 51797 62022 51835 62047
rect 51887 62022 52015 62047
rect 52067 62022 52105 62047
rect 54085 62081 54223 62127
rect 54269 62087 54540 62127
rect 54269 62081 54440 62087
rect 54085 62041 54440 62081
rect 54486 62041 54540 62087
rect 50044 61974 51657 62011
rect 51789 61976 51802 62022
rect 53776 61976 53789 62022
rect 50044 61917 50160 61974
rect 44901 61798 44939 61815
rect 44991 61798 45151 61815
rect 45203 61798 45241 61815
rect 44799 61752 44812 61798
rect 44858 61752 44925 61798
rect 44991 61763 45038 61798
rect 44971 61752 45038 61763
rect 45084 61752 45151 61798
rect 45203 61763 45264 61798
rect 45197 61752 45264 61763
rect 45310 61752 45323 61798
rect 48557 61762 48622 61902
rect 48668 61762 48687 61902
rect 49820 61885 50160 61917
rect 48765 61839 48778 61885
rect 48824 61839 48881 61885
rect 48927 61839 48984 61885
rect 49030 61839 49087 61885
rect 49133 61839 49190 61885
rect 49236 61839 49293 61885
rect 49339 61839 49396 61885
rect 49442 61839 49499 61885
rect 49545 61839 49602 61885
rect 49852 61839 50160 61885
rect 51589 61922 51657 61974
rect 51797 61954 52105 61976
rect 49820 61798 50160 61839
rect 50262 61815 50812 61856
rect 48557 61759 48687 61762
rect 44901 61723 45241 61752
rect 48557 61707 48596 61759
rect 48648 61707 48687 61759
rect 50262 61763 50300 61815
rect 50352 61798 50511 61815
rect 50563 61798 50722 61815
rect 50352 61763 50467 61798
rect 50563 61763 50571 61798
rect 50262 61752 50467 61763
rect 50513 61752 50571 61763
rect 50617 61752 50674 61798
rect 50720 61763 50722 61798
rect 50774 61798 50812 61815
rect 50774 61763 50777 61798
rect 50720 61752 50777 61763
rect 50823 61752 50880 61798
rect 50926 61752 50983 61798
rect 51029 61752 51086 61798
rect 51132 61752 51189 61798
rect 51235 61752 51292 61798
rect 51338 61752 51395 61798
rect 51441 61752 51454 61798
rect 50262 61723 50812 61752
rect 48557 61666 48687 61707
rect 48905 61661 49877 61692
rect 48765 61615 48778 61661
rect 48824 61615 48881 61661
rect 48927 61652 48984 61661
rect 48927 61615 48943 61652
rect 49030 61615 49087 61661
rect 49133 61652 49190 61661
rect 49133 61615 49154 61652
rect 49236 61615 49293 61661
rect 49339 61652 49396 61661
rect 49339 61615 49365 61652
rect 49442 61615 49499 61661
rect 49545 61652 49602 61661
rect 49545 61615 49576 61652
rect 49852 61615 49877 61661
rect 48905 61600 48943 61615
rect 48995 61600 49154 61615
rect 49206 61600 49365 61615
rect 49417 61600 49576 61615
rect 49628 61600 49787 61615
rect 49839 61600 49877 61615
rect 44605 61528 44812 61574
rect 44858 61528 44925 61574
rect 44971 61528 45038 61574
rect 45084 61528 45151 61574
rect 45197 61528 45264 61574
rect 45310 61528 45323 61574
rect 48905 61560 49877 61600
rect 51035 61577 51343 61617
rect 51035 61574 51073 61577
rect 51125 61574 51253 61577
rect 51305 61574 51343 61577
rect 43362 61491 43524 61498
rect 43362 61445 43373 61491
rect 43513 61445 43524 61491
rect 43362 61434 43524 61445
rect 45584 61514 48546 61550
rect 50454 61528 50467 61574
rect 50513 61528 50571 61574
rect 50617 61528 50674 61574
rect 50720 61528 50777 61574
rect 50823 61528 50880 61574
rect 50926 61528 50983 61574
rect 51029 61528 51073 61574
rect 51132 61528 51189 61574
rect 51235 61528 51253 61574
rect 51338 61528 51395 61574
rect 51441 61528 51454 61574
rect 45584 61468 45619 61514
rect 45665 61468 45777 61514
rect 45823 61468 45935 61514
rect 45981 61468 46093 61514
rect 46139 61468 46251 61514
rect 46297 61468 46409 61514
rect 46455 61468 46568 61514
rect 46614 61468 46726 61514
rect 46772 61468 46884 61514
rect 46930 61468 47042 61514
rect 47088 61468 47200 61514
rect 47246 61468 47358 61514
rect 47404 61468 47516 61514
rect 47562 61468 47675 61514
rect 47721 61468 47833 61514
rect 47879 61468 47991 61514
rect 48037 61468 48149 61514
rect 48195 61468 48307 61514
rect 48353 61468 48465 61514
rect 48511 61468 48546 61514
rect 51035 61525 51073 61528
rect 51125 61525 51253 61528
rect 51305 61525 51343 61528
rect 51035 61484 51343 61525
rect 51589 61500 51600 61922
rect 51646 61500 51657 61922
rect 54085 61923 54540 62041
rect 54085 61877 54440 61923
rect 54486 61877 54540 61923
rect 54085 61849 54540 61877
rect 53585 61798 54540 61849
rect 51789 61752 51802 61798
rect 53776 61760 54540 61798
rect 53776 61752 54440 61760
rect 53585 61730 54440 61752
rect 54085 61714 54440 61730
rect 54486 61714 54540 61760
rect 54085 61638 54540 61714
rect 51797 61584 52105 61624
rect 51797 61574 51835 61584
rect 51887 61574 52015 61584
rect 52067 61574 52105 61584
rect 54085 61592 54223 61638
rect 54269 61597 54540 61638
rect 54269 61592 54440 61597
rect 51789 61528 51802 61574
rect 53776 61528 53789 61574
rect 54085 61551 54440 61592
rect 54486 61551 54540 61597
rect 51589 61489 51657 61500
rect 51797 61491 52105 61528
rect 40215 61387 40523 61394
rect 40788 61387 42986 61401
rect 43753 61387 44514 61394
rect 39492 61364 42986 61387
rect 43704 61364 44514 61387
rect 39492 61353 44514 61364
rect 39492 61350 40253 61353
rect 39492 61304 39740 61350
rect 39786 61304 39862 61350
rect 39908 61304 39985 61350
rect 40031 61304 40108 61350
rect 40154 61304 40253 61350
rect 39492 61301 40253 61304
rect 40305 61301 40433 61353
rect 40485 61350 43790 61353
rect 40485 61304 40836 61350
rect 40882 61304 40994 61350
rect 41040 61304 41152 61350
rect 41198 61304 41310 61350
rect 41356 61304 41469 61350
rect 41515 61304 41627 61350
rect 41673 61304 41785 61350
rect 41831 61304 41943 61350
rect 41989 61304 42101 61350
rect 42147 61304 42259 61350
rect 42305 61304 42418 61350
rect 42464 61304 42576 61350
rect 42622 61304 42734 61350
rect 42780 61304 42892 61350
rect 42938 61304 43739 61350
rect 43785 61304 43790 61350
rect 40485 61301 43790 61304
rect 43842 61350 44001 61353
rect 43842 61304 43906 61350
rect 43952 61304 44001 61350
rect 43842 61301 44001 61304
rect 44053 61350 44213 61353
rect 44265 61350 44424 61353
rect 44053 61304 44071 61350
rect 44117 61304 44213 61350
rect 44282 61304 44424 61350
rect 44053 61301 44213 61304
rect 44265 61301 44424 61304
rect 44476 61301 44514 61353
rect 39492 61290 44514 61301
rect 39492 61267 42986 61290
rect 43704 61267 44514 61290
rect 39492 60815 39608 61267
rect 40215 61260 40523 61267
rect 40788 61253 42986 61267
rect 43753 61260 44514 61267
rect 44796 61387 45346 61394
rect 45584 61387 48546 61468
rect 54085 61474 54540 61551
rect 54085 61428 54223 61474
rect 54269 61434 54540 61474
rect 54269 61428 54440 61434
rect 54085 61394 54440 61428
rect 48800 61387 49982 61394
rect 50308 61387 50859 61394
rect 44796 61353 49982 61387
rect 44796 61350 44834 61353
rect 44886 61350 45045 61353
rect 45097 61350 45256 61353
rect 45308 61350 48838 61353
rect 44796 61304 44812 61350
rect 44886 61304 44925 61350
rect 44971 61304 45038 61350
rect 45097 61304 45151 61350
rect 45197 61304 45256 61350
rect 45310 61304 45619 61350
rect 45665 61304 45777 61350
rect 45823 61304 45935 61350
rect 45981 61304 46093 61350
rect 46139 61304 46251 61350
rect 46297 61304 46409 61350
rect 46455 61304 46568 61350
rect 46614 61304 46726 61350
rect 46772 61304 46884 61350
rect 46930 61304 47042 61350
rect 47088 61304 47200 61350
rect 47246 61304 47358 61350
rect 47404 61304 47516 61350
rect 47562 61304 47675 61350
rect 47721 61304 47833 61350
rect 47879 61304 47991 61350
rect 48037 61304 48149 61350
rect 48195 61304 48307 61350
rect 48353 61304 48465 61350
rect 48511 61304 48838 61350
rect 44796 61301 44834 61304
rect 44886 61301 45045 61304
rect 45097 61301 45256 61304
rect 45308 61301 48838 61304
rect 48890 61301 49048 61353
rect 49100 61301 49259 61353
rect 49311 61301 49471 61353
rect 49523 61301 49682 61353
rect 49734 61301 49892 61353
rect 49944 61301 49982 61353
rect 44796 61267 49982 61301
rect 50307 61353 50859 61387
rect 50307 61301 50346 61353
rect 50398 61350 50557 61353
rect 50609 61350 50768 61353
rect 50820 61350 50859 61353
rect 52278 61388 54440 61394
rect 54486 61388 54540 61434
rect 55927 62087 57736 62201
rect 55927 62044 56267 62087
rect 55927 61998 55961 62044
rect 56007 62041 56267 62044
rect 56313 62041 57736 62087
rect 56007 61998 57736 62041
rect 55927 61923 57736 61998
rect 55927 61881 56267 61923
rect 55927 61835 55961 61881
rect 56007 61877 56267 61881
rect 56313 61877 57736 61923
rect 56007 61835 57736 61877
rect 55927 61760 57736 61835
rect 55927 61717 56267 61760
rect 55927 61671 55961 61717
rect 56007 61714 56267 61717
rect 56313 61714 57736 61760
rect 56007 61671 57736 61714
rect 55927 61597 57736 61671
rect 55927 61554 56267 61597
rect 55927 61508 55961 61554
rect 56007 61551 56267 61554
rect 56313 61551 57736 61597
rect 56007 61508 57736 61551
rect 55927 61434 57736 61508
rect 52278 61353 54540 61388
rect 52278 61350 52316 61353
rect 52368 61350 52527 61353
rect 52579 61350 52738 61353
rect 52790 61350 52948 61353
rect 53000 61350 53159 61353
rect 53211 61350 53371 61353
rect 53423 61350 53582 61353
rect 53634 61350 53792 61353
rect 50398 61304 50467 61350
rect 50513 61304 50557 61350
rect 50617 61304 50674 61350
rect 50720 61304 50768 61350
rect 50823 61304 50880 61350
rect 50926 61304 50983 61350
rect 51029 61304 51086 61350
rect 51132 61304 51189 61350
rect 51235 61304 51292 61350
rect 51338 61304 51395 61350
rect 51441 61304 51454 61350
rect 51789 61304 51802 61350
rect 53776 61304 53792 61350
rect 50398 61301 50557 61304
rect 50609 61301 50768 61304
rect 50820 61301 50859 61304
rect 50307 61267 50859 61301
rect 44796 61260 45346 61267
rect 43362 61209 43524 61220
rect 39737 61126 39866 61155
rect 40246 61137 40362 61174
rect 43362 61163 43373 61209
rect 43513 61163 43524 61209
rect 43362 61156 43524 61163
rect 39727 61080 39740 61126
rect 39786 61115 39862 61126
rect 39827 61080 39862 61115
rect 39908 61080 39985 61126
rect 40031 61080 40108 61126
rect 40154 61080 40167 61126
rect 40246 61091 40281 61137
rect 40327 61091 40362 61137
rect 39737 61063 39775 61080
rect 39827 61063 39866 61080
rect 39737 61036 39866 61063
rect 39737 61023 39865 61036
rect 39923 60900 40085 60940
rect 39923 60848 39994 60900
rect 40046 60848 40085 60900
rect 39008 60769 39021 60815
rect 39067 60769 39144 60815
rect 39190 60769 39267 60815
rect 39313 60769 39326 60815
rect 39492 60769 39641 60815
rect 39687 60769 39730 60815
rect 39014 60737 39323 60769
rect 39492 60737 39608 60769
rect 37853 60625 38161 60630
rect 36438 60591 36953 60625
rect 37439 60591 38161 60625
rect 38658 60605 38726 60727
rect 39923 60717 40085 60848
rect 39809 60714 40085 60717
rect 39809 60706 39994 60714
rect 39809 60660 39844 60706
rect 39890 60662 39994 60706
rect 40046 60693 40085 60714
rect 40246 60693 40362 61091
rect 40718 61115 43524 61156
rect 45584 61186 48546 61267
rect 48800 61260 49982 61267
rect 50308 61260 50859 61267
rect 52278 61301 52316 61304
rect 52368 61301 52527 61304
rect 52579 61301 52738 61304
rect 52790 61301 52948 61304
rect 53000 61301 53159 61304
rect 53211 61301 53371 61304
rect 53423 61301 53582 61304
rect 53634 61301 53792 61304
rect 53844 61301 54003 61353
rect 54055 61301 54214 61353
rect 54266 61301 54540 61353
rect 52278 61266 54540 61301
rect 52278 61260 54440 61266
rect 45584 61140 45619 61186
rect 45665 61140 45777 61186
rect 45823 61140 45935 61186
rect 45981 61140 46093 61186
rect 46139 61140 46251 61186
rect 46297 61140 46409 61186
rect 46455 61140 46568 61186
rect 46614 61140 46726 61186
rect 46772 61140 46884 61186
rect 46930 61140 47042 61186
rect 47088 61140 47200 61186
rect 47246 61140 47358 61186
rect 47404 61140 47516 61186
rect 47562 61140 47675 61186
rect 47721 61140 47833 61186
rect 47879 61140 47991 61186
rect 48037 61140 48149 61186
rect 48195 61140 48307 61186
rect 48353 61140 48465 61186
rect 48511 61140 48546 61186
rect 54085 61226 54440 61260
rect 54085 61180 54223 61226
rect 54269 61220 54440 61226
rect 54486 61220 54540 61266
rect 54758 61353 55840 61394
rect 54758 61350 54855 61353
rect 54758 61304 54793 61350
rect 54839 61304 54855 61350
rect 54758 61301 54855 61304
rect 54907 61350 55066 61353
rect 54907 61304 54956 61350
rect 55002 61304 55066 61350
rect 54907 61301 55066 61304
rect 55118 61350 55278 61353
rect 55330 61350 55489 61353
rect 55164 61304 55278 61350
rect 55330 61304 55439 61350
rect 55485 61304 55489 61350
rect 55118 61301 55278 61304
rect 55330 61301 55489 61304
rect 55541 61350 55840 61353
rect 55541 61304 55599 61350
rect 55645 61304 55760 61350
rect 55806 61304 55840 61350
rect 55541 61301 55840 61304
rect 54758 61261 55840 61301
rect 55927 61388 56267 61434
rect 56313 61388 57736 61434
rect 55927 61266 57736 61388
rect 54817 61260 55579 61261
rect 54269 61180 54540 61220
rect 40718 61063 41935 61115
rect 41987 61063 43524 61115
rect 40718 61022 43524 61063
rect 44605 61080 44812 61126
rect 44858 61080 44925 61126
rect 44971 61080 45038 61126
rect 45084 61080 45151 61126
rect 45197 61080 45264 61126
rect 45310 61080 45323 61126
rect 45584 61104 48546 61140
rect 51035 61129 51343 61170
rect 51035 61126 51073 61129
rect 51125 61126 51253 61129
rect 51305 61126 51343 61129
rect 51589 61154 51657 61165
rect 44341 61014 44509 61025
rect 44341 60968 44358 61014
rect 44498 60968 44509 61014
rect 44341 60924 44509 60968
rect 42229 60884 44509 60924
rect 42229 60832 42312 60884
rect 42364 60832 44509 60884
rect 42229 60791 44509 60832
rect 44605 60693 44721 61080
rect 48905 61054 49877 61094
rect 50454 61080 50467 61126
rect 50513 61080 50571 61126
rect 50617 61080 50674 61126
rect 50720 61080 50777 61126
rect 50823 61080 50880 61126
rect 50926 61080 50983 61126
rect 51029 61080 51073 61126
rect 51132 61080 51189 61126
rect 51235 61080 51253 61126
rect 51338 61080 51395 61126
rect 51441 61080 51454 61126
rect 48905 61039 48943 61054
rect 48995 61039 49154 61054
rect 49206 61039 49365 61054
rect 49417 61039 49576 61054
rect 49628 61039 49787 61054
rect 49839 61039 49877 61054
rect 48765 60993 48778 61039
rect 48824 60993 48881 61039
rect 48927 61002 48943 61039
rect 48927 60993 48984 61002
rect 49030 60993 49087 61039
rect 49133 61002 49154 61039
rect 49133 60993 49190 61002
rect 49236 60993 49293 61039
rect 49339 61002 49365 61039
rect 49339 60993 49396 61002
rect 49442 60993 49499 61039
rect 49545 61002 49576 61039
rect 49545 60993 49602 61002
rect 49852 60993 49877 61039
rect 51035 61077 51073 61080
rect 51125 61077 51253 61080
rect 51305 61077 51343 61080
rect 51035 61037 51343 61077
rect 48557 60947 48687 60988
rect 48905 60962 49877 60993
rect 44901 60902 45241 60931
rect 44799 60856 44812 60902
rect 44858 60856 44925 60902
rect 44971 60891 45038 60902
rect 44991 60856 45038 60891
rect 45084 60856 45151 60902
rect 45197 60891 45264 60902
rect 45203 60856 45264 60891
rect 45310 60856 45323 60902
rect 48557 60895 48596 60947
rect 48648 60895 48687 60947
rect 48557 60892 48687 60895
rect 44901 60839 44939 60856
rect 44991 60839 45151 60856
rect 45203 60839 45241 60856
rect 44901 60798 45241 60839
rect 45400 60783 48379 60816
rect 45400 60737 45464 60783
rect 45604 60775 48379 60783
rect 45604 60737 47108 60775
rect 45400 60723 47108 60737
rect 47160 60723 48379 60775
rect 40046 60678 44918 60693
rect 45400 60682 48379 60723
rect 48557 60752 48622 60892
rect 48668 60752 48687 60892
rect 50262 60902 50812 60931
rect 50262 60891 50467 60902
rect 50513 60891 50571 60902
rect 49820 60815 50160 60856
rect 48765 60769 48778 60815
rect 48824 60769 48881 60815
rect 48927 60769 48984 60815
rect 49030 60769 49087 60815
rect 49133 60769 49190 60815
rect 49236 60769 49293 60815
rect 49339 60769 49396 60815
rect 49442 60769 49499 60815
rect 49545 60769 49602 60815
rect 49852 60769 50160 60815
rect 50262 60839 50300 60891
rect 50352 60856 50467 60891
rect 50563 60856 50571 60891
rect 50617 60856 50674 60902
rect 50720 60891 50777 60902
rect 50720 60856 50722 60891
rect 50352 60839 50511 60856
rect 50563 60839 50722 60856
rect 50774 60856 50777 60891
rect 50823 60856 50880 60902
rect 50926 60856 50983 60902
rect 51029 60856 51086 60902
rect 51132 60856 51189 60902
rect 51235 60856 51292 60902
rect 51338 60856 51395 60902
rect 51441 60856 51454 60902
rect 50774 60839 50812 60856
rect 50262 60798 50812 60839
rect 48557 60729 48687 60752
rect 49820 60737 50160 60769
rect 40046 60662 44812 60678
rect 39890 60660 44812 60662
rect 39809 60657 44812 60660
rect 39809 60611 43739 60657
rect 43785 60611 43906 60657
rect 43952 60611 44071 60657
rect 44117 60611 44236 60657
rect 44282 60632 44812 60657
rect 44858 60632 44925 60678
rect 44971 60632 45038 60678
rect 45084 60632 45151 60678
rect 45197 60632 45264 60678
rect 45310 60632 45323 60678
rect 48557 60677 48596 60729
rect 48648 60677 48687 60729
rect 48557 60637 48687 60677
rect 50044 60680 50160 60737
rect 51589 60732 51600 61154
rect 51646 60732 51657 61154
rect 51797 61126 52105 61163
rect 51789 61080 51802 61126
rect 53776 61080 53789 61126
rect 54085 61103 54540 61180
rect 51797 61070 51835 61080
rect 51887 61070 52015 61080
rect 52067 61070 52105 61080
rect 51797 61030 52105 61070
rect 54085 61062 54440 61103
rect 54085 61016 54223 61062
rect 54269 61057 54440 61062
rect 54486 61057 54540 61103
rect 54269 61016 54540 61057
rect 54085 60940 54540 61016
rect 54085 60924 54440 60940
rect 53585 60902 54440 60924
rect 51789 60856 51802 60902
rect 53776 60894 54440 60902
rect 54486 60894 54540 60940
rect 53776 60856 54540 60894
rect 53585 60805 54540 60856
rect 51589 60680 51657 60732
rect 54085 60777 54540 60805
rect 54085 60731 54440 60777
rect 54486 60731 54540 60777
rect 50044 60643 51657 60680
rect 51797 60678 52105 60700
rect 44282 60611 44918 60632
rect 38658 60591 39723 60605
rect 30683 60567 30855 60573
rect 30583 60527 30855 60567
rect 30901 60527 31040 60573
rect 33484 60560 34643 60589
rect 35260 60545 35273 60591
rect 35523 60545 35543 60591
rect 35626 60545 35683 60591
rect 35729 60545 35754 60591
rect 35832 60545 35889 60591
rect 35935 60545 35965 60591
rect 36038 60545 36095 60591
rect 36141 60545 36176 60591
rect 36244 60545 36301 60591
rect 36347 60545 36360 60591
rect 36438 60545 36854 60591
rect 36900 60545 36971 60591
rect 37017 60545 37088 60591
rect 37134 60545 37206 60591
rect 37252 60545 37324 60591
rect 37370 60545 37442 60591
rect 37488 60589 37909 60591
rect 37488 60545 37891 60589
rect 37955 60545 38026 60591
rect 38072 60589 38143 60591
rect 38123 60545 38143 60589
rect 38189 60545 38261 60591
rect 38307 60545 38379 60591
rect 38425 60545 38497 60591
rect 38543 60545 38556 60591
rect 38658 60545 39021 60591
rect 39067 60545 39144 60591
rect 39190 60545 39267 60591
rect 39313 60545 39641 60591
rect 39687 60545 39730 60591
rect 39809 60573 44918 60611
rect 48905 60591 49877 60631
rect 48765 60545 48778 60591
rect 48824 60545 48881 60591
rect 48927 60545 48943 60591
rect 49030 60545 49087 60591
rect 49133 60545 49154 60591
rect 49236 60545 49293 60591
rect 49339 60545 49365 60591
rect 49442 60545 49499 60591
rect 49545 60545 49576 60591
rect 49852 60545 49877 60591
rect 50044 60597 50516 60643
rect 50562 60597 50703 60643
rect 50749 60597 50890 60643
rect 50936 60597 51076 60643
rect 51122 60597 51263 60643
rect 51309 60597 51657 60643
rect 51789 60632 51802 60678
rect 53776 60632 53789 60678
rect 50044 60587 51657 60597
rect 50481 60560 51657 60587
rect 51797 60607 51835 60632
rect 51887 60607 52015 60632
rect 52067 60607 52105 60632
rect 51797 60567 52105 60607
rect 54085 60613 54540 60731
rect 54085 60573 54440 60613
rect 30583 60494 31040 60527
rect 35294 60539 35332 60545
rect 35384 60539 35543 60545
rect 35595 60539 35754 60545
rect 35806 60539 35965 60545
rect 36017 60539 36176 60545
rect 36228 60539 36266 60545
rect 34870 60494 35025 60501
rect 35294 60499 36266 60539
rect 36438 60505 36953 60545
rect 37439 60537 37891 60545
rect 37943 60537 38071 60545
rect 38123 60537 38161 60545
rect 37439 60505 38161 60537
rect 37853 60497 38161 60505
rect 27387 60401 27790 60453
rect 27842 60401 28001 60453
rect 28053 60401 28212 60453
rect 28264 60401 28423 60453
rect 28475 60401 28634 60453
rect 28686 60450 28845 60453
rect 28686 60404 28810 60450
rect 28686 60401 28845 60404
rect 28897 60401 29056 60453
rect 29108 60401 29196 60453
rect 27387 60287 29196 60401
rect 29283 60453 30365 60494
rect 29283 60450 29582 60453
rect 29283 60404 29317 60450
rect 29363 60404 29478 60450
rect 29524 60404 29582 60450
rect 29283 60401 29582 60404
rect 29634 60450 29793 60453
rect 29845 60450 30005 60453
rect 29634 60404 29638 60450
rect 29684 60404 29793 60450
rect 29845 60404 29959 60450
rect 29634 60401 29793 60404
rect 29845 60401 30005 60404
rect 30057 60450 30216 60453
rect 30057 60404 30121 60450
rect 30167 60404 30216 60450
rect 30057 60401 30216 60404
rect 30268 60450 30365 60453
rect 30268 60404 30284 60450
rect 30330 60404 30365 60450
rect 30268 60401 30365 60404
rect 29283 60361 30365 60401
rect 30583 60453 32842 60494
rect 30583 60450 30854 60453
rect 30583 60404 30637 60450
rect 30683 60404 30854 60450
rect 30583 60401 30854 60404
rect 30906 60401 31065 60453
rect 31117 60401 31276 60453
rect 31328 60401 31486 60453
rect 31538 60401 31697 60453
rect 31749 60401 31909 60453
rect 31961 60401 32120 60453
rect 32172 60401 32330 60453
rect 32382 60401 32541 60453
rect 32593 60401 32752 60453
rect 32804 60401 32842 60453
rect 29544 60360 30306 60361
rect 30583 60360 32842 60401
rect 34717 60453 35025 60494
rect 38658 60485 39723 60545
rect 48905 60539 48943 60545
rect 48995 60539 49154 60545
rect 49206 60539 49365 60545
rect 49417 60539 49576 60545
rect 49628 60539 49787 60545
rect 49839 60539 49877 60545
rect 48905 60499 49877 60539
rect 54085 60527 54223 60573
rect 54269 60567 54440 60573
rect 54486 60567 54540 60613
rect 54269 60527 54540 60567
rect 50099 60494 50255 60501
rect 54085 60494 54540 60527
rect 55927 61220 56267 61266
rect 56313 61220 57736 61266
rect 55927 61144 57736 61220
rect 55927 61098 55961 61144
rect 56007 61103 57736 61144
rect 56007 61098 56267 61103
rect 55927 61057 56267 61098
rect 56313 61057 57736 61103
rect 55927 60981 57736 61057
rect 55927 60935 55961 60981
rect 56007 60940 57736 60981
rect 56007 60935 56267 60940
rect 55927 60894 56267 60935
rect 56313 60894 57736 60940
rect 55927 60817 57736 60894
rect 55927 60771 55961 60817
rect 56007 60777 57736 60817
rect 56007 60771 56267 60777
rect 55927 60731 56267 60771
rect 56313 60731 57736 60777
rect 55927 60654 57736 60731
rect 55927 60608 55961 60654
rect 56007 60613 57736 60654
rect 56007 60608 56267 60613
rect 55927 60567 56267 60608
rect 56313 60567 57736 60613
rect 34717 60401 34755 60453
rect 34807 60450 34935 60453
rect 34807 60404 34916 60450
rect 34807 60401 34935 60404
rect 34987 60401 35025 60453
rect 34717 60360 35025 60401
rect 50099 60453 50408 60494
rect 50099 60401 50138 60453
rect 50190 60450 50318 60453
rect 50206 60404 50318 60450
rect 50190 60401 50318 60404
rect 50370 60401 50408 60453
rect 27387 60241 28810 60287
rect 28856 60244 29196 60287
rect 28856 60241 29116 60244
rect 27387 60198 29116 60241
rect 29162 60198 29196 60244
rect 27387 60123 29196 60198
rect 27387 60077 28810 60123
rect 28856 60081 29196 60123
rect 28856 60077 29116 60081
rect 27387 60035 29116 60077
rect 29162 60035 29196 60081
rect 27387 59960 29196 60035
rect 27387 59914 28810 59960
rect 28856 59917 29196 59960
rect 28856 59914 29116 59917
rect 27387 59871 29116 59914
rect 29162 59871 29196 59917
rect 27387 59797 29196 59871
rect 27387 59751 28810 59797
rect 28856 59754 29196 59797
rect 28856 59751 29116 59754
rect 27387 59708 29116 59751
rect 29162 59708 29196 59754
rect 27387 59634 29196 59708
rect 27387 59588 28810 59634
rect 28856 59588 29196 59634
rect 30583 60327 31040 60360
rect 34870 60353 35025 60360
rect 30583 60287 30855 60327
rect 30583 60241 30637 60287
rect 30683 60281 30855 60287
rect 30901 60281 31040 60327
rect 35294 60315 36266 60355
rect 37853 60349 38161 60357
rect 35294 60309 35332 60315
rect 35384 60309 35543 60315
rect 35595 60309 35754 60315
rect 35806 60309 35965 60315
rect 36017 60309 36176 60315
rect 36228 60309 36266 60315
rect 36438 60309 36953 60349
rect 37439 60317 38161 60349
rect 37439 60309 37891 60317
rect 37943 60309 38071 60317
rect 38123 60309 38161 60317
rect 38658 60309 39723 60369
rect 50099 60360 50408 60401
rect 52278 60453 54540 60494
rect 52278 60401 52316 60453
rect 52368 60401 52527 60453
rect 52579 60401 52738 60453
rect 52790 60401 52948 60453
rect 53000 60401 53159 60453
rect 53211 60401 53371 60453
rect 53423 60401 53582 60453
rect 53634 60401 53792 60453
rect 53844 60401 54003 60453
rect 54055 60401 54214 60453
rect 54266 60450 54540 60453
rect 54266 60404 54440 60450
rect 54486 60404 54540 60450
rect 54266 60401 54540 60404
rect 52278 60360 54540 60401
rect 54758 60453 55840 60494
rect 54758 60450 54855 60453
rect 54758 60404 54793 60450
rect 54839 60404 54855 60450
rect 54758 60401 54855 60404
rect 54907 60450 55066 60453
rect 54907 60404 54956 60450
rect 55002 60404 55066 60450
rect 54907 60401 55066 60404
rect 55118 60450 55278 60453
rect 55330 60450 55489 60453
rect 55164 60404 55278 60450
rect 55330 60404 55439 60450
rect 55485 60404 55489 60450
rect 55118 60401 55278 60404
rect 55330 60401 55489 60404
rect 55541 60450 55840 60453
rect 55541 60404 55599 60450
rect 55645 60404 55760 60450
rect 55806 60404 55840 60450
rect 55541 60401 55840 60404
rect 54758 60361 55840 60401
rect 55927 60453 57736 60567
rect 55927 60401 56015 60453
rect 56067 60401 56226 60453
rect 56278 60450 56437 60453
rect 56313 60404 56437 60450
rect 56278 60401 56437 60404
rect 56489 60401 56648 60453
rect 56700 60401 56859 60453
rect 56911 60401 57070 60453
rect 57122 60401 57281 60453
rect 57333 60401 57736 60453
rect 54817 60360 55579 60361
rect 48905 60315 49877 60355
rect 50099 60353 50255 60360
rect 48905 60309 48943 60315
rect 48995 60309 49154 60315
rect 49206 60309 49365 60315
rect 49417 60309 49576 60315
rect 49628 60309 49787 60315
rect 49839 60309 49877 60315
rect 30683 60241 31040 60281
rect 33484 60265 34643 60294
rect 30583 60164 31040 60241
rect 33019 60225 33327 60265
rect 33019 60222 33057 60225
rect 33109 60222 33237 60225
rect 33289 60222 33327 60225
rect 33484 60257 35082 60265
rect 35260 60263 35273 60309
rect 35523 60263 35543 60309
rect 35626 60263 35683 60309
rect 35729 60263 35754 60309
rect 35832 60263 35889 60309
rect 35935 60263 35965 60309
rect 36038 60263 36095 60309
rect 36141 60263 36176 60309
rect 36244 60263 36301 60309
rect 36347 60263 36360 60309
rect 36438 60263 36854 60309
rect 36900 60263 36971 60309
rect 37017 60263 37088 60309
rect 37134 60263 37206 60309
rect 37252 60263 37324 60309
rect 37370 60263 37442 60309
rect 37488 60265 37891 60309
rect 37488 60263 37909 60265
rect 37955 60263 38026 60309
rect 38123 60265 38143 60309
rect 38072 60263 38143 60265
rect 38189 60263 38261 60309
rect 38307 60263 38379 60309
rect 38425 60263 38497 60309
rect 38543 60263 38556 60309
rect 38658 60263 39021 60309
rect 39067 60263 39144 60309
rect 39190 60263 39267 60309
rect 39313 60263 39641 60309
rect 39687 60263 39730 60309
rect 31336 60176 31349 60222
rect 33323 60176 33336 60222
rect 33484 60211 33816 60257
rect 33862 60211 34002 60257
rect 34048 60211 34189 60257
rect 34235 60211 34376 60257
rect 34422 60211 34562 60257
rect 34608 60211 35082 60257
rect 35294 60223 36266 60263
rect 36438 60229 36953 60263
rect 37439 60229 38161 60263
rect 30583 60123 30855 60164
rect 30583 60077 30637 60123
rect 30683 60118 30855 60123
rect 30901 60118 31040 60164
rect 33019 60173 33057 60176
rect 33109 60173 33237 60176
rect 33289 60173 33327 60176
rect 33019 60132 33327 60173
rect 33484 60174 35082 60211
rect 30683 60077 31040 60118
rect 30583 60049 31040 60077
rect 33484 60092 33552 60174
rect 30583 60001 31493 60049
rect 30583 59960 30855 60001
rect 30583 59914 30637 59960
rect 30683 59955 30855 59960
rect 30901 59998 31493 60001
rect 30901 59955 31349 59998
rect 30683 59952 31349 59955
rect 33323 59952 33336 59998
rect 30683 59930 31493 59952
rect 30683 59914 31040 59930
rect 30583 59838 31040 59914
rect 30583 59797 30855 59838
rect 30583 59751 30637 59797
rect 30683 59792 30855 59797
rect 30901 59792 31040 59838
rect 30683 59751 31040 59792
rect 33019 59777 33327 59817
rect 33019 59774 33057 59777
rect 33109 59774 33237 59777
rect 33289 59774 33327 59777
rect 30583 59674 31040 59751
rect 31336 59728 31349 59774
rect 33323 59728 33336 59774
rect 33019 59725 33057 59728
rect 33109 59725 33237 59728
rect 33289 59725 33327 59728
rect 33019 59684 33327 59725
rect 30583 59634 30855 59674
rect 27387 59466 29196 59588
rect 27387 59420 28810 59466
rect 28856 59420 29196 59466
rect 29283 59553 30365 59594
rect 29283 59550 29582 59553
rect 29283 59504 29317 59550
rect 29363 59504 29478 59550
rect 29524 59504 29582 59550
rect 29283 59501 29582 59504
rect 29634 59550 29793 59553
rect 29845 59550 30005 59553
rect 29634 59504 29638 59550
rect 29684 59504 29793 59550
rect 29845 59504 29959 59550
rect 29634 59501 29793 59504
rect 29845 59501 30005 59504
rect 30057 59550 30216 59553
rect 30057 59504 30121 59550
rect 30167 59504 30216 59550
rect 30057 59501 30216 59504
rect 30268 59550 30365 59553
rect 30268 59504 30284 59550
rect 30330 59504 30365 59550
rect 30268 59501 30365 59504
rect 29283 59461 30365 59501
rect 30583 59588 30637 59634
rect 30683 59628 30855 59634
rect 30901 59628 31040 59674
rect 33484 59670 33495 60092
rect 33541 59670 33552 60092
rect 34964 60117 35082 60174
rect 36438 60129 36554 60229
rect 37853 60224 38161 60229
rect 38658 60249 39723 60263
rect 34964 60085 36360 60117
rect 34228 60015 34718 60056
rect 34228 59998 34267 60015
rect 34319 59998 34447 60015
rect 34499 59998 34627 60015
rect 33671 59952 33684 59998
rect 33730 59952 33787 59998
rect 33833 59952 33890 59998
rect 33936 59952 33993 59998
rect 34039 59952 34096 59998
rect 34142 59952 34199 59998
rect 34245 59963 34267 59998
rect 34245 59952 34302 59963
rect 34348 59952 34405 59998
rect 34499 59963 34508 59998
rect 34451 59952 34508 59963
rect 34554 59952 34612 59998
rect 34679 59963 34718 60015
rect 34964 60039 35273 60085
rect 35523 60039 35580 60085
rect 35626 60039 35683 60085
rect 35729 60039 35786 60085
rect 35832 60039 35889 60085
rect 35935 60039 35992 60085
rect 36038 60039 36095 60085
rect 36141 60039 36198 60085
rect 36244 60039 36301 60085
rect 36347 60039 36360 60085
rect 34964 59995 36360 60039
rect 34658 59952 34718 59963
rect 34228 59923 34718 59952
rect 36438 59989 36475 60129
rect 36521 59989 36554 60129
rect 35294 59861 36266 59895
rect 36438 59886 36554 59989
rect 36640 60129 36773 60149
rect 36640 60090 36697 60129
rect 36640 60038 36678 60090
rect 36640 59989 36697 60038
rect 36743 59989 36773 60129
rect 38658 60127 38726 60249
rect 39809 60243 44918 60281
rect 48765 60263 48778 60309
rect 48824 60263 48881 60309
rect 48927 60263 48943 60309
rect 49030 60263 49087 60309
rect 49133 60263 49154 60309
rect 49236 60263 49293 60309
rect 49339 60263 49365 60309
rect 49442 60263 49499 60309
rect 49545 60263 49576 60309
rect 49852 60263 49877 60309
rect 54085 60327 54540 60360
rect 50481 60267 51657 60294
rect 39809 60197 43739 60243
rect 43785 60197 43906 60243
rect 43952 60197 44071 60243
rect 44117 60197 44236 60243
rect 44282 60222 44918 60243
rect 48905 60223 49877 60263
rect 50044 60257 51657 60267
rect 44282 60197 44812 60222
rect 39809 60194 44812 60197
rect 39809 60148 39844 60194
rect 39890 60192 44812 60194
rect 39890 60148 39994 60192
rect 39809 60140 39994 60148
rect 40046 60176 44812 60192
rect 44858 60176 44925 60222
rect 44971 60176 45038 60222
rect 45084 60176 45151 60222
rect 45197 60176 45264 60222
rect 45310 60176 45323 60222
rect 48557 60177 48687 60217
rect 40046 60161 44918 60176
rect 40046 60140 40085 60161
rect 39809 60137 40085 60140
rect 36924 60117 37685 60124
rect 36923 60085 37931 60117
rect 36841 60039 36854 60085
rect 36900 60083 36971 60085
rect 36900 60039 36961 60083
rect 37017 60039 37088 60085
rect 37134 60083 37206 60085
rect 37134 60039 37172 60083
rect 37252 60039 37324 60085
rect 37370 60083 37442 60085
rect 37370 60039 37384 60083
rect 36923 60031 36961 60039
rect 37013 60031 37172 60039
rect 37224 60031 37384 60039
rect 37436 60039 37442 60083
rect 37488 60083 37909 60085
rect 37488 60039 37595 60083
rect 37436 60031 37595 60039
rect 37647 60039 37909 60083
rect 37955 60039 38026 60085
rect 38072 60039 38143 60085
rect 38189 60039 38261 60085
rect 38307 60039 38379 60085
rect 38425 60039 38497 60085
rect 38543 60039 38556 60085
rect 37647 60031 37931 60039
rect 36923 59998 37931 60031
rect 36923 59997 37685 59998
rect 36924 59991 37685 59997
rect 36640 59966 36773 59989
rect 38658 59987 38669 60127
rect 38715 59987 38726 60127
rect 39014 60085 39323 60117
rect 39492 60085 39608 60117
rect 39008 60039 39021 60085
rect 39067 60039 39144 60085
rect 39190 60039 39267 60085
rect 39313 60039 39326 60085
rect 39492 60039 39641 60085
rect 39687 60039 39730 60085
rect 38658 59976 38726 59987
rect 36438 59861 36953 59886
rect 37439 59883 37931 59886
rect 37439 59861 38161 59883
rect 35260 59815 35273 59861
rect 35523 59855 35580 59861
rect 35523 59815 35543 59855
rect 35626 59815 35683 59861
rect 35729 59855 35786 59861
rect 35729 59815 35754 59855
rect 35832 59815 35889 59861
rect 35935 59855 35992 59861
rect 35935 59815 35965 59855
rect 36038 59815 36095 59861
rect 36141 59855 36198 59861
rect 36141 59815 36176 59855
rect 36244 59815 36301 59861
rect 36347 59815 36360 59861
rect 36438 59815 36854 59861
rect 36900 59815 36971 59861
rect 37017 59815 37088 59861
rect 37134 59815 37206 59861
rect 37252 59815 37324 59861
rect 37370 59815 37442 59861
rect 37488 59843 37909 59861
rect 37488 59815 37891 59843
rect 37955 59815 38026 59861
rect 38072 59843 38143 59861
rect 38123 59815 38143 59843
rect 38189 59815 38261 59861
rect 38307 59815 38379 59861
rect 38425 59815 38497 59861
rect 38543 59815 38556 59861
rect 33781 59774 34089 59809
rect 35294 59803 35332 59815
rect 35384 59803 35543 59815
rect 35595 59803 35754 59815
rect 35806 59803 35965 59815
rect 36017 59803 36176 59815
rect 36228 59803 36266 59815
rect 33671 59728 33684 59774
rect 33730 59728 33787 59774
rect 33833 59769 33890 59774
rect 33871 59728 33890 59769
rect 33936 59728 33993 59774
rect 34039 59769 34096 59774
rect 34051 59728 34096 59769
rect 34142 59728 34199 59774
rect 34245 59728 34302 59774
rect 34348 59728 34405 59774
rect 34451 59728 34508 59774
rect 34554 59728 34612 59774
rect 34658 59728 34671 59774
rect 35294 59763 36266 59803
rect 36438 59766 36953 59815
rect 37439 59791 37891 59815
rect 37943 59791 38071 59815
rect 38123 59791 38161 59815
rect 37439 59766 38161 59791
rect 37853 59750 38161 59766
rect 33781 59717 33819 59728
rect 33871 59717 33999 59728
rect 34051 59717 34089 59728
rect 33781 59676 34089 59717
rect 33484 59659 33552 59670
rect 30683 59594 31040 59628
rect 30683 59588 32842 59594
rect 30583 59553 32842 59588
rect 34247 59587 35008 59594
rect 30583 59501 30854 59553
rect 30906 59501 31065 59553
rect 31117 59501 31276 59553
rect 31328 59550 31486 59553
rect 31538 59550 31697 59553
rect 31749 59550 31909 59553
rect 31961 59550 32120 59553
rect 32172 59550 32330 59553
rect 32382 59550 32541 59553
rect 32593 59550 32752 59553
rect 32804 59550 32842 59553
rect 34246 59553 35008 59587
rect 34246 59550 34284 59553
rect 34336 59550 34495 59553
rect 34547 59550 34707 59553
rect 31328 59504 31349 59550
rect 33323 59504 33336 59550
rect 33671 59504 33684 59550
rect 33730 59504 33787 59550
rect 33833 59504 33890 59550
rect 33936 59504 33993 59550
rect 34039 59504 34096 59550
rect 34142 59504 34199 59550
rect 34245 59504 34284 59550
rect 34348 59504 34405 59550
rect 34451 59504 34495 59550
rect 34554 59504 34612 59550
rect 34658 59504 34707 59550
rect 31328 59501 31486 59504
rect 31538 59501 31697 59504
rect 31749 59501 31909 59504
rect 31961 59501 32120 59504
rect 32172 59501 32330 59504
rect 32382 59501 32541 59504
rect 32593 59501 32752 59504
rect 32804 59501 32842 59504
rect 30583 59466 32842 59501
rect 34246 59501 34284 59504
rect 34336 59501 34495 59504
rect 34547 59501 34707 59504
rect 34759 59501 34918 59553
rect 34970 59501 35008 59553
rect 34246 59467 35008 59501
rect 29544 59460 30306 59461
rect 27387 59344 29196 59420
rect 27387 59303 29116 59344
rect 27387 59257 28810 59303
rect 28856 59298 29116 59303
rect 29162 59298 29196 59344
rect 28856 59257 29196 59298
rect 27387 59181 29196 59257
rect 27387 59140 29116 59181
rect 27387 59094 28810 59140
rect 28856 59135 29116 59140
rect 29162 59135 29196 59181
rect 28856 59094 29196 59135
rect 27387 59017 29196 59094
rect 27387 58977 29116 59017
rect 27387 58931 28810 58977
rect 28856 58971 29116 58977
rect 29162 58971 29196 59017
rect 28856 58931 29196 58971
rect 27387 58854 29196 58931
rect 27387 58813 29116 58854
rect 27387 58767 28810 58813
rect 28856 58808 29116 58813
rect 29162 58808 29196 58854
rect 28856 58767 29196 58808
rect 27387 58653 29196 58767
rect 30583 59420 30637 59466
rect 30683 59460 32842 59466
rect 34247 59460 35008 59467
rect 35182 59587 36364 59594
rect 35182 59553 36958 59587
rect 35182 59501 35220 59553
rect 35272 59501 35430 59553
rect 35482 59501 35641 59553
rect 35693 59501 35853 59553
rect 35905 59501 36064 59553
rect 36116 59501 36274 59553
rect 36326 59550 36958 59553
rect 36326 59504 36489 59550
rect 36723 59504 36958 59550
rect 36326 59501 36958 59504
rect 35182 59467 36958 59501
rect 37946 59553 38842 59594
rect 37946 59550 38330 59553
rect 38382 59550 38541 59553
rect 37946 59504 37957 59550
rect 38473 59504 38541 59550
rect 37946 59501 38330 59504
rect 38382 59501 38541 59504
rect 38593 59501 38752 59553
rect 38804 59501 38842 59553
rect 35182 59460 36364 59467
rect 37946 59460 38842 59501
rect 39014 59553 39323 60039
rect 39014 59501 39052 59553
rect 39104 59550 39232 59553
rect 39108 59504 39220 59550
rect 39104 59501 39232 59504
rect 39284 59501 39323 59553
rect 30683 59426 31040 59460
rect 30683 59420 30855 59426
rect 30583 59380 30855 59420
rect 30901 59380 31040 59426
rect 30583 59303 31040 59380
rect 33484 59384 33552 59395
rect 33019 59329 33327 59370
rect 33019 59326 33057 59329
rect 33109 59326 33237 59329
rect 33289 59326 33327 59329
rect 30583 59257 30637 59303
rect 30683 59262 31040 59303
rect 31336 59280 31349 59326
rect 33323 59280 33336 59326
rect 30683 59257 30855 59262
rect 30583 59216 30855 59257
rect 30901 59216 31040 59262
rect 33019 59277 33057 59280
rect 33109 59277 33237 59280
rect 33289 59277 33327 59280
rect 33019 59237 33327 59277
rect 30583 59140 31040 59216
rect 30583 59094 30637 59140
rect 30683 59124 31040 59140
rect 30683 59102 31493 59124
rect 30683 59099 31349 59102
rect 30683 59094 30855 59099
rect 30583 59053 30855 59094
rect 30901 59056 31349 59099
rect 33323 59056 33336 59102
rect 30901 59053 31493 59056
rect 30583 59005 31493 59053
rect 30583 58977 31040 59005
rect 30583 58931 30637 58977
rect 30683 58936 31040 58977
rect 30683 58931 30855 58936
rect 30583 58890 30855 58931
rect 30901 58890 31040 58936
rect 33484 58962 33495 59384
rect 33541 58962 33552 59384
rect 33781 59337 34089 59378
rect 33781 59326 33819 59337
rect 33871 59326 33999 59337
rect 34051 59326 34089 59337
rect 33671 59280 33684 59326
rect 33730 59280 33787 59326
rect 33871 59285 33890 59326
rect 33833 59280 33890 59285
rect 33936 59280 33993 59326
rect 34051 59285 34096 59326
rect 34039 59280 34096 59285
rect 34142 59280 34199 59326
rect 34245 59280 34302 59326
rect 34348 59280 34405 59326
rect 34451 59280 34508 59326
rect 34554 59280 34612 59326
rect 34658 59280 34671 59326
rect 33781 59245 34089 59280
rect 35294 59251 36266 59291
rect 37853 59288 38161 59304
rect 35294 59239 35332 59251
rect 35384 59239 35543 59251
rect 35595 59239 35754 59251
rect 35806 59239 35965 59251
rect 36017 59239 36176 59251
rect 36228 59239 36266 59251
rect 36438 59239 36953 59288
rect 37439 59263 38161 59288
rect 37439 59239 37891 59263
rect 37943 59239 38071 59263
rect 38123 59239 38161 59263
rect 35260 59193 35273 59239
rect 35523 59199 35543 59239
rect 35523 59193 35580 59199
rect 35626 59193 35683 59239
rect 35729 59199 35754 59239
rect 35729 59193 35786 59199
rect 35832 59193 35889 59239
rect 35935 59199 35965 59239
rect 35935 59193 35992 59199
rect 36038 59193 36095 59239
rect 36141 59199 36176 59239
rect 36141 59193 36198 59199
rect 36244 59193 36301 59239
rect 36347 59193 36360 59239
rect 36438 59193 36854 59239
rect 36900 59193 36971 59239
rect 37017 59193 37088 59239
rect 37134 59193 37206 59239
rect 37252 59193 37324 59239
rect 37370 59193 37442 59239
rect 37488 59211 37891 59239
rect 37488 59193 37909 59211
rect 37955 59193 38026 59239
rect 38123 59211 38143 59239
rect 38072 59193 38143 59211
rect 38189 59193 38261 59239
rect 38307 59193 38379 59239
rect 38425 59193 38497 59239
rect 38543 59193 38556 59239
rect 35294 59159 36266 59193
rect 36438 59168 36953 59193
rect 37439 59171 38161 59193
rect 37439 59168 37931 59171
rect 34228 59102 34718 59131
rect 33671 59056 33684 59102
rect 33730 59056 33787 59102
rect 33833 59056 33890 59102
rect 33936 59056 33993 59102
rect 34039 59056 34096 59102
rect 34142 59056 34199 59102
rect 34245 59091 34302 59102
rect 34245 59056 34267 59091
rect 34348 59056 34405 59102
rect 34451 59091 34508 59102
rect 34499 59056 34508 59091
rect 34554 59056 34612 59102
rect 34658 59091 34718 59102
rect 34228 59039 34267 59056
rect 34319 59039 34447 59056
rect 34499 59039 34627 59056
rect 34679 59039 34718 59091
rect 36438 59065 36554 59168
rect 34228 58998 34718 59039
rect 34964 59015 36360 59059
rect 30583 58813 31040 58890
rect 33019 58881 33327 58922
rect 33019 58878 33057 58881
rect 33109 58878 33237 58881
rect 33289 58878 33327 58881
rect 33484 58880 33552 58962
rect 34964 58969 35273 59015
rect 35523 58969 35580 59015
rect 35626 58969 35683 59015
rect 35729 58969 35786 59015
rect 35832 58969 35889 59015
rect 35935 58969 35992 59015
rect 36038 58969 36095 59015
rect 36141 58969 36198 59015
rect 36244 58969 36301 59015
rect 36347 58969 36360 59015
rect 34964 58937 36360 58969
rect 34964 58880 35082 58937
rect 31336 58832 31349 58878
rect 33323 58832 33336 58878
rect 33484 58843 35082 58880
rect 30583 58767 30637 58813
rect 30683 58773 31040 58813
rect 33019 58829 33057 58832
rect 33109 58829 33237 58832
rect 33289 58829 33327 58832
rect 33019 58789 33327 58829
rect 33484 58797 33816 58843
rect 33862 58797 34002 58843
rect 34048 58797 34189 58843
rect 34235 58797 34376 58843
rect 34422 58797 34562 58843
rect 34608 58797 35082 58843
rect 36438 58925 36475 59065
rect 36521 58925 36554 59065
rect 33484 58789 35082 58797
rect 35294 58791 36266 58831
rect 36438 58825 36554 58925
rect 36640 59065 36773 59088
rect 36640 59016 36697 59065
rect 36640 58964 36678 59016
rect 36640 58925 36697 58964
rect 36743 58925 36773 59065
rect 38658 59067 38726 59078
rect 36924 59057 37685 59063
rect 36923 59056 37685 59057
rect 36923 59023 37931 59056
rect 36923 59015 36961 59023
rect 37013 59015 37172 59023
rect 37224 59015 37384 59023
rect 36841 58969 36854 59015
rect 36900 58971 36961 59015
rect 36900 58969 36971 58971
rect 37017 58969 37088 59015
rect 37134 58971 37172 59015
rect 37134 58969 37206 58971
rect 37252 58969 37324 59015
rect 37370 58971 37384 59015
rect 37436 59015 37595 59023
rect 37436 58971 37442 59015
rect 37370 58969 37442 58971
rect 37488 58971 37595 59015
rect 37647 59015 37931 59023
rect 37647 58971 37909 59015
rect 37488 58969 37909 58971
rect 37955 58969 38026 59015
rect 38072 58969 38143 59015
rect 38189 58969 38261 59015
rect 38307 58969 38379 59015
rect 38425 58969 38497 59015
rect 38543 58969 38556 59015
rect 36923 58937 37931 58969
rect 36924 58930 37685 58937
rect 36640 58905 36773 58925
rect 38658 58927 38669 59067
rect 38715 58927 38726 59067
rect 39014 59015 39323 59501
rect 39492 59587 39608 60039
rect 39923 60006 40085 60137
rect 39923 59954 39994 60006
rect 40046 59954 40085 60006
rect 39923 59914 40085 59954
rect 39737 59818 39865 59831
rect 39737 59791 39866 59818
rect 39737 59774 39775 59791
rect 39827 59774 39866 59791
rect 39727 59728 39740 59774
rect 39827 59739 39862 59774
rect 39786 59728 39862 59739
rect 39908 59728 39985 59774
rect 40031 59728 40108 59774
rect 40154 59728 40167 59774
rect 40246 59763 40362 60161
rect 42229 60022 44509 60063
rect 42229 59970 42312 60022
rect 42364 59970 44509 60022
rect 42229 59930 44509 59970
rect 44341 59886 44509 59930
rect 44341 59840 44358 59886
rect 44498 59840 44509 59886
rect 39737 59699 39866 59728
rect 40246 59717 40281 59763
rect 40327 59717 40362 59763
rect 40246 59680 40362 59717
rect 40718 59791 43524 59832
rect 44341 59829 44509 59840
rect 40718 59739 41935 59791
rect 41987 59739 43524 59791
rect 40718 59698 43524 59739
rect 44605 59774 44721 60161
rect 45400 60131 48379 60172
rect 45400 60117 47486 60131
rect 45400 60071 45464 60117
rect 45604 60079 47486 60117
rect 47538 60079 48379 60131
rect 45604 60071 48379 60079
rect 44901 60015 45241 60056
rect 45400 60038 48379 60071
rect 48557 60125 48596 60177
rect 48648 60125 48687 60177
rect 48557 60102 48687 60125
rect 50044 60211 50516 60257
rect 50562 60211 50703 60257
rect 50749 60211 50890 60257
rect 50936 60211 51076 60257
rect 51122 60211 51263 60257
rect 51309 60211 51657 60257
rect 51797 60247 52105 60287
rect 51797 60222 51835 60247
rect 51887 60222 52015 60247
rect 52067 60222 52105 60247
rect 54085 60281 54223 60327
rect 54269 60287 54540 60327
rect 54269 60281 54440 60287
rect 54085 60241 54440 60281
rect 54486 60241 54540 60287
rect 50044 60174 51657 60211
rect 51789 60176 51802 60222
rect 53776 60176 53789 60222
rect 50044 60117 50160 60174
rect 44901 59998 44939 60015
rect 44991 59998 45151 60015
rect 45203 59998 45241 60015
rect 44799 59952 44812 59998
rect 44858 59952 44925 59998
rect 44991 59963 45038 59998
rect 44971 59952 45038 59963
rect 45084 59952 45151 59998
rect 45203 59963 45264 59998
rect 45197 59952 45264 59963
rect 45310 59952 45323 59998
rect 48557 59962 48622 60102
rect 48668 59962 48687 60102
rect 49820 60085 50160 60117
rect 48765 60039 48778 60085
rect 48824 60039 48881 60085
rect 48927 60039 48984 60085
rect 49030 60039 49087 60085
rect 49133 60039 49190 60085
rect 49236 60039 49293 60085
rect 49339 60039 49396 60085
rect 49442 60039 49499 60085
rect 49545 60039 49602 60085
rect 49852 60039 50160 60085
rect 51589 60122 51657 60174
rect 51797 60154 52105 60176
rect 49820 59998 50160 60039
rect 50262 60015 50812 60056
rect 48557 59959 48687 59962
rect 44901 59923 45241 59952
rect 48557 59907 48596 59959
rect 48648 59907 48687 59959
rect 50262 59963 50300 60015
rect 50352 59998 50511 60015
rect 50563 59998 50722 60015
rect 50352 59963 50467 59998
rect 50563 59963 50571 59998
rect 50262 59952 50467 59963
rect 50513 59952 50571 59963
rect 50617 59952 50674 59998
rect 50720 59963 50722 59998
rect 50774 59998 50812 60015
rect 50774 59963 50777 59998
rect 50720 59952 50777 59963
rect 50823 59952 50880 59998
rect 50926 59952 50983 59998
rect 51029 59952 51086 59998
rect 51132 59952 51189 59998
rect 51235 59952 51292 59998
rect 51338 59952 51395 59998
rect 51441 59952 51454 59998
rect 50262 59923 50812 59952
rect 48557 59866 48687 59907
rect 48905 59861 49877 59892
rect 48765 59815 48778 59861
rect 48824 59815 48881 59861
rect 48927 59852 48984 59861
rect 48927 59815 48943 59852
rect 49030 59815 49087 59861
rect 49133 59852 49190 59861
rect 49133 59815 49154 59852
rect 49236 59815 49293 59861
rect 49339 59852 49396 59861
rect 49339 59815 49365 59852
rect 49442 59815 49499 59861
rect 49545 59852 49602 59861
rect 49545 59815 49576 59852
rect 49852 59815 49877 59861
rect 48905 59800 48943 59815
rect 48995 59800 49154 59815
rect 49206 59800 49365 59815
rect 49417 59800 49576 59815
rect 49628 59800 49787 59815
rect 49839 59800 49877 59815
rect 44605 59728 44812 59774
rect 44858 59728 44925 59774
rect 44971 59728 45038 59774
rect 45084 59728 45151 59774
rect 45197 59728 45264 59774
rect 45310 59728 45323 59774
rect 48905 59760 49877 59800
rect 51035 59777 51343 59817
rect 51035 59774 51073 59777
rect 51125 59774 51253 59777
rect 51305 59774 51343 59777
rect 43362 59691 43524 59698
rect 43362 59645 43373 59691
rect 43513 59645 43524 59691
rect 43362 59634 43524 59645
rect 45584 59714 48546 59750
rect 50454 59728 50467 59774
rect 50513 59728 50571 59774
rect 50617 59728 50674 59774
rect 50720 59728 50777 59774
rect 50823 59728 50880 59774
rect 50926 59728 50983 59774
rect 51029 59728 51073 59774
rect 51132 59728 51189 59774
rect 51235 59728 51253 59774
rect 51338 59728 51395 59774
rect 51441 59728 51454 59774
rect 45584 59668 45619 59714
rect 45665 59668 45777 59714
rect 45823 59668 45935 59714
rect 45981 59668 46093 59714
rect 46139 59668 46251 59714
rect 46297 59668 46409 59714
rect 46455 59668 46568 59714
rect 46614 59668 46726 59714
rect 46772 59668 46884 59714
rect 46930 59668 47042 59714
rect 47088 59668 47200 59714
rect 47246 59668 47358 59714
rect 47404 59668 47516 59714
rect 47562 59668 47675 59714
rect 47721 59668 47833 59714
rect 47879 59668 47991 59714
rect 48037 59668 48149 59714
rect 48195 59668 48307 59714
rect 48353 59668 48465 59714
rect 48511 59668 48546 59714
rect 51035 59725 51073 59728
rect 51125 59725 51253 59728
rect 51305 59725 51343 59728
rect 51035 59684 51343 59725
rect 51589 59700 51600 60122
rect 51646 59700 51657 60122
rect 54085 60123 54540 60241
rect 54085 60077 54440 60123
rect 54486 60077 54540 60123
rect 54085 60049 54540 60077
rect 53585 59998 54540 60049
rect 51789 59952 51802 59998
rect 53776 59960 54540 59998
rect 53776 59952 54440 59960
rect 53585 59930 54440 59952
rect 54085 59914 54440 59930
rect 54486 59914 54540 59960
rect 54085 59838 54540 59914
rect 51797 59784 52105 59824
rect 51797 59774 51835 59784
rect 51887 59774 52015 59784
rect 52067 59774 52105 59784
rect 54085 59792 54223 59838
rect 54269 59797 54540 59838
rect 54269 59792 54440 59797
rect 51789 59728 51802 59774
rect 53776 59728 53789 59774
rect 54085 59751 54440 59792
rect 54486 59751 54540 59797
rect 51589 59689 51657 59700
rect 51797 59691 52105 59728
rect 40215 59587 40523 59594
rect 40788 59587 42986 59601
rect 43753 59587 44514 59594
rect 39492 59564 42986 59587
rect 43704 59564 44514 59587
rect 39492 59553 44514 59564
rect 39492 59550 40253 59553
rect 39492 59504 39740 59550
rect 39786 59504 39862 59550
rect 39908 59504 39985 59550
rect 40031 59504 40108 59550
rect 40154 59504 40253 59550
rect 39492 59501 40253 59504
rect 40305 59501 40433 59553
rect 40485 59550 43790 59553
rect 40485 59504 40836 59550
rect 40882 59504 40994 59550
rect 41040 59504 41152 59550
rect 41198 59504 41310 59550
rect 41356 59504 41469 59550
rect 41515 59504 41627 59550
rect 41673 59504 41785 59550
rect 41831 59504 41943 59550
rect 41989 59504 42101 59550
rect 42147 59504 42259 59550
rect 42305 59504 42418 59550
rect 42464 59504 42576 59550
rect 42622 59504 42734 59550
rect 42780 59504 42892 59550
rect 42938 59504 43739 59550
rect 43785 59504 43790 59550
rect 40485 59501 43790 59504
rect 43842 59550 44001 59553
rect 43842 59504 43906 59550
rect 43952 59504 44001 59550
rect 43842 59501 44001 59504
rect 44053 59550 44213 59553
rect 44265 59550 44424 59553
rect 44053 59504 44071 59550
rect 44117 59504 44213 59550
rect 44282 59504 44424 59550
rect 44053 59501 44213 59504
rect 44265 59501 44424 59504
rect 44476 59501 44514 59553
rect 39492 59490 44514 59501
rect 39492 59467 42986 59490
rect 43704 59467 44514 59490
rect 39492 59015 39608 59467
rect 40215 59460 40523 59467
rect 40788 59453 42986 59467
rect 43753 59460 44514 59467
rect 44796 59587 45346 59594
rect 45584 59587 48546 59668
rect 54085 59674 54540 59751
rect 54085 59628 54223 59674
rect 54269 59634 54540 59674
rect 54269 59628 54440 59634
rect 54085 59594 54440 59628
rect 48800 59587 49982 59594
rect 50308 59587 50859 59594
rect 44796 59553 49982 59587
rect 44796 59550 44834 59553
rect 44886 59550 45045 59553
rect 45097 59550 45256 59553
rect 45308 59550 48838 59553
rect 44796 59504 44812 59550
rect 44886 59504 44925 59550
rect 44971 59504 45038 59550
rect 45097 59504 45151 59550
rect 45197 59504 45256 59550
rect 45310 59504 45619 59550
rect 45665 59504 45777 59550
rect 45823 59504 45935 59550
rect 45981 59504 46093 59550
rect 46139 59504 46251 59550
rect 46297 59504 46409 59550
rect 46455 59504 46568 59550
rect 46614 59504 46726 59550
rect 46772 59504 46884 59550
rect 46930 59504 47042 59550
rect 47088 59504 47200 59550
rect 47246 59504 47358 59550
rect 47404 59504 47516 59550
rect 47562 59504 47675 59550
rect 47721 59504 47833 59550
rect 47879 59504 47991 59550
rect 48037 59504 48149 59550
rect 48195 59504 48307 59550
rect 48353 59504 48465 59550
rect 48511 59504 48838 59550
rect 44796 59501 44834 59504
rect 44886 59501 45045 59504
rect 45097 59501 45256 59504
rect 45308 59501 48838 59504
rect 48890 59501 49048 59553
rect 49100 59501 49259 59553
rect 49311 59501 49471 59553
rect 49523 59501 49682 59553
rect 49734 59501 49892 59553
rect 49944 59501 49982 59553
rect 44796 59467 49982 59501
rect 50307 59553 50859 59587
rect 50307 59501 50346 59553
rect 50398 59550 50557 59553
rect 50609 59550 50768 59553
rect 50820 59550 50859 59553
rect 52278 59588 54440 59594
rect 54486 59588 54540 59634
rect 55927 60287 57736 60401
rect 55927 60244 56267 60287
rect 55927 60198 55961 60244
rect 56007 60241 56267 60244
rect 56313 60241 57736 60287
rect 56007 60198 57736 60241
rect 55927 60123 57736 60198
rect 55927 60081 56267 60123
rect 55927 60035 55961 60081
rect 56007 60077 56267 60081
rect 56313 60077 57736 60123
rect 56007 60035 57736 60077
rect 55927 59960 57736 60035
rect 55927 59917 56267 59960
rect 55927 59871 55961 59917
rect 56007 59914 56267 59917
rect 56313 59914 57736 59960
rect 56007 59871 57736 59914
rect 55927 59797 57736 59871
rect 55927 59754 56267 59797
rect 55927 59708 55961 59754
rect 56007 59751 56267 59754
rect 56313 59751 57736 59797
rect 56007 59708 57736 59751
rect 55927 59634 57736 59708
rect 52278 59553 54540 59588
rect 52278 59550 52316 59553
rect 52368 59550 52527 59553
rect 52579 59550 52738 59553
rect 52790 59550 52948 59553
rect 53000 59550 53159 59553
rect 53211 59550 53371 59553
rect 53423 59550 53582 59553
rect 53634 59550 53792 59553
rect 50398 59504 50467 59550
rect 50513 59504 50557 59550
rect 50617 59504 50674 59550
rect 50720 59504 50768 59550
rect 50823 59504 50880 59550
rect 50926 59504 50983 59550
rect 51029 59504 51086 59550
rect 51132 59504 51189 59550
rect 51235 59504 51292 59550
rect 51338 59504 51395 59550
rect 51441 59504 51454 59550
rect 51789 59504 51802 59550
rect 53776 59504 53792 59550
rect 50398 59501 50557 59504
rect 50609 59501 50768 59504
rect 50820 59501 50859 59504
rect 50307 59467 50859 59501
rect 44796 59460 45346 59467
rect 43362 59409 43524 59420
rect 39737 59326 39866 59355
rect 40246 59337 40362 59374
rect 43362 59363 43373 59409
rect 43513 59363 43524 59409
rect 43362 59356 43524 59363
rect 39727 59280 39740 59326
rect 39786 59315 39862 59326
rect 39827 59280 39862 59315
rect 39908 59280 39985 59326
rect 40031 59280 40108 59326
rect 40154 59280 40167 59326
rect 40246 59291 40281 59337
rect 40327 59291 40362 59337
rect 39737 59263 39775 59280
rect 39827 59263 39866 59280
rect 39737 59236 39866 59263
rect 39737 59223 39865 59236
rect 39923 59100 40085 59140
rect 39923 59048 39994 59100
rect 40046 59048 40085 59100
rect 39008 58969 39021 59015
rect 39067 58969 39144 59015
rect 39190 58969 39267 59015
rect 39313 58969 39326 59015
rect 39492 58969 39641 59015
rect 39687 58969 39730 59015
rect 39014 58937 39323 58969
rect 39492 58937 39608 58969
rect 37853 58825 38161 58830
rect 36438 58791 36953 58825
rect 37439 58791 38161 58825
rect 38658 58805 38726 58927
rect 39923 58917 40085 59048
rect 39809 58914 40085 58917
rect 39809 58906 39994 58914
rect 39809 58860 39844 58906
rect 39890 58862 39994 58906
rect 40046 58893 40085 58914
rect 40246 58893 40362 59291
rect 40718 59315 43524 59356
rect 45584 59386 48546 59467
rect 48800 59460 49982 59467
rect 50308 59460 50859 59467
rect 52278 59501 52316 59504
rect 52368 59501 52527 59504
rect 52579 59501 52738 59504
rect 52790 59501 52948 59504
rect 53000 59501 53159 59504
rect 53211 59501 53371 59504
rect 53423 59501 53582 59504
rect 53634 59501 53792 59504
rect 53844 59501 54003 59553
rect 54055 59501 54214 59553
rect 54266 59501 54540 59553
rect 52278 59466 54540 59501
rect 52278 59460 54440 59466
rect 45584 59340 45619 59386
rect 45665 59340 45777 59386
rect 45823 59340 45935 59386
rect 45981 59340 46093 59386
rect 46139 59340 46251 59386
rect 46297 59340 46409 59386
rect 46455 59340 46568 59386
rect 46614 59340 46726 59386
rect 46772 59340 46884 59386
rect 46930 59340 47042 59386
rect 47088 59340 47200 59386
rect 47246 59340 47358 59386
rect 47404 59340 47516 59386
rect 47562 59340 47675 59386
rect 47721 59340 47833 59386
rect 47879 59340 47991 59386
rect 48037 59340 48149 59386
rect 48195 59340 48307 59386
rect 48353 59340 48465 59386
rect 48511 59340 48546 59386
rect 54085 59426 54440 59460
rect 54085 59380 54223 59426
rect 54269 59420 54440 59426
rect 54486 59420 54540 59466
rect 54758 59553 55840 59594
rect 54758 59550 54855 59553
rect 54758 59504 54793 59550
rect 54839 59504 54855 59550
rect 54758 59501 54855 59504
rect 54907 59550 55066 59553
rect 54907 59504 54956 59550
rect 55002 59504 55066 59550
rect 54907 59501 55066 59504
rect 55118 59550 55278 59553
rect 55330 59550 55489 59553
rect 55164 59504 55278 59550
rect 55330 59504 55439 59550
rect 55485 59504 55489 59550
rect 55118 59501 55278 59504
rect 55330 59501 55489 59504
rect 55541 59550 55840 59553
rect 55541 59504 55599 59550
rect 55645 59504 55760 59550
rect 55806 59504 55840 59550
rect 55541 59501 55840 59504
rect 54758 59461 55840 59501
rect 55927 59588 56267 59634
rect 56313 59588 57736 59634
rect 55927 59466 57736 59588
rect 54817 59460 55579 59461
rect 54269 59380 54540 59420
rect 40718 59263 41935 59315
rect 41987 59263 43524 59315
rect 40718 59222 43524 59263
rect 44605 59280 44812 59326
rect 44858 59280 44925 59326
rect 44971 59280 45038 59326
rect 45084 59280 45151 59326
rect 45197 59280 45264 59326
rect 45310 59280 45323 59326
rect 45584 59304 48546 59340
rect 51035 59329 51343 59370
rect 51035 59326 51073 59329
rect 51125 59326 51253 59329
rect 51305 59326 51343 59329
rect 51589 59354 51657 59365
rect 44341 59214 44509 59225
rect 44341 59168 44358 59214
rect 44498 59168 44509 59214
rect 44341 59124 44509 59168
rect 42229 59084 44509 59124
rect 42229 59032 42312 59084
rect 42364 59032 44509 59084
rect 42229 58991 44509 59032
rect 44605 58893 44721 59280
rect 48905 59254 49877 59294
rect 50454 59280 50467 59326
rect 50513 59280 50571 59326
rect 50617 59280 50674 59326
rect 50720 59280 50777 59326
rect 50823 59280 50880 59326
rect 50926 59280 50983 59326
rect 51029 59280 51073 59326
rect 51132 59280 51189 59326
rect 51235 59280 51253 59326
rect 51338 59280 51395 59326
rect 51441 59280 51454 59326
rect 48905 59239 48943 59254
rect 48995 59239 49154 59254
rect 49206 59239 49365 59254
rect 49417 59239 49576 59254
rect 49628 59239 49787 59254
rect 49839 59239 49877 59254
rect 48765 59193 48778 59239
rect 48824 59193 48881 59239
rect 48927 59202 48943 59239
rect 48927 59193 48984 59202
rect 49030 59193 49087 59239
rect 49133 59202 49154 59239
rect 49133 59193 49190 59202
rect 49236 59193 49293 59239
rect 49339 59202 49365 59239
rect 49339 59193 49396 59202
rect 49442 59193 49499 59239
rect 49545 59202 49576 59239
rect 49545 59193 49602 59202
rect 49852 59193 49877 59239
rect 51035 59277 51073 59280
rect 51125 59277 51253 59280
rect 51305 59277 51343 59280
rect 51035 59237 51343 59277
rect 48557 59147 48687 59188
rect 48905 59162 49877 59193
rect 44901 59102 45241 59131
rect 44799 59056 44812 59102
rect 44858 59056 44925 59102
rect 44971 59091 45038 59102
rect 44991 59056 45038 59091
rect 45084 59056 45151 59102
rect 45197 59091 45264 59102
rect 45203 59056 45264 59091
rect 45310 59056 45323 59102
rect 48557 59095 48596 59147
rect 48648 59095 48687 59147
rect 48557 59092 48687 59095
rect 44901 59039 44939 59056
rect 44991 59039 45151 59056
rect 45203 59039 45241 59056
rect 44901 58998 45241 59039
rect 45400 58983 48379 59016
rect 45400 58937 45464 58983
rect 45604 58975 48379 58983
rect 45604 58937 47864 58975
rect 45400 58923 47864 58937
rect 47916 58923 48379 58975
rect 40046 58878 44918 58893
rect 45400 58882 48379 58923
rect 48557 58952 48622 59092
rect 48668 58952 48687 59092
rect 50262 59102 50812 59131
rect 50262 59091 50467 59102
rect 50513 59091 50571 59102
rect 49820 59015 50160 59056
rect 48765 58969 48778 59015
rect 48824 58969 48881 59015
rect 48927 58969 48984 59015
rect 49030 58969 49087 59015
rect 49133 58969 49190 59015
rect 49236 58969 49293 59015
rect 49339 58969 49396 59015
rect 49442 58969 49499 59015
rect 49545 58969 49602 59015
rect 49852 58969 50160 59015
rect 50262 59039 50300 59091
rect 50352 59056 50467 59091
rect 50563 59056 50571 59091
rect 50617 59056 50674 59102
rect 50720 59091 50777 59102
rect 50720 59056 50722 59091
rect 50352 59039 50511 59056
rect 50563 59039 50722 59056
rect 50774 59056 50777 59091
rect 50823 59056 50880 59102
rect 50926 59056 50983 59102
rect 51029 59056 51086 59102
rect 51132 59056 51189 59102
rect 51235 59056 51292 59102
rect 51338 59056 51395 59102
rect 51441 59056 51454 59102
rect 50774 59039 50812 59056
rect 50262 58998 50812 59039
rect 48557 58929 48687 58952
rect 49820 58937 50160 58969
rect 40046 58862 44812 58878
rect 39890 58860 44812 58862
rect 39809 58857 44812 58860
rect 39809 58811 43739 58857
rect 43785 58811 43906 58857
rect 43952 58811 44071 58857
rect 44117 58811 44236 58857
rect 44282 58832 44812 58857
rect 44858 58832 44925 58878
rect 44971 58832 45038 58878
rect 45084 58832 45151 58878
rect 45197 58832 45264 58878
rect 45310 58832 45323 58878
rect 48557 58877 48596 58929
rect 48648 58877 48687 58929
rect 48557 58837 48687 58877
rect 50044 58880 50160 58937
rect 51589 58932 51600 59354
rect 51646 58932 51657 59354
rect 51797 59326 52105 59363
rect 51789 59280 51802 59326
rect 53776 59280 53789 59326
rect 54085 59303 54540 59380
rect 51797 59270 51835 59280
rect 51887 59270 52015 59280
rect 52067 59270 52105 59280
rect 51797 59230 52105 59270
rect 54085 59262 54440 59303
rect 54085 59216 54223 59262
rect 54269 59257 54440 59262
rect 54486 59257 54540 59303
rect 54269 59216 54540 59257
rect 54085 59140 54540 59216
rect 54085 59124 54440 59140
rect 53585 59102 54440 59124
rect 51789 59056 51802 59102
rect 53776 59094 54440 59102
rect 54486 59094 54540 59140
rect 53776 59056 54540 59094
rect 53585 59005 54540 59056
rect 51589 58880 51657 58932
rect 54085 58977 54540 59005
rect 54085 58931 54440 58977
rect 54486 58931 54540 58977
rect 50044 58843 51657 58880
rect 51797 58878 52105 58900
rect 44282 58811 44918 58832
rect 38658 58791 39723 58805
rect 30683 58767 30855 58773
rect 30583 58727 30855 58767
rect 30901 58727 31040 58773
rect 33484 58760 34643 58789
rect 35260 58745 35273 58791
rect 35523 58745 35543 58791
rect 35626 58745 35683 58791
rect 35729 58745 35754 58791
rect 35832 58745 35889 58791
rect 35935 58745 35965 58791
rect 36038 58745 36095 58791
rect 36141 58745 36176 58791
rect 36244 58745 36301 58791
rect 36347 58745 36360 58791
rect 36438 58745 36854 58791
rect 36900 58745 36971 58791
rect 37017 58745 37088 58791
rect 37134 58745 37206 58791
rect 37252 58745 37324 58791
rect 37370 58745 37442 58791
rect 37488 58789 37909 58791
rect 37488 58745 37891 58789
rect 37955 58745 38026 58791
rect 38072 58789 38143 58791
rect 38123 58745 38143 58789
rect 38189 58745 38261 58791
rect 38307 58745 38379 58791
rect 38425 58745 38497 58791
rect 38543 58745 38556 58791
rect 38658 58745 39021 58791
rect 39067 58745 39144 58791
rect 39190 58745 39267 58791
rect 39313 58745 39641 58791
rect 39687 58745 39730 58791
rect 39809 58773 44918 58811
rect 48905 58791 49877 58831
rect 48765 58745 48778 58791
rect 48824 58745 48881 58791
rect 48927 58745 48943 58791
rect 49030 58745 49087 58791
rect 49133 58745 49154 58791
rect 49236 58745 49293 58791
rect 49339 58745 49365 58791
rect 49442 58745 49499 58791
rect 49545 58745 49576 58791
rect 49852 58745 49877 58791
rect 50044 58797 50516 58843
rect 50562 58797 50703 58843
rect 50749 58797 50890 58843
rect 50936 58797 51076 58843
rect 51122 58797 51263 58843
rect 51309 58797 51657 58843
rect 51789 58832 51802 58878
rect 53776 58832 53789 58878
rect 50044 58787 51657 58797
rect 50481 58760 51657 58787
rect 51797 58807 51835 58832
rect 51887 58807 52015 58832
rect 52067 58807 52105 58832
rect 51797 58767 52105 58807
rect 54085 58813 54540 58931
rect 54085 58773 54440 58813
rect 30583 58694 31040 58727
rect 35294 58739 35332 58745
rect 35384 58739 35543 58745
rect 35595 58739 35754 58745
rect 35806 58739 35965 58745
rect 36017 58739 36176 58745
rect 36228 58739 36266 58745
rect 34870 58694 35025 58701
rect 35294 58699 36266 58739
rect 36438 58705 36953 58745
rect 37439 58737 37891 58745
rect 37943 58737 38071 58745
rect 38123 58737 38161 58745
rect 37439 58705 38161 58737
rect 37853 58697 38161 58705
rect 27387 58601 27790 58653
rect 27842 58601 28001 58653
rect 28053 58601 28212 58653
rect 28264 58601 28423 58653
rect 28475 58601 28634 58653
rect 28686 58650 28845 58653
rect 28686 58604 28810 58650
rect 28686 58601 28845 58604
rect 28897 58601 29056 58653
rect 29108 58601 29196 58653
rect 27387 58487 29196 58601
rect 29283 58653 30365 58694
rect 29283 58650 29582 58653
rect 29283 58604 29317 58650
rect 29363 58604 29478 58650
rect 29524 58604 29582 58650
rect 29283 58601 29582 58604
rect 29634 58650 29793 58653
rect 29845 58650 30005 58653
rect 29634 58604 29638 58650
rect 29684 58604 29793 58650
rect 29845 58604 29959 58650
rect 29634 58601 29793 58604
rect 29845 58601 30005 58604
rect 30057 58650 30216 58653
rect 30057 58604 30121 58650
rect 30167 58604 30216 58650
rect 30057 58601 30216 58604
rect 30268 58650 30365 58653
rect 30268 58604 30284 58650
rect 30330 58604 30365 58650
rect 30268 58601 30365 58604
rect 29283 58561 30365 58601
rect 30583 58653 32842 58694
rect 30583 58650 30854 58653
rect 30583 58604 30637 58650
rect 30683 58604 30854 58650
rect 30583 58601 30854 58604
rect 30906 58601 31065 58653
rect 31117 58601 31276 58653
rect 31328 58601 31486 58653
rect 31538 58601 31697 58653
rect 31749 58601 31909 58653
rect 31961 58601 32120 58653
rect 32172 58601 32330 58653
rect 32382 58601 32541 58653
rect 32593 58601 32752 58653
rect 32804 58601 32842 58653
rect 29544 58560 30306 58561
rect 30583 58560 32842 58601
rect 34717 58653 35025 58694
rect 38658 58685 39723 58745
rect 48905 58739 48943 58745
rect 48995 58739 49154 58745
rect 49206 58739 49365 58745
rect 49417 58739 49576 58745
rect 49628 58739 49787 58745
rect 49839 58739 49877 58745
rect 48905 58699 49877 58739
rect 54085 58727 54223 58773
rect 54269 58767 54440 58773
rect 54486 58767 54540 58813
rect 54269 58727 54540 58767
rect 50099 58694 50255 58701
rect 54085 58694 54540 58727
rect 55927 59420 56267 59466
rect 56313 59420 57736 59466
rect 55927 59344 57736 59420
rect 55927 59298 55961 59344
rect 56007 59303 57736 59344
rect 56007 59298 56267 59303
rect 55927 59257 56267 59298
rect 56313 59257 57736 59303
rect 55927 59181 57736 59257
rect 55927 59135 55961 59181
rect 56007 59140 57736 59181
rect 56007 59135 56267 59140
rect 55927 59094 56267 59135
rect 56313 59094 57736 59140
rect 55927 59017 57736 59094
rect 55927 58971 55961 59017
rect 56007 58977 57736 59017
rect 56007 58971 56267 58977
rect 55927 58931 56267 58971
rect 56313 58931 57736 58977
rect 55927 58854 57736 58931
rect 55927 58808 55961 58854
rect 56007 58813 57736 58854
rect 56007 58808 56267 58813
rect 55927 58767 56267 58808
rect 56313 58767 57736 58813
rect 34717 58601 34755 58653
rect 34807 58650 34935 58653
rect 34807 58604 34916 58650
rect 34807 58601 34935 58604
rect 34987 58601 35025 58653
rect 34717 58560 35025 58601
rect 50099 58653 50408 58694
rect 50099 58601 50138 58653
rect 50190 58650 50318 58653
rect 50206 58604 50318 58650
rect 50190 58601 50318 58604
rect 50370 58601 50408 58653
rect 27387 58441 28810 58487
rect 28856 58444 29196 58487
rect 28856 58441 29116 58444
rect 27387 58398 29116 58441
rect 29162 58398 29196 58444
rect 27387 58323 29196 58398
rect 27387 58277 28810 58323
rect 28856 58281 29196 58323
rect 28856 58277 29116 58281
rect 27387 58235 29116 58277
rect 29162 58235 29196 58281
rect 27387 58160 29196 58235
rect 27387 58114 28810 58160
rect 28856 58117 29196 58160
rect 28856 58114 29116 58117
rect 27387 58071 29116 58114
rect 29162 58071 29196 58117
rect 27387 57997 29196 58071
rect 27387 57951 28810 57997
rect 28856 57954 29196 57997
rect 28856 57951 29116 57954
rect 27387 57908 29116 57951
rect 29162 57908 29196 57954
rect 27387 57834 29196 57908
rect 27387 57788 28810 57834
rect 28856 57788 29196 57834
rect 30583 58527 31040 58560
rect 34870 58553 35025 58560
rect 30583 58487 30855 58527
rect 30583 58441 30637 58487
rect 30683 58481 30855 58487
rect 30901 58481 31040 58527
rect 35294 58515 36266 58555
rect 37853 58549 38161 58557
rect 35294 58509 35332 58515
rect 35384 58509 35543 58515
rect 35595 58509 35754 58515
rect 35806 58509 35965 58515
rect 36017 58509 36176 58515
rect 36228 58509 36266 58515
rect 36438 58509 36953 58549
rect 37439 58517 38161 58549
rect 37439 58509 37891 58517
rect 37943 58509 38071 58517
rect 38123 58509 38161 58517
rect 38658 58509 39723 58569
rect 50099 58560 50408 58601
rect 52278 58653 54540 58694
rect 52278 58601 52316 58653
rect 52368 58601 52527 58653
rect 52579 58601 52738 58653
rect 52790 58601 52948 58653
rect 53000 58601 53159 58653
rect 53211 58601 53371 58653
rect 53423 58601 53582 58653
rect 53634 58601 53792 58653
rect 53844 58601 54003 58653
rect 54055 58601 54214 58653
rect 54266 58650 54540 58653
rect 54266 58604 54440 58650
rect 54486 58604 54540 58650
rect 54266 58601 54540 58604
rect 52278 58560 54540 58601
rect 54758 58653 55840 58694
rect 54758 58650 54855 58653
rect 54758 58604 54793 58650
rect 54839 58604 54855 58650
rect 54758 58601 54855 58604
rect 54907 58650 55066 58653
rect 54907 58604 54956 58650
rect 55002 58604 55066 58650
rect 54907 58601 55066 58604
rect 55118 58650 55278 58653
rect 55330 58650 55489 58653
rect 55164 58604 55278 58650
rect 55330 58604 55439 58650
rect 55485 58604 55489 58650
rect 55118 58601 55278 58604
rect 55330 58601 55489 58604
rect 55541 58650 55840 58653
rect 55541 58604 55599 58650
rect 55645 58604 55760 58650
rect 55806 58604 55840 58650
rect 55541 58601 55840 58604
rect 54758 58561 55840 58601
rect 55927 58653 57736 58767
rect 55927 58601 56015 58653
rect 56067 58601 56226 58653
rect 56278 58650 56437 58653
rect 56313 58604 56437 58650
rect 56278 58601 56437 58604
rect 56489 58601 56648 58653
rect 56700 58601 56859 58653
rect 56911 58601 57070 58653
rect 57122 58601 57281 58653
rect 57333 58601 57736 58653
rect 54817 58560 55579 58561
rect 48905 58515 49877 58555
rect 50099 58553 50255 58560
rect 48905 58509 48943 58515
rect 48995 58509 49154 58515
rect 49206 58509 49365 58515
rect 49417 58509 49576 58515
rect 49628 58509 49787 58515
rect 49839 58509 49877 58515
rect 30683 58441 31040 58481
rect 33484 58465 34643 58494
rect 30583 58364 31040 58441
rect 33019 58425 33327 58465
rect 33019 58422 33057 58425
rect 33109 58422 33237 58425
rect 33289 58422 33327 58425
rect 33484 58457 35082 58465
rect 35260 58463 35273 58509
rect 35523 58463 35543 58509
rect 35626 58463 35683 58509
rect 35729 58463 35754 58509
rect 35832 58463 35889 58509
rect 35935 58463 35965 58509
rect 36038 58463 36095 58509
rect 36141 58463 36176 58509
rect 36244 58463 36301 58509
rect 36347 58463 36360 58509
rect 36438 58463 36854 58509
rect 36900 58463 36971 58509
rect 37017 58463 37088 58509
rect 37134 58463 37206 58509
rect 37252 58463 37324 58509
rect 37370 58463 37442 58509
rect 37488 58465 37891 58509
rect 37488 58463 37909 58465
rect 37955 58463 38026 58509
rect 38123 58465 38143 58509
rect 38072 58463 38143 58465
rect 38189 58463 38261 58509
rect 38307 58463 38379 58509
rect 38425 58463 38497 58509
rect 38543 58463 38556 58509
rect 38658 58463 39021 58509
rect 39067 58463 39144 58509
rect 39190 58463 39267 58509
rect 39313 58463 39641 58509
rect 39687 58463 39730 58509
rect 31336 58376 31349 58422
rect 33323 58376 33336 58422
rect 33484 58411 33816 58457
rect 33862 58411 34002 58457
rect 34048 58411 34189 58457
rect 34235 58411 34376 58457
rect 34422 58411 34562 58457
rect 34608 58411 35082 58457
rect 35294 58423 36266 58463
rect 36438 58429 36953 58463
rect 37439 58429 38161 58463
rect 30583 58323 30855 58364
rect 30583 58277 30637 58323
rect 30683 58318 30855 58323
rect 30901 58318 31040 58364
rect 33019 58373 33057 58376
rect 33109 58373 33237 58376
rect 33289 58373 33327 58376
rect 33019 58332 33327 58373
rect 33484 58374 35082 58411
rect 30683 58277 31040 58318
rect 30583 58249 31040 58277
rect 33484 58292 33552 58374
rect 30583 58201 31493 58249
rect 30583 58160 30855 58201
rect 30583 58114 30637 58160
rect 30683 58155 30855 58160
rect 30901 58198 31493 58201
rect 30901 58155 31349 58198
rect 30683 58152 31349 58155
rect 33323 58152 33336 58198
rect 30683 58130 31493 58152
rect 30683 58114 31040 58130
rect 30583 58038 31040 58114
rect 30583 57997 30855 58038
rect 30583 57951 30637 57997
rect 30683 57992 30855 57997
rect 30901 57992 31040 58038
rect 30683 57951 31040 57992
rect 33019 57977 33327 58017
rect 33019 57974 33057 57977
rect 33109 57974 33237 57977
rect 33289 57974 33327 57977
rect 30583 57874 31040 57951
rect 31336 57928 31349 57974
rect 33323 57928 33336 57974
rect 33019 57925 33057 57928
rect 33109 57925 33237 57928
rect 33289 57925 33327 57928
rect 33019 57884 33327 57925
rect 30583 57834 30855 57874
rect 27387 57666 29196 57788
rect 27387 57620 28810 57666
rect 28856 57620 29196 57666
rect 29283 57753 30365 57794
rect 29283 57750 29582 57753
rect 29283 57704 29317 57750
rect 29363 57704 29478 57750
rect 29524 57704 29582 57750
rect 29283 57701 29582 57704
rect 29634 57750 29793 57753
rect 29845 57750 30005 57753
rect 29634 57704 29638 57750
rect 29684 57704 29793 57750
rect 29845 57704 29959 57750
rect 29634 57701 29793 57704
rect 29845 57701 30005 57704
rect 30057 57750 30216 57753
rect 30057 57704 30121 57750
rect 30167 57704 30216 57750
rect 30057 57701 30216 57704
rect 30268 57750 30365 57753
rect 30268 57704 30284 57750
rect 30330 57704 30365 57750
rect 30268 57701 30365 57704
rect 29283 57661 30365 57701
rect 30583 57788 30637 57834
rect 30683 57828 30855 57834
rect 30901 57828 31040 57874
rect 33484 57870 33495 58292
rect 33541 57870 33552 58292
rect 34964 58317 35082 58374
rect 36438 58329 36554 58429
rect 37853 58424 38161 58429
rect 38658 58449 39723 58463
rect 34964 58285 36360 58317
rect 34228 58215 34718 58256
rect 34228 58198 34267 58215
rect 34319 58198 34447 58215
rect 34499 58198 34627 58215
rect 33671 58152 33684 58198
rect 33730 58152 33787 58198
rect 33833 58152 33890 58198
rect 33936 58152 33993 58198
rect 34039 58152 34096 58198
rect 34142 58152 34199 58198
rect 34245 58163 34267 58198
rect 34245 58152 34302 58163
rect 34348 58152 34405 58198
rect 34499 58163 34508 58198
rect 34451 58152 34508 58163
rect 34554 58152 34612 58198
rect 34679 58163 34718 58215
rect 34964 58239 35273 58285
rect 35523 58239 35580 58285
rect 35626 58239 35683 58285
rect 35729 58239 35786 58285
rect 35832 58239 35889 58285
rect 35935 58239 35992 58285
rect 36038 58239 36095 58285
rect 36141 58239 36198 58285
rect 36244 58239 36301 58285
rect 36347 58239 36360 58285
rect 34964 58195 36360 58239
rect 34658 58152 34718 58163
rect 34228 58123 34718 58152
rect 36438 58189 36475 58329
rect 36521 58189 36554 58329
rect 35294 58061 36266 58095
rect 36438 58086 36554 58189
rect 36640 58329 36773 58349
rect 36640 58290 36697 58329
rect 36640 58238 36678 58290
rect 36640 58189 36697 58238
rect 36743 58189 36773 58329
rect 38658 58327 38726 58449
rect 39809 58443 44918 58481
rect 48765 58463 48778 58509
rect 48824 58463 48881 58509
rect 48927 58463 48943 58509
rect 49030 58463 49087 58509
rect 49133 58463 49154 58509
rect 49236 58463 49293 58509
rect 49339 58463 49365 58509
rect 49442 58463 49499 58509
rect 49545 58463 49576 58509
rect 49852 58463 49877 58509
rect 54085 58527 54540 58560
rect 50481 58467 51657 58494
rect 39809 58397 43739 58443
rect 43785 58397 43906 58443
rect 43952 58397 44071 58443
rect 44117 58397 44236 58443
rect 44282 58422 44918 58443
rect 48905 58423 49877 58463
rect 50044 58457 51657 58467
rect 44282 58397 44812 58422
rect 39809 58394 44812 58397
rect 39809 58348 39844 58394
rect 39890 58392 44812 58394
rect 39890 58348 39994 58392
rect 39809 58340 39994 58348
rect 40046 58376 44812 58392
rect 44858 58376 44925 58422
rect 44971 58376 45038 58422
rect 45084 58376 45151 58422
rect 45197 58376 45264 58422
rect 45310 58376 45323 58422
rect 48557 58377 48687 58417
rect 40046 58361 44918 58376
rect 40046 58340 40085 58361
rect 39809 58337 40085 58340
rect 36924 58317 37685 58324
rect 36923 58285 37931 58317
rect 36841 58239 36854 58285
rect 36900 58283 36971 58285
rect 36900 58239 36961 58283
rect 37017 58239 37088 58285
rect 37134 58283 37206 58285
rect 37134 58239 37172 58283
rect 37252 58239 37324 58285
rect 37370 58283 37442 58285
rect 37370 58239 37384 58283
rect 36923 58231 36961 58239
rect 37013 58231 37172 58239
rect 37224 58231 37384 58239
rect 37436 58239 37442 58283
rect 37488 58283 37909 58285
rect 37488 58239 37595 58283
rect 37436 58231 37595 58239
rect 37647 58239 37909 58283
rect 37955 58239 38026 58285
rect 38072 58239 38143 58285
rect 38189 58239 38261 58285
rect 38307 58239 38379 58285
rect 38425 58239 38497 58285
rect 38543 58239 38556 58285
rect 37647 58231 37931 58239
rect 36923 58198 37931 58231
rect 36923 58197 37685 58198
rect 36924 58191 37685 58197
rect 36640 58166 36773 58189
rect 38658 58187 38669 58327
rect 38715 58187 38726 58327
rect 39014 58285 39323 58317
rect 39492 58285 39608 58317
rect 39008 58239 39021 58285
rect 39067 58239 39144 58285
rect 39190 58239 39267 58285
rect 39313 58239 39326 58285
rect 39492 58239 39641 58285
rect 39687 58239 39730 58285
rect 38658 58176 38726 58187
rect 36438 58061 36953 58086
rect 37439 58083 37931 58086
rect 37439 58061 38161 58083
rect 35260 58015 35273 58061
rect 35523 58055 35580 58061
rect 35523 58015 35543 58055
rect 35626 58015 35683 58061
rect 35729 58055 35786 58061
rect 35729 58015 35754 58055
rect 35832 58015 35889 58061
rect 35935 58055 35992 58061
rect 35935 58015 35965 58055
rect 36038 58015 36095 58061
rect 36141 58055 36198 58061
rect 36141 58015 36176 58055
rect 36244 58015 36301 58061
rect 36347 58015 36360 58061
rect 36438 58015 36854 58061
rect 36900 58015 36971 58061
rect 37017 58015 37088 58061
rect 37134 58015 37206 58061
rect 37252 58015 37324 58061
rect 37370 58015 37442 58061
rect 37488 58043 37909 58061
rect 37488 58015 37891 58043
rect 37955 58015 38026 58061
rect 38072 58043 38143 58061
rect 38123 58015 38143 58043
rect 38189 58015 38261 58061
rect 38307 58015 38379 58061
rect 38425 58015 38497 58061
rect 38543 58015 38556 58061
rect 33781 57974 34089 58009
rect 35294 58003 35332 58015
rect 35384 58003 35543 58015
rect 35595 58003 35754 58015
rect 35806 58003 35965 58015
rect 36017 58003 36176 58015
rect 36228 58003 36266 58015
rect 33671 57928 33684 57974
rect 33730 57928 33787 57974
rect 33833 57969 33890 57974
rect 33871 57928 33890 57969
rect 33936 57928 33993 57974
rect 34039 57969 34096 57974
rect 34051 57928 34096 57969
rect 34142 57928 34199 57974
rect 34245 57928 34302 57974
rect 34348 57928 34405 57974
rect 34451 57928 34508 57974
rect 34554 57928 34612 57974
rect 34658 57928 34671 57974
rect 35294 57963 36266 58003
rect 36438 57966 36953 58015
rect 37439 57991 37891 58015
rect 37943 57991 38071 58015
rect 38123 57991 38161 58015
rect 37439 57966 38161 57991
rect 37853 57950 38161 57966
rect 33781 57917 33819 57928
rect 33871 57917 33999 57928
rect 34051 57917 34089 57928
rect 33781 57876 34089 57917
rect 33484 57859 33552 57870
rect 30683 57794 31040 57828
rect 30683 57788 32842 57794
rect 30583 57753 32842 57788
rect 34247 57787 35008 57794
rect 30583 57701 30854 57753
rect 30906 57701 31065 57753
rect 31117 57701 31276 57753
rect 31328 57750 31486 57753
rect 31538 57750 31697 57753
rect 31749 57750 31909 57753
rect 31961 57750 32120 57753
rect 32172 57750 32330 57753
rect 32382 57750 32541 57753
rect 32593 57750 32752 57753
rect 32804 57750 32842 57753
rect 34246 57753 35008 57787
rect 34246 57750 34284 57753
rect 34336 57750 34495 57753
rect 34547 57750 34707 57753
rect 31328 57704 31349 57750
rect 33323 57704 33336 57750
rect 33671 57704 33684 57750
rect 33730 57704 33787 57750
rect 33833 57704 33890 57750
rect 33936 57704 33993 57750
rect 34039 57704 34096 57750
rect 34142 57704 34199 57750
rect 34245 57704 34284 57750
rect 34348 57704 34405 57750
rect 34451 57704 34495 57750
rect 34554 57704 34612 57750
rect 34658 57704 34707 57750
rect 31328 57701 31486 57704
rect 31538 57701 31697 57704
rect 31749 57701 31909 57704
rect 31961 57701 32120 57704
rect 32172 57701 32330 57704
rect 32382 57701 32541 57704
rect 32593 57701 32752 57704
rect 32804 57701 32842 57704
rect 30583 57666 32842 57701
rect 34246 57701 34284 57704
rect 34336 57701 34495 57704
rect 34547 57701 34707 57704
rect 34759 57701 34918 57753
rect 34970 57701 35008 57753
rect 34246 57667 35008 57701
rect 29544 57660 30306 57661
rect 27387 57544 29196 57620
rect 27387 57503 29116 57544
rect 27387 57457 28810 57503
rect 28856 57498 29116 57503
rect 29162 57498 29196 57544
rect 28856 57457 29196 57498
rect 27387 57381 29196 57457
rect 27387 57340 29116 57381
rect 27387 57294 28810 57340
rect 28856 57335 29116 57340
rect 29162 57335 29196 57381
rect 28856 57294 29196 57335
rect 27387 57217 29196 57294
rect 27387 57177 29116 57217
rect 27387 57131 28810 57177
rect 28856 57171 29116 57177
rect 29162 57171 29196 57217
rect 28856 57131 29196 57171
rect 27387 57054 29196 57131
rect 27387 57013 29116 57054
rect 27387 56967 28810 57013
rect 28856 57008 29116 57013
rect 29162 57008 29196 57054
rect 28856 56967 29196 57008
rect 27387 56853 29196 56967
rect 30583 57620 30637 57666
rect 30683 57660 32842 57666
rect 34247 57660 35008 57667
rect 35182 57787 36364 57794
rect 35182 57753 36958 57787
rect 35182 57701 35220 57753
rect 35272 57701 35430 57753
rect 35482 57701 35641 57753
rect 35693 57701 35853 57753
rect 35905 57701 36064 57753
rect 36116 57701 36274 57753
rect 36326 57750 36958 57753
rect 36326 57704 36489 57750
rect 36723 57704 36958 57750
rect 36326 57701 36958 57704
rect 35182 57667 36958 57701
rect 37946 57753 38842 57794
rect 37946 57750 38330 57753
rect 38382 57750 38541 57753
rect 37946 57704 37957 57750
rect 38473 57704 38541 57750
rect 37946 57701 38330 57704
rect 38382 57701 38541 57704
rect 38593 57701 38752 57753
rect 38804 57701 38842 57753
rect 35182 57660 36364 57667
rect 37946 57660 38842 57701
rect 39014 57753 39323 58239
rect 39014 57701 39052 57753
rect 39104 57750 39232 57753
rect 39108 57704 39220 57750
rect 39104 57701 39232 57704
rect 39284 57701 39323 57753
rect 30683 57626 31040 57660
rect 30683 57620 30855 57626
rect 30583 57580 30855 57620
rect 30901 57580 31040 57626
rect 30583 57503 31040 57580
rect 33484 57584 33552 57595
rect 33019 57529 33327 57570
rect 33019 57526 33057 57529
rect 33109 57526 33237 57529
rect 33289 57526 33327 57529
rect 30583 57457 30637 57503
rect 30683 57462 31040 57503
rect 31336 57480 31349 57526
rect 33323 57480 33336 57526
rect 30683 57457 30855 57462
rect 30583 57416 30855 57457
rect 30901 57416 31040 57462
rect 33019 57477 33057 57480
rect 33109 57477 33237 57480
rect 33289 57477 33327 57480
rect 33019 57437 33327 57477
rect 30583 57340 31040 57416
rect 30583 57294 30637 57340
rect 30683 57324 31040 57340
rect 30683 57302 31493 57324
rect 30683 57299 31349 57302
rect 30683 57294 30855 57299
rect 30583 57253 30855 57294
rect 30901 57256 31349 57299
rect 33323 57256 33336 57302
rect 30901 57253 31493 57256
rect 30583 57205 31493 57253
rect 30583 57177 31040 57205
rect 30583 57131 30637 57177
rect 30683 57136 31040 57177
rect 30683 57131 30855 57136
rect 30583 57090 30855 57131
rect 30901 57090 31040 57136
rect 33484 57162 33495 57584
rect 33541 57162 33552 57584
rect 33781 57537 34089 57578
rect 33781 57526 33819 57537
rect 33871 57526 33999 57537
rect 34051 57526 34089 57537
rect 33671 57480 33684 57526
rect 33730 57480 33787 57526
rect 33871 57485 33890 57526
rect 33833 57480 33890 57485
rect 33936 57480 33993 57526
rect 34051 57485 34096 57526
rect 34039 57480 34096 57485
rect 34142 57480 34199 57526
rect 34245 57480 34302 57526
rect 34348 57480 34405 57526
rect 34451 57480 34508 57526
rect 34554 57480 34612 57526
rect 34658 57480 34671 57526
rect 33781 57445 34089 57480
rect 35294 57451 36266 57491
rect 37853 57488 38161 57504
rect 35294 57439 35332 57451
rect 35384 57439 35543 57451
rect 35595 57439 35754 57451
rect 35806 57439 35965 57451
rect 36017 57439 36176 57451
rect 36228 57439 36266 57451
rect 36438 57439 36953 57488
rect 37439 57463 38161 57488
rect 37439 57439 37891 57463
rect 37943 57439 38071 57463
rect 38123 57439 38161 57463
rect 35260 57393 35273 57439
rect 35523 57399 35543 57439
rect 35523 57393 35580 57399
rect 35626 57393 35683 57439
rect 35729 57399 35754 57439
rect 35729 57393 35786 57399
rect 35832 57393 35889 57439
rect 35935 57399 35965 57439
rect 35935 57393 35992 57399
rect 36038 57393 36095 57439
rect 36141 57399 36176 57439
rect 36141 57393 36198 57399
rect 36244 57393 36301 57439
rect 36347 57393 36360 57439
rect 36438 57393 36854 57439
rect 36900 57393 36971 57439
rect 37017 57393 37088 57439
rect 37134 57393 37206 57439
rect 37252 57393 37324 57439
rect 37370 57393 37442 57439
rect 37488 57411 37891 57439
rect 37488 57393 37909 57411
rect 37955 57393 38026 57439
rect 38123 57411 38143 57439
rect 38072 57393 38143 57411
rect 38189 57393 38261 57439
rect 38307 57393 38379 57439
rect 38425 57393 38497 57439
rect 38543 57393 38556 57439
rect 35294 57359 36266 57393
rect 36438 57368 36953 57393
rect 37439 57371 38161 57393
rect 37439 57368 37931 57371
rect 34228 57302 34718 57331
rect 33671 57256 33684 57302
rect 33730 57256 33787 57302
rect 33833 57256 33890 57302
rect 33936 57256 33993 57302
rect 34039 57256 34096 57302
rect 34142 57256 34199 57302
rect 34245 57291 34302 57302
rect 34245 57256 34267 57291
rect 34348 57256 34405 57302
rect 34451 57291 34508 57302
rect 34499 57256 34508 57291
rect 34554 57256 34612 57302
rect 34658 57291 34718 57302
rect 34228 57239 34267 57256
rect 34319 57239 34447 57256
rect 34499 57239 34627 57256
rect 34679 57239 34718 57291
rect 36438 57265 36554 57368
rect 34228 57198 34718 57239
rect 34964 57215 36360 57259
rect 30583 57013 31040 57090
rect 33019 57081 33327 57122
rect 33019 57078 33057 57081
rect 33109 57078 33237 57081
rect 33289 57078 33327 57081
rect 33484 57080 33552 57162
rect 34964 57169 35273 57215
rect 35523 57169 35580 57215
rect 35626 57169 35683 57215
rect 35729 57169 35786 57215
rect 35832 57169 35889 57215
rect 35935 57169 35992 57215
rect 36038 57169 36095 57215
rect 36141 57169 36198 57215
rect 36244 57169 36301 57215
rect 36347 57169 36360 57215
rect 34964 57137 36360 57169
rect 34964 57080 35082 57137
rect 31336 57032 31349 57078
rect 33323 57032 33336 57078
rect 33484 57043 35082 57080
rect 30583 56967 30637 57013
rect 30683 56973 31040 57013
rect 33019 57029 33057 57032
rect 33109 57029 33237 57032
rect 33289 57029 33327 57032
rect 33019 56989 33327 57029
rect 33484 56997 33816 57043
rect 33862 56997 34002 57043
rect 34048 56997 34189 57043
rect 34235 56997 34376 57043
rect 34422 56997 34562 57043
rect 34608 56997 35082 57043
rect 36438 57125 36475 57265
rect 36521 57125 36554 57265
rect 33484 56989 35082 56997
rect 35294 56991 36266 57031
rect 36438 57025 36554 57125
rect 36640 57265 36773 57288
rect 36640 57216 36697 57265
rect 36640 57164 36678 57216
rect 36640 57125 36697 57164
rect 36743 57125 36773 57265
rect 38658 57267 38726 57278
rect 36924 57257 37685 57263
rect 36923 57256 37685 57257
rect 36923 57223 37931 57256
rect 36923 57215 36961 57223
rect 37013 57215 37172 57223
rect 37224 57215 37384 57223
rect 36841 57169 36854 57215
rect 36900 57171 36961 57215
rect 36900 57169 36971 57171
rect 37017 57169 37088 57215
rect 37134 57171 37172 57215
rect 37134 57169 37206 57171
rect 37252 57169 37324 57215
rect 37370 57171 37384 57215
rect 37436 57215 37595 57223
rect 37436 57171 37442 57215
rect 37370 57169 37442 57171
rect 37488 57171 37595 57215
rect 37647 57215 37931 57223
rect 37647 57171 37909 57215
rect 37488 57169 37909 57171
rect 37955 57169 38026 57215
rect 38072 57169 38143 57215
rect 38189 57169 38261 57215
rect 38307 57169 38379 57215
rect 38425 57169 38497 57215
rect 38543 57169 38556 57215
rect 36923 57137 37931 57169
rect 36924 57130 37685 57137
rect 36640 57105 36773 57125
rect 38658 57127 38669 57267
rect 38715 57127 38726 57267
rect 39014 57215 39323 57701
rect 39492 57787 39608 58239
rect 39923 58206 40085 58337
rect 39923 58154 39994 58206
rect 40046 58154 40085 58206
rect 39923 58114 40085 58154
rect 39737 58018 39865 58031
rect 39737 57991 39866 58018
rect 39737 57974 39775 57991
rect 39827 57974 39866 57991
rect 39727 57928 39740 57974
rect 39827 57939 39862 57974
rect 39786 57928 39862 57939
rect 39908 57928 39985 57974
rect 40031 57928 40108 57974
rect 40154 57928 40167 57974
rect 40246 57963 40362 58361
rect 42229 58222 44509 58263
rect 42229 58170 42312 58222
rect 42364 58170 44509 58222
rect 42229 58130 44509 58170
rect 44341 58086 44509 58130
rect 44341 58040 44358 58086
rect 44498 58040 44509 58086
rect 39737 57899 39866 57928
rect 40246 57917 40281 57963
rect 40327 57917 40362 57963
rect 40246 57880 40362 57917
rect 40718 57991 43524 58032
rect 44341 58029 44509 58040
rect 40718 57939 41935 57991
rect 41987 57939 43524 57991
rect 40718 57898 43524 57939
rect 44605 57974 44721 58361
rect 45400 58331 48379 58372
rect 45400 58317 48241 58331
rect 45400 58271 45464 58317
rect 45604 58279 48241 58317
rect 48293 58279 48379 58331
rect 45604 58271 48379 58279
rect 44901 58215 45241 58256
rect 45400 58238 48379 58271
rect 48557 58325 48596 58377
rect 48648 58325 48687 58377
rect 48557 58302 48687 58325
rect 50044 58411 50516 58457
rect 50562 58411 50703 58457
rect 50749 58411 50890 58457
rect 50936 58411 51076 58457
rect 51122 58411 51263 58457
rect 51309 58411 51657 58457
rect 51797 58447 52105 58487
rect 51797 58422 51835 58447
rect 51887 58422 52015 58447
rect 52067 58422 52105 58447
rect 54085 58481 54223 58527
rect 54269 58487 54540 58527
rect 54269 58481 54440 58487
rect 54085 58441 54440 58481
rect 54486 58441 54540 58487
rect 50044 58374 51657 58411
rect 51789 58376 51802 58422
rect 53776 58376 53789 58422
rect 50044 58317 50160 58374
rect 44901 58198 44939 58215
rect 44991 58198 45151 58215
rect 45203 58198 45241 58215
rect 44799 58152 44812 58198
rect 44858 58152 44925 58198
rect 44991 58163 45038 58198
rect 44971 58152 45038 58163
rect 45084 58152 45151 58198
rect 45203 58163 45264 58198
rect 45197 58152 45264 58163
rect 45310 58152 45323 58198
rect 48557 58162 48622 58302
rect 48668 58162 48687 58302
rect 49820 58285 50160 58317
rect 48765 58239 48778 58285
rect 48824 58239 48881 58285
rect 48927 58239 48984 58285
rect 49030 58239 49087 58285
rect 49133 58239 49190 58285
rect 49236 58239 49293 58285
rect 49339 58239 49396 58285
rect 49442 58239 49499 58285
rect 49545 58239 49602 58285
rect 49852 58239 50160 58285
rect 51589 58322 51657 58374
rect 51797 58354 52105 58376
rect 49820 58198 50160 58239
rect 50262 58215 50812 58256
rect 48557 58159 48687 58162
rect 44901 58123 45241 58152
rect 48557 58107 48596 58159
rect 48648 58107 48687 58159
rect 50262 58163 50300 58215
rect 50352 58198 50511 58215
rect 50563 58198 50722 58215
rect 50352 58163 50467 58198
rect 50563 58163 50571 58198
rect 50262 58152 50467 58163
rect 50513 58152 50571 58163
rect 50617 58152 50674 58198
rect 50720 58163 50722 58198
rect 50774 58198 50812 58215
rect 50774 58163 50777 58198
rect 50720 58152 50777 58163
rect 50823 58152 50880 58198
rect 50926 58152 50983 58198
rect 51029 58152 51086 58198
rect 51132 58152 51189 58198
rect 51235 58152 51292 58198
rect 51338 58152 51395 58198
rect 51441 58152 51454 58198
rect 50262 58123 50812 58152
rect 48557 58066 48687 58107
rect 48905 58061 49877 58092
rect 48765 58015 48778 58061
rect 48824 58015 48881 58061
rect 48927 58052 48984 58061
rect 48927 58015 48943 58052
rect 49030 58015 49087 58061
rect 49133 58052 49190 58061
rect 49133 58015 49154 58052
rect 49236 58015 49293 58061
rect 49339 58052 49396 58061
rect 49339 58015 49365 58052
rect 49442 58015 49499 58061
rect 49545 58052 49602 58061
rect 49545 58015 49576 58052
rect 49852 58015 49877 58061
rect 48905 58000 48943 58015
rect 48995 58000 49154 58015
rect 49206 58000 49365 58015
rect 49417 58000 49576 58015
rect 49628 58000 49787 58015
rect 49839 58000 49877 58015
rect 44605 57928 44812 57974
rect 44858 57928 44925 57974
rect 44971 57928 45038 57974
rect 45084 57928 45151 57974
rect 45197 57928 45264 57974
rect 45310 57928 45323 57974
rect 48905 57960 49877 58000
rect 51035 57977 51343 58017
rect 51035 57974 51073 57977
rect 51125 57974 51253 57977
rect 51305 57974 51343 57977
rect 43362 57891 43524 57898
rect 43362 57845 43373 57891
rect 43513 57845 43524 57891
rect 43362 57834 43524 57845
rect 45584 57914 48546 57950
rect 50454 57928 50467 57974
rect 50513 57928 50571 57974
rect 50617 57928 50674 57974
rect 50720 57928 50777 57974
rect 50823 57928 50880 57974
rect 50926 57928 50983 57974
rect 51029 57928 51073 57974
rect 51132 57928 51189 57974
rect 51235 57928 51253 57974
rect 51338 57928 51395 57974
rect 51441 57928 51454 57974
rect 45584 57868 45619 57914
rect 45665 57868 45777 57914
rect 45823 57868 45935 57914
rect 45981 57868 46093 57914
rect 46139 57868 46251 57914
rect 46297 57868 46409 57914
rect 46455 57868 46568 57914
rect 46614 57868 46726 57914
rect 46772 57868 46884 57914
rect 46930 57868 47042 57914
rect 47088 57868 47200 57914
rect 47246 57868 47358 57914
rect 47404 57868 47516 57914
rect 47562 57868 47675 57914
rect 47721 57868 47833 57914
rect 47879 57868 47991 57914
rect 48037 57868 48149 57914
rect 48195 57868 48307 57914
rect 48353 57868 48465 57914
rect 48511 57868 48546 57914
rect 51035 57925 51073 57928
rect 51125 57925 51253 57928
rect 51305 57925 51343 57928
rect 51035 57884 51343 57925
rect 51589 57900 51600 58322
rect 51646 57900 51657 58322
rect 54085 58323 54540 58441
rect 54085 58277 54440 58323
rect 54486 58277 54540 58323
rect 54085 58249 54540 58277
rect 53585 58198 54540 58249
rect 51789 58152 51802 58198
rect 53776 58160 54540 58198
rect 53776 58152 54440 58160
rect 53585 58130 54440 58152
rect 54085 58114 54440 58130
rect 54486 58114 54540 58160
rect 54085 58038 54540 58114
rect 51797 57984 52105 58024
rect 51797 57974 51835 57984
rect 51887 57974 52015 57984
rect 52067 57974 52105 57984
rect 54085 57992 54223 58038
rect 54269 57997 54540 58038
rect 54269 57992 54440 57997
rect 51789 57928 51802 57974
rect 53776 57928 53789 57974
rect 54085 57951 54440 57992
rect 54486 57951 54540 57997
rect 51589 57889 51657 57900
rect 51797 57891 52105 57928
rect 40215 57787 40523 57794
rect 40788 57787 42986 57801
rect 43753 57787 44514 57794
rect 39492 57764 42986 57787
rect 43704 57764 44514 57787
rect 39492 57753 44514 57764
rect 39492 57750 40253 57753
rect 39492 57704 39740 57750
rect 39786 57704 39862 57750
rect 39908 57704 39985 57750
rect 40031 57704 40108 57750
rect 40154 57704 40253 57750
rect 39492 57701 40253 57704
rect 40305 57701 40433 57753
rect 40485 57750 43790 57753
rect 40485 57704 40836 57750
rect 40882 57704 40994 57750
rect 41040 57704 41152 57750
rect 41198 57704 41310 57750
rect 41356 57704 41469 57750
rect 41515 57704 41627 57750
rect 41673 57704 41785 57750
rect 41831 57704 41943 57750
rect 41989 57704 42101 57750
rect 42147 57704 42259 57750
rect 42305 57704 42418 57750
rect 42464 57704 42576 57750
rect 42622 57704 42734 57750
rect 42780 57704 42892 57750
rect 42938 57704 43739 57750
rect 43785 57704 43790 57750
rect 40485 57701 43790 57704
rect 43842 57750 44001 57753
rect 43842 57704 43906 57750
rect 43952 57704 44001 57750
rect 43842 57701 44001 57704
rect 44053 57750 44213 57753
rect 44265 57750 44424 57753
rect 44053 57704 44071 57750
rect 44117 57704 44213 57750
rect 44282 57704 44424 57750
rect 44053 57701 44213 57704
rect 44265 57701 44424 57704
rect 44476 57701 44514 57753
rect 39492 57690 44514 57701
rect 39492 57667 42986 57690
rect 43704 57667 44514 57690
rect 39492 57215 39608 57667
rect 40215 57660 40523 57667
rect 40788 57653 42986 57667
rect 43753 57660 44514 57667
rect 44796 57787 45346 57794
rect 45584 57787 48546 57868
rect 54085 57874 54540 57951
rect 54085 57828 54223 57874
rect 54269 57834 54540 57874
rect 54269 57828 54440 57834
rect 54085 57794 54440 57828
rect 48800 57787 49982 57794
rect 50308 57787 50859 57794
rect 44796 57753 49982 57787
rect 44796 57750 44834 57753
rect 44886 57750 45045 57753
rect 45097 57750 45256 57753
rect 45308 57750 48838 57753
rect 44796 57704 44812 57750
rect 44886 57704 44925 57750
rect 44971 57704 45038 57750
rect 45097 57704 45151 57750
rect 45197 57704 45256 57750
rect 45310 57704 45619 57750
rect 45665 57704 45777 57750
rect 45823 57704 45935 57750
rect 45981 57704 46093 57750
rect 46139 57704 46251 57750
rect 46297 57704 46409 57750
rect 46455 57704 46568 57750
rect 46614 57704 46726 57750
rect 46772 57704 46884 57750
rect 46930 57704 47042 57750
rect 47088 57704 47200 57750
rect 47246 57704 47358 57750
rect 47404 57704 47516 57750
rect 47562 57704 47675 57750
rect 47721 57704 47833 57750
rect 47879 57704 47991 57750
rect 48037 57704 48149 57750
rect 48195 57704 48307 57750
rect 48353 57704 48465 57750
rect 48511 57704 48838 57750
rect 44796 57701 44834 57704
rect 44886 57701 45045 57704
rect 45097 57701 45256 57704
rect 45308 57701 48838 57704
rect 48890 57701 49048 57753
rect 49100 57701 49259 57753
rect 49311 57701 49471 57753
rect 49523 57701 49682 57753
rect 49734 57701 49892 57753
rect 49944 57701 49982 57753
rect 44796 57667 49982 57701
rect 50307 57753 50859 57787
rect 50307 57701 50346 57753
rect 50398 57750 50557 57753
rect 50609 57750 50768 57753
rect 50820 57750 50859 57753
rect 52278 57788 54440 57794
rect 54486 57788 54540 57834
rect 55927 58487 57736 58601
rect 55927 58444 56267 58487
rect 55927 58398 55961 58444
rect 56007 58441 56267 58444
rect 56313 58441 57736 58487
rect 56007 58398 57736 58441
rect 55927 58323 57736 58398
rect 55927 58281 56267 58323
rect 55927 58235 55961 58281
rect 56007 58277 56267 58281
rect 56313 58277 57736 58323
rect 56007 58235 57736 58277
rect 55927 58160 57736 58235
rect 55927 58117 56267 58160
rect 55927 58071 55961 58117
rect 56007 58114 56267 58117
rect 56313 58114 57736 58160
rect 56007 58071 57736 58114
rect 55927 57997 57736 58071
rect 55927 57954 56267 57997
rect 55927 57908 55961 57954
rect 56007 57951 56267 57954
rect 56313 57951 57736 57997
rect 56007 57908 57736 57951
rect 55927 57834 57736 57908
rect 52278 57753 54540 57788
rect 52278 57750 52316 57753
rect 52368 57750 52527 57753
rect 52579 57750 52738 57753
rect 52790 57750 52948 57753
rect 53000 57750 53159 57753
rect 53211 57750 53371 57753
rect 53423 57750 53582 57753
rect 53634 57750 53792 57753
rect 50398 57704 50467 57750
rect 50513 57704 50557 57750
rect 50617 57704 50674 57750
rect 50720 57704 50768 57750
rect 50823 57704 50880 57750
rect 50926 57704 50983 57750
rect 51029 57704 51086 57750
rect 51132 57704 51189 57750
rect 51235 57704 51292 57750
rect 51338 57704 51395 57750
rect 51441 57704 51454 57750
rect 51789 57704 51802 57750
rect 53776 57704 53792 57750
rect 50398 57701 50557 57704
rect 50609 57701 50768 57704
rect 50820 57701 50859 57704
rect 50307 57667 50859 57701
rect 44796 57660 45346 57667
rect 43362 57609 43524 57620
rect 39737 57526 39866 57555
rect 40246 57537 40362 57574
rect 43362 57563 43373 57609
rect 43513 57563 43524 57609
rect 43362 57556 43524 57563
rect 39727 57480 39740 57526
rect 39786 57515 39862 57526
rect 39827 57480 39862 57515
rect 39908 57480 39985 57526
rect 40031 57480 40108 57526
rect 40154 57480 40167 57526
rect 40246 57491 40281 57537
rect 40327 57491 40362 57537
rect 39737 57463 39775 57480
rect 39827 57463 39866 57480
rect 39737 57436 39866 57463
rect 39737 57423 39865 57436
rect 39923 57300 40085 57340
rect 39923 57248 39994 57300
rect 40046 57248 40085 57300
rect 39008 57169 39021 57215
rect 39067 57169 39144 57215
rect 39190 57169 39267 57215
rect 39313 57169 39326 57215
rect 39492 57169 39641 57215
rect 39687 57169 39730 57215
rect 39014 57137 39323 57169
rect 39492 57137 39608 57169
rect 37853 57025 38161 57030
rect 36438 56991 36953 57025
rect 37439 56991 38161 57025
rect 38658 57005 38726 57127
rect 39923 57117 40085 57248
rect 39809 57114 40085 57117
rect 39809 57106 39994 57114
rect 39809 57060 39844 57106
rect 39890 57062 39994 57106
rect 40046 57093 40085 57114
rect 40246 57093 40362 57491
rect 40718 57515 43524 57556
rect 45584 57586 48546 57667
rect 48800 57660 49982 57667
rect 50308 57660 50859 57667
rect 52278 57701 52316 57704
rect 52368 57701 52527 57704
rect 52579 57701 52738 57704
rect 52790 57701 52948 57704
rect 53000 57701 53159 57704
rect 53211 57701 53371 57704
rect 53423 57701 53582 57704
rect 53634 57701 53792 57704
rect 53844 57701 54003 57753
rect 54055 57701 54214 57753
rect 54266 57701 54540 57753
rect 52278 57666 54540 57701
rect 52278 57660 54440 57666
rect 45584 57540 45619 57586
rect 45665 57540 45777 57586
rect 45823 57540 45935 57586
rect 45981 57540 46093 57586
rect 46139 57540 46251 57586
rect 46297 57540 46409 57586
rect 46455 57540 46568 57586
rect 46614 57540 46726 57586
rect 46772 57540 46884 57586
rect 46930 57540 47042 57586
rect 47088 57540 47200 57586
rect 47246 57540 47358 57586
rect 47404 57540 47516 57586
rect 47562 57540 47675 57586
rect 47721 57540 47833 57586
rect 47879 57540 47991 57586
rect 48037 57540 48149 57586
rect 48195 57540 48307 57586
rect 48353 57540 48465 57586
rect 48511 57540 48546 57586
rect 54085 57626 54440 57660
rect 54085 57580 54223 57626
rect 54269 57620 54440 57626
rect 54486 57620 54540 57666
rect 54758 57753 55840 57794
rect 54758 57750 54855 57753
rect 54758 57704 54793 57750
rect 54839 57704 54855 57750
rect 54758 57701 54855 57704
rect 54907 57750 55066 57753
rect 54907 57704 54956 57750
rect 55002 57704 55066 57750
rect 54907 57701 55066 57704
rect 55118 57750 55278 57753
rect 55330 57750 55489 57753
rect 55164 57704 55278 57750
rect 55330 57704 55439 57750
rect 55485 57704 55489 57750
rect 55118 57701 55278 57704
rect 55330 57701 55489 57704
rect 55541 57750 55840 57753
rect 55541 57704 55599 57750
rect 55645 57704 55760 57750
rect 55806 57704 55840 57750
rect 55541 57701 55840 57704
rect 54758 57661 55840 57701
rect 55927 57788 56267 57834
rect 56313 57788 57736 57834
rect 55927 57666 57736 57788
rect 54817 57660 55579 57661
rect 54269 57580 54540 57620
rect 40718 57463 41935 57515
rect 41987 57463 43524 57515
rect 40718 57422 43524 57463
rect 44605 57480 44812 57526
rect 44858 57480 44925 57526
rect 44971 57480 45038 57526
rect 45084 57480 45151 57526
rect 45197 57480 45264 57526
rect 45310 57480 45323 57526
rect 45584 57504 48546 57540
rect 51035 57529 51343 57570
rect 51035 57526 51073 57529
rect 51125 57526 51253 57529
rect 51305 57526 51343 57529
rect 51589 57554 51657 57565
rect 44341 57414 44509 57425
rect 44341 57368 44358 57414
rect 44498 57368 44509 57414
rect 44341 57324 44509 57368
rect 42229 57284 44509 57324
rect 42229 57232 42690 57284
rect 42742 57232 44509 57284
rect 42229 57191 44509 57232
rect 44605 57093 44721 57480
rect 48905 57454 49877 57494
rect 50454 57480 50467 57526
rect 50513 57480 50571 57526
rect 50617 57480 50674 57526
rect 50720 57480 50777 57526
rect 50823 57480 50880 57526
rect 50926 57480 50983 57526
rect 51029 57480 51073 57526
rect 51132 57480 51189 57526
rect 51235 57480 51253 57526
rect 51338 57480 51395 57526
rect 51441 57480 51454 57526
rect 48905 57439 48943 57454
rect 48995 57439 49154 57454
rect 49206 57439 49365 57454
rect 49417 57439 49576 57454
rect 49628 57439 49787 57454
rect 49839 57439 49877 57454
rect 48765 57393 48778 57439
rect 48824 57393 48881 57439
rect 48927 57402 48943 57439
rect 48927 57393 48984 57402
rect 49030 57393 49087 57439
rect 49133 57402 49154 57439
rect 49133 57393 49190 57402
rect 49236 57393 49293 57439
rect 49339 57402 49365 57439
rect 49339 57393 49396 57402
rect 49442 57393 49499 57439
rect 49545 57402 49576 57439
rect 49545 57393 49602 57402
rect 49852 57393 49877 57439
rect 51035 57477 51073 57480
rect 51125 57477 51253 57480
rect 51305 57477 51343 57480
rect 51035 57437 51343 57477
rect 48557 57347 48687 57388
rect 48905 57362 49877 57393
rect 44901 57302 45241 57331
rect 44799 57256 44812 57302
rect 44858 57256 44925 57302
rect 44971 57291 45038 57302
rect 44991 57256 45038 57291
rect 45084 57256 45151 57302
rect 45197 57291 45264 57302
rect 45203 57256 45264 57291
rect 45310 57256 45323 57302
rect 48557 57295 48596 57347
rect 48648 57295 48687 57347
rect 48557 57292 48687 57295
rect 44901 57239 44939 57256
rect 44991 57239 45151 57256
rect 45203 57239 45241 57256
rect 44901 57198 45241 57239
rect 45400 57183 48379 57216
rect 45400 57137 45464 57183
rect 45604 57175 48379 57183
rect 45400 57123 45597 57137
rect 45649 57123 48379 57175
rect 40046 57078 44918 57093
rect 45400 57082 48379 57123
rect 48557 57152 48622 57292
rect 48668 57152 48687 57292
rect 50262 57302 50812 57331
rect 50262 57291 50467 57302
rect 50513 57291 50571 57302
rect 49820 57215 50160 57256
rect 48765 57169 48778 57215
rect 48824 57169 48881 57215
rect 48927 57169 48984 57215
rect 49030 57169 49087 57215
rect 49133 57169 49190 57215
rect 49236 57169 49293 57215
rect 49339 57169 49396 57215
rect 49442 57169 49499 57215
rect 49545 57169 49602 57215
rect 49852 57169 50160 57215
rect 50262 57239 50300 57291
rect 50352 57256 50467 57291
rect 50563 57256 50571 57291
rect 50617 57256 50674 57302
rect 50720 57291 50777 57302
rect 50720 57256 50722 57291
rect 50352 57239 50511 57256
rect 50563 57239 50722 57256
rect 50774 57256 50777 57291
rect 50823 57256 50880 57302
rect 50926 57256 50983 57302
rect 51029 57256 51086 57302
rect 51132 57256 51189 57302
rect 51235 57256 51292 57302
rect 51338 57256 51395 57302
rect 51441 57256 51454 57302
rect 50774 57239 50812 57256
rect 50262 57198 50812 57239
rect 48557 57129 48687 57152
rect 49820 57137 50160 57169
rect 40046 57062 44812 57078
rect 39890 57060 44812 57062
rect 39809 57057 44812 57060
rect 39809 57011 43739 57057
rect 43785 57011 43906 57057
rect 43952 57011 44071 57057
rect 44117 57011 44236 57057
rect 44282 57032 44812 57057
rect 44858 57032 44925 57078
rect 44971 57032 45038 57078
rect 45084 57032 45151 57078
rect 45197 57032 45264 57078
rect 45310 57032 45323 57078
rect 48557 57077 48596 57129
rect 48648 57077 48687 57129
rect 48557 57037 48687 57077
rect 50044 57080 50160 57137
rect 51589 57132 51600 57554
rect 51646 57132 51657 57554
rect 51797 57526 52105 57563
rect 51789 57480 51802 57526
rect 53776 57480 53789 57526
rect 54085 57503 54540 57580
rect 51797 57470 51835 57480
rect 51887 57470 52015 57480
rect 52067 57470 52105 57480
rect 51797 57430 52105 57470
rect 54085 57462 54440 57503
rect 54085 57416 54223 57462
rect 54269 57457 54440 57462
rect 54486 57457 54540 57503
rect 54269 57416 54540 57457
rect 54085 57340 54540 57416
rect 54085 57324 54440 57340
rect 53585 57302 54440 57324
rect 51789 57256 51802 57302
rect 53776 57294 54440 57302
rect 54486 57294 54540 57340
rect 53776 57256 54540 57294
rect 53585 57205 54540 57256
rect 51589 57080 51657 57132
rect 54085 57177 54540 57205
rect 54085 57131 54440 57177
rect 54486 57131 54540 57177
rect 50044 57043 51657 57080
rect 51797 57078 52105 57100
rect 44282 57011 44918 57032
rect 38658 56991 39723 57005
rect 30683 56967 30855 56973
rect 30583 56927 30855 56967
rect 30901 56927 31040 56973
rect 33484 56960 34643 56989
rect 35260 56945 35273 56991
rect 35523 56945 35543 56991
rect 35626 56945 35683 56991
rect 35729 56945 35754 56991
rect 35832 56945 35889 56991
rect 35935 56945 35965 56991
rect 36038 56945 36095 56991
rect 36141 56945 36176 56991
rect 36244 56945 36301 56991
rect 36347 56945 36360 56991
rect 36438 56945 36854 56991
rect 36900 56945 36971 56991
rect 37017 56945 37088 56991
rect 37134 56945 37206 56991
rect 37252 56945 37324 56991
rect 37370 56945 37442 56991
rect 37488 56989 37909 56991
rect 37488 56945 37891 56989
rect 37955 56945 38026 56991
rect 38072 56989 38143 56991
rect 38123 56945 38143 56989
rect 38189 56945 38261 56991
rect 38307 56945 38379 56991
rect 38425 56945 38497 56991
rect 38543 56945 38556 56991
rect 38658 56945 39021 56991
rect 39067 56945 39144 56991
rect 39190 56945 39267 56991
rect 39313 56945 39641 56991
rect 39687 56945 39730 56991
rect 39809 56973 44918 57011
rect 48905 56991 49877 57031
rect 48765 56945 48778 56991
rect 48824 56945 48881 56991
rect 48927 56945 48943 56991
rect 49030 56945 49087 56991
rect 49133 56945 49154 56991
rect 49236 56945 49293 56991
rect 49339 56945 49365 56991
rect 49442 56945 49499 56991
rect 49545 56945 49576 56991
rect 49852 56945 49877 56991
rect 50044 56997 50516 57043
rect 50562 56997 50703 57043
rect 50749 56997 50890 57043
rect 50936 56997 51076 57043
rect 51122 56997 51263 57043
rect 51309 56997 51657 57043
rect 51789 57032 51802 57078
rect 53776 57032 53789 57078
rect 50044 56987 51657 56997
rect 50481 56960 51657 56987
rect 51797 57007 51835 57032
rect 51887 57007 52015 57032
rect 52067 57007 52105 57032
rect 51797 56967 52105 57007
rect 54085 57013 54540 57131
rect 54085 56973 54440 57013
rect 30583 56894 31040 56927
rect 35294 56939 35332 56945
rect 35384 56939 35543 56945
rect 35595 56939 35754 56945
rect 35806 56939 35965 56945
rect 36017 56939 36176 56945
rect 36228 56939 36266 56945
rect 34870 56894 35025 56901
rect 35294 56899 36266 56939
rect 36438 56905 36953 56945
rect 37439 56937 37891 56945
rect 37943 56937 38071 56945
rect 38123 56937 38161 56945
rect 37439 56905 38161 56937
rect 37853 56897 38161 56905
rect 27387 56801 27790 56853
rect 27842 56801 28001 56853
rect 28053 56801 28212 56853
rect 28264 56801 28423 56853
rect 28475 56801 28634 56853
rect 28686 56850 28845 56853
rect 28686 56804 28810 56850
rect 28686 56801 28845 56804
rect 28897 56801 29056 56853
rect 29108 56801 29196 56853
rect 27387 56687 29196 56801
rect 29283 56853 30365 56894
rect 29283 56850 29582 56853
rect 29283 56804 29317 56850
rect 29363 56804 29478 56850
rect 29524 56804 29582 56850
rect 29283 56801 29582 56804
rect 29634 56850 29793 56853
rect 29845 56850 30005 56853
rect 29634 56804 29638 56850
rect 29684 56804 29793 56850
rect 29845 56804 29959 56850
rect 29634 56801 29793 56804
rect 29845 56801 30005 56804
rect 30057 56850 30216 56853
rect 30057 56804 30121 56850
rect 30167 56804 30216 56850
rect 30057 56801 30216 56804
rect 30268 56850 30365 56853
rect 30268 56804 30284 56850
rect 30330 56804 30365 56850
rect 30268 56801 30365 56804
rect 29283 56761 30365 56801
rect 30583 56853 32842 56894
rect 30583 56850 30854 56853
rect 30583 56804 30637 56850
rect 30683 56804 30854 56850
rect 30583 56801 30854 56804
rect 30906 56801 31065 56853
rect 31117 56801 31276 56853
rect 31328 56801 31486 56853
rect 31538 56801 31697 56853
rect 31749 56801 31909 56853
rect 31961 56801 32120 56853
rect 32172 56801 32330 56853
rect 32382 56801 32541 56853
rect 32593 56801 32752 56853
rect 32804 56801 32842 56853
rect 29544 56760 30306 56761
rect 30583 56760 32842 56801
rect 34717 56853 35025 56894
rect 38658 56885 39723 56945
rect 48905 56939 48943 56945
rect 48995 56939 49154 56945
rect 49206 56939 49365 56945
rect 49417 56939 49576 56945
rect 49628 56939 49787 56945
rect 49839 56939 49877 56945
rect 48905 56899 49877 56939
rect 54085 56927 54223 56973
rect 54269 56967 54440 56973
rect 54486 56967 54540 57013
rect 54269 56927 54540 56967
rect 50099 56894 50255 56901
rect 54085 56894 54540 56927
rect 55927 57620 56267 57666
rect 56313 57620 57736 57666
rect 55927 57544 57736 57620
rect 55927 57498 55961 57544
rect 56007 57503 57736 57544
rect 56007 57498 56267 57503
rect 55927 57457 56267 57498
rect 56313 57457 57736 57503
rect 55927 57381 57736 57457
rect 55927 57335 55961 57381
rect 56007 57340 57736 57381
rect 56007 57335 56267 57340
rect 55927 57294 56267 57335
rect 56313 57294 57736 57340
rect 55927 57217 57736 57294
rect 55927 57171 55961 57217
rect 56007 57177 57736 57217
rect 56007 57171 56267 57177
rect 55927 57131 56267 57171
rect 56313 57131 57736 57177
rect 55927 57054 57736 57131
rect 55927 57008 55961 57054
rect 56007 57013 57736 57054
rect 56007 57008 56267 57013
rect 55927 56967 56267 57008
rect 56313 56967 57736 57013
rect 34717 56801 34755 56853
rect 34807 56850 34935 56853
rect 34807 56804 34916 56850
rect 34807 56801 34935 56804
rect 34987 56801 35025 56853
rect 34717 56760 35025 56801
rect 50099 56853 50408 56894
rect 50099 56801 50138 56853
rect 50190 56850 50318 56853
rect 50206 56804 50318 56850
rect 50190 56801 50318 56804
rect 50370 56801 50408 56853
rect 27387 56641 28810 56687
rect 28856 56644 29196 56687
rect 28856 56641 29116 56644
rect 27387 56598 29116 56641
rect 29162 56598 29196 56644
rect 27387 56523 29196 56598
rect 27387 56477 28810 56523
rect 28856 56481 29196 56523
rect 28856 56477 29116 56481
rect 27387 56435 29116 56477
rect 29162 56435 29196 56481
rect 27387 56360 29196 56435
rect 27387 56314 28810 56360
rect 28856 56317 29196 56360
rect 28856 56314 29116 56317
rect 27387 56271 29116 56314
rect 29162 56271 29196 56317
rect 27387 56197 29196 56271
rect 27387 56151 28810 56197
rect 28856 56154 29196 56197
rect 28856 56151 29116 56154
rect 27387 56108 29116 56151
rect 29162 56108 29196 56154
rect 27387 56034 29196 56108
rect 27387 55988 28810 56034
rect 28856 55988 29196 56034
rect 30583 56727 31040 56760
rect 34870 56753 35025 56760
rect 30583 56687 30855 56727
rect 30583 56641 30637 56687
rect 30683 56681 30855 56687
rect 30901 56681 31040 56727
rect 35294 56715 36266 56755
rect 37853 56749 38161 56757
rect 35294 56709 35332 56715
rect 35384 56709 35543 56715
rect 35595 56709 35754 56715
rect 35806 56709 35965 56715
rect 36017 56709 36176 56715
rect 36228 56709 36266 56715
rect 36438 56709 36953 56749
rect 37439 56717 38161 56749
rect 37439 56709 37891 56717
rect 37943 56709 38071 56717
rect 38123 56709 38161 56717
rect 38658 56709 39723 56769
rect 50099 56760 50408 56801
rect 52278 56853 54540 56894
rect 52278 56801 52316 56853
rect 52368 56801 52527 56853
rect 52579 56801 52738 56853
rect 52790 56801 52948 56853
rect 53000 56801 53159 56853
rect 53211 56801 53371 56853
rect 53423 56801 53582 56853
rect 53634 56801 53792 56853
rect 53844 56801 54003 56853
rect 54055 56801 54214 56853
rect 54266 56850 54540 56853
rect 54266 56804 54440 56850
rect 54486 56804 54540 56850
rect 54266 56801 54540 56804
rect 52278 56760 54540 56801
rect 54758 56853 55840 56894
rect 54758 56850 54855 56853
rect 54758 56804 54793 56850
rect 54839 56804 54855 56850
rect 54758 56801 54855 56804
rect 54907 56850 55066 56853
rect 54907 56804 54956 56850
rect 55002 56804 55066 56850
rect 54907 56801 55066 56804
rect 55118 56850 55278 56853
rect 55330 56850 55489 56853
rect 55164 56804 55278 56850
rect 55330 56804 55439 56850
rect 55485 56804 55489 56850
rect 55118 56801 55278 56804
rect 55330 56801 55489 56804
rect 55541 56850 55840 56853
rect 55541 56804 55599 56850
rect 55645 56804 55760 56850
rect 55806 56804 55840 56850
rect 55541 56801 55840 56804
rect 54758 56761 55840 56801
rect 55927 56853 57736 56967
rect 55927 56801 56015 56853
rect 56067 56801 56226 56853
rect 56278 56850 56437 56853
rect 56313 56804 56437 56850
rect 56278 56801 56437 56804
rect 56489 56801 56648 56853
rect 56700 56801 56859 56853
rect 56911 56801 57070 56853
rect 57122 56801 57281 56853
rect 57333 56801 57736 56853
rect 54817 56760 55579 56761
rect 48905 56715 49877 56755
rect 50099 56753 50255 56760
rect 48905 56709 48943 56715
rect 48995 56709 49154 56715
rect 49206 56709 49365 56715
rect 49417 56709 49576 56715
rect 49628 56709 49787 56715
rect 49839 56709 49877 56715
rect 30683 56641 31040 56681
rect 33484 56665 34643 56694
rect 30583 56564 31040 56641
rect 33019 56625 33327 56665
rect 33019 56622 33057 56625
rect 33109 56622 33237 56625
rect 33289 56622 33327 56625
rect 33484 56657 35082 56665
rect 35260 56663 35273 56709
rect 35523 56663 35543 56709
rect 35626 56663 35683 56709
rect 35729 56663 35754 56709
rect 35832 56663 35889 56709
rect 35935 56663 35965 56709
rect 36038 56663 36095 56709
rect 36141 56663 36176 56709
rect 36244 56663 36301 56709
rect 36347 56663 36360 56709
rect 36438 56663 36854 56709
rect 36900 56663 36971 56709
rect 37017 56663 37088 56709
rect 37134 56663 37206 56709
rect 37252 56663 37324 56709
rect 37370 56663 37442 56709
rect 37488 56665 37891 56709
rect 37488 56663 37909 56665
rect 37955 56663 38026 56709
rect 38123 56665 38143 56709
rect 38072 56663 38143 56665
rect 38189 56663 38261 56709
rect 38307 56663 38379 56709
rect 38425 56663 38497 56709
rect 38543 56663 38556 56709
rect 38658 56663 39021 56709
rect 39067 56663 39144 56709
rect 39190 56663 39267 56709
rect 39313 56663 39641 56709
rect 39687 56663 39730 56709
rect 31336 56576 31349 56622
rect 33323 56576 33336 56622
rect 33484 56611 33816 56657
rect 33862 56611 34002 56657
rect 34048 56611 34189 56657
rect 34235 56611 34376 56657
rect 34422 56611 34562 56657
rect 34608 56611 35082 56657
rect 35294 56623 36266 56663
rect 36438 56629 36953 56663
rect 37439 56629 38161 56663
rect 30583 56523 30855 56564
rect 30583 56477 30637 56523
rect 30683 56518 30855 56523
rect 30901 56518 31040 56564
rect 33019 56573 33057 56576
rect 33109 56573 33237 56576
rect 33289 56573 33327 56576
rect 33019 56532 33327 56573
rect 33484 56574 35082 56611
rect 30683 56477 31040 56518
rect 30583 56449 31040 56477
rect 33484 56492 33552 56574
rect 30583 56401 31493 56449
rect 30583 56360 30855 56401
rect 30583 56314 30637 56360
rect 30683 56355 30855 56360
rect 30901 56398 31493 56401
rect 30901 56355 31349 56398
rect 30683 56352 31349 56355
rect 33323 56352 33336 56398
rect 30683 56330 31493 56352
rect 30683 56314 31040 56330
rect 30583 56238 31040 56314
rect 30583 56197 30855 56238
rect 30583 56151 30637 56197
rect 30683 56192 30855 56197
rect 30901 56192 31040 56238
rect 30683 56151 31040 56192
rect 33019 56177 33327 56217
rect 33019 56174 33057 56177
rect 33109 56174 33237 56177
rect 33289 56174 33327 56177
rect 30583 56074 31040 56151
rect 31336 56128 31349 56174
rect 33323 56128 33336 56174
rect 33019 56125 33057 56128
rect 33109 56125 33237 56128
rect 33289 56125 33327 56128
rect 33019 56084 33327 56125
rect 30583 56034 30855 56074
rect 27387 55866 29196 55988
rect 27387 55820 28810 55866
rect 28856 55820 29196 55866
rect 29283 55953 30365 55994
rect 29283 55950 29582 55953
rect 29283 55904 29317 55950
rect 29363 55904 29478 55950
rect 29524 55904 29582 55950
rect 29283 55901 29582 55904
rect 29634 55950 29793 55953
rect 29845 55950 30005 55953
rect 29634 55904 29638 55950
rect 29684 55904 29793 55950
rect 29845 55904 29959 55950
rect 29634 55901 29793 55904
rect 29845 55901 30005 55904
rect 30057 55950 30216 55953
rect 30057 55904 30121 55950
rect 30167 55904 30216 55950
rect 30057 55901 30216 55904
rect 30268 55950 30365 55953
rect 30268 55904 30284 55950
rect 30330 55904 30365 55950
rect 30268 55901 30365 55904
rect 29283 55861 30365 55901
rect 30583 55988 30637 56034
rect 30683 56028 30855 56034
rect 30901 56028 31040 56074
rect 33484 56070 33495 56492
rect 33541 56070 33552 56492
rect 34964 56517 35082 56574
rect 36438 56529 36554 56629
rect 37853 56624 38161 56629
rect 38658 56649 39723 56663
rect 34964 56485 36360 56517
rect 34228 56415 34718 56456
rect 34228 56398 34267 56415
rect 34319 56398 34447 56415
rect 34499 56398 34627 56415
rect 33671 56352 33684 56398
rect 33730 56352 33787 56398
rect 33833 56352 33890 56398
rect 33936 56352 33993 56398
rect 34039 56352 34096 56398
rect 34142 56352 34199 56398
rect 34245 56363 34267 56398
rect 34245 56352 34302 56363
rect 34348 56352 34405 56398
rect 34499 56363 34508 56398
rect 34451 56352 34508 56363
rect 34554 56352 34612 56398
rect 34679 56363 34718 56415
rect 34964 56439 35273 56485
rect 35523 56439 35580 56485
rect 35626 56439 35683 56485
rect 35729 56439 35786 56485
rect 35832 56439 35889 56485
rect 35935 56439 35992 56485
rect 36038 56439 36095 56485
rect 36141 56439 36198 56485
rect 36244 56439 36301 56485
rect 36347 56439 36360 56485
rect 34964 56395 36360 56439
rect 34658 56352 34718 56363
rect 34228 56323 34718 56352
rect 36438 56389 36475 56529
rect 36521 56389 36554 56529
rect 35294 56261 36266 56295
rect 36438 56286 36554 56389
rect 36640 56529 36773 56549
rect 36640 56490 36697 56529
rect 36640 56438 36678 56490
rect 36640 56389 36697 56438
rect 36743 56389 36773 56529
rect 38658 56527 38726 56649
rect 39809 56643 44918 56681
rect 48765 56663 48778 56709
rect 48824 56663 48881 56709
rect 48927 56663 48943 56709
rect 49030 56663 49087 56709
rect 49133 56663 49154 56709
rect 49236 56663 49293 56709
rect 49339 56663 49365 56709
rect 49442 56663 49499 56709
rect 49545 56663 49576 56709
rect 49852 56663 49877 56709
rect 54085 56727 54540 56760
rect 50481 56667 51657 56694
rect 39809 56597 43739 56643
rect 43785 56597 43906 56643
rect 43952 56597 44071 56643
rect 44117 56597 44236 56643
rect 44282 56622 44918 56643
rect 48905 56623 49877 56663
rect 50044 56657 51657 56667
rect 44282 56597 44812 56622
rect 39809 56594 44812 56597
rect 39809 56548 39844 56594
rect 39890 56592 44812 56594
rect 39890 56548 39994 56592
rect 39809 56540 39994 56548
rect 40046 56576 44812 56592
rect 44858 56576 44925 56622
rect 44971 56576 45038 56622
rect 45084 56576 45151 56622
rect 45197 56576 45264 56622
rect 45310 56576 45323 56622
rect 48557 56577 48687 56617
rect 40046 56561 44918 56576
rect 40046 56540 40085 56561
rect 39809 56537 40085 56540
rect 36924 56517 37685 56524
rect 36923 56485 37931 56517
rect 36841 56439 36854 56485
rect 36900 56483 36971 56485
rect 36900 56439 36961 56483
rect 37017 56439 37088 56485
rect 37134 56483 37206 56485
rect 37134 56439 37172 56483
rect 37252 56439 37324 56485
rect 37370 56483 37442 56485
rect 37370 56439 37384 56483
rect 36923 56431 36961 56439
rect 37013 56431 37172 56439
rect 37224 56431 37384 56439
rect 37436 56439 37442 56483
rect 37488 56483 37909 56485
rect 37488 56439 37595 56483
rect 37436 56431 37595 56439
rect 37647 56439 37909 56483
rect 37955 56439 38026 56485
rect 38072 56439 38143 56485
rect 38189 56439 38261 56485
rect 38307 56439 38379 56485
rect 38425 56439 38497 56485
rect 38543 56439 38556 56485
rect 37647 56431 37931 56439
rect 36923 56398 37931 56431
rect 36923 56397 37685 56398
rect 36924 56391 37685 56397
rect 36640 56366 36773 56389
rect 38658 56387 38669 56527
rect 38715 56387 38726 56527
rect 39014 56485 39323 56517
rect 39492 56485 39608 56517
rect 39008 56439 39021 56485
rect 39067 56439 39144 56485
rect 39190 56439 39267 56485
rect 39313 56439 39326 56485
rect 39492 56439 39641 56485
rect 39687 56439 39730 56485
rect 38658 56376 38726 56387
rect 36438 56261 36953 56286
rect 37439 56283 37931 56286
rect 37439 56261 38161 56283
rect 35260 56215 35273 56261
rect 35523 56255 35580 56261
rect 35523 56215 35543 56255
rect 35626 56215 35683 56261
rect 35729 56255 35786 56261
rect 35729 56215 35754 56255
rect 35832 56215 35889 56261
rect 35935 56255 35992 56261
rect 35935 56215 35965 56255
rect 36038 56215 36095 56261
rect 36141 56255 36198 56261
rect 36141 56215 36176 56255
rect 36244 56215 36301 56261
rect 36347 56215 36360 56261
rect 36438 56215 36854 56261
rect 36900 56215 36971 56261
rect 37017 56215 37088 56261
rect 37134 56215 37206 56261
rect 37252 56215 37324 56261
rect 37370 56215 37442 56261
rect 37488 56243 37909 56261
rect 37488 56215 37891 56243
rect 37955 56215 38026 56261
rect 38072 56243 38143 56261
rect 38123 56215 38143 56243
rect 38189 56215 38261 56261
rect 38307 56215 38379 56261
rect 38425 56215 38497 56261
rect 38543 56215 38556 56261
rect 33781 56174 34089 56209
rect 35294 56203 35332 56215
rect 35384 56203 35543 56215
rect 35595 56203 35754 56215
rect 35806 56203 35965 56215
rect 36017 56203 36176 56215
rect 36228 56203 36266 56215
rect 33671 56128 33684 56174
rect 33730 56128 33787 56174
rect 33833 56169 33890 56174
rect 33871 56128 33890 56169
rect 33936 56128 33993 56174
rect 34039 56169 34096 56174
rect 34051 56128 34096 56169
rect 34142 56128 34199 56174
rect 34245 56128 34302 56174
rect 34348 56128 34405 56174
rect 34451 56128 34508 56174
rect 34554 56128 34612 56174
rect 34658 56128 34671 56174
rect 35294 56163 36266 56203
rect 36438 56166 36953 56215
rect 37439 56191 37891 56215
rect 37943 56191 38071 56215
rect 38123 56191 38161 56215
rect 37439 56166 38161 56191
rect 37853 56150 38161 56166
rect 33781 56117 33819 56128
rect 33871 56117 33999 56128
rect 34051 56117 34089 56128
rect 33781 56076 34089 56117
rect 33484 56059 33552 56070
rect 30683 55994 31040 56028
rect 30683 55988 32842 55994
rect 30583 55953 32842 55988
rect 34247 55987 35008 55994
rect 30583 55901 30854 55953
rect 30906 55901 31065 55953
rect 31117 55901 31276 55953
rect 31328 55950 31486 55953
rect 31538 55950 31697 55953
rect 31749 55950 31909 55953
rect 31961 55950 32120 55953
rect 32172 55950 32330 55953
rect 32382 55950 32541 55953
rect 32593 55950 32752 55953
rect 32804 55950 32842 55953
rect 34246 55953 35008 55987
rect 34246 55950 34284 55953
rect 34336 55950 34495 55953
rect 34547 55950 34707 55953
rect 31328 55904 31349 55950
rect 33323 55904 33336 55950
rect 33671 55904 33684 55950
rect 33730 55904 33787 55950
rect 33833 55904 33890 55950
rect 33936 55904 33993 55950
rect 34039 55904 34096 55950
rect 34142 55904 34199 55950
rect 34245 55904 34284 55950
rect 34348 55904 34405 55950
rect 34451 55904 34495 55950
rect 34554 55904 34612 55950
rect 34658 55904 34707 55950
rect 31328 55901 31486 55904
rect 31538 55901 31697 55904
rect 31749 55901 31909 55904
rect 31961 55901 32120 55904
rect 32172 55901 32330 55904
rect 32382 55901 32541 55904
rect 32593 55901 32752 55904
rect 32804 55901 32842 55904
rect 30583 55866 32842 55901
rect 34246 55901 34284 55904
rect 34336 55901 34495 55904
rect 34547 55901 34707 55904
rect 34759 55901 34918 55953
rect 34970 55901 35008 55953
rect 34246 55867 35008 55901
rect 29544 55860 30306 55861
rect 27387 55744 29196 55820
rect 27387 55703 29116 55744
rect 27387 55657 28810 55703
rect 28856 55698 29116 55703
rect 29162 55698 29196 55744
rect 28856 55657 29196 55698
rect 27387 55581 29196 55657
rect 27387 55540 29116 55581
rect 27387 55494 28810 55540
rect 28856 55535 29116 55540
rect 29162 55535 29196 55581
rect 28856 55494 29196 55535
rect 27387 55417 29196 55494
rect 27387 55377 29116 55417
rect 27387 55331 28810 55377
rect 28856 55371 29116 55377
rect 29162 55371 29196 55417
rect 28856 55331 29196 55371
rect 27387 55254 29196 55331
rect 27387 55213 29116 55254
rect 27387 55167 28810 55213
rect 28856 55208 29116 55213
rect 29162 55208 29196 55254
rect 28856 55167 29196 55208
rect 27387 55053 29196 55167
rect 30583 55820 30637 55866
rect 30683 55860 32842 55866
rect 34247 55860 35008 55867
rect 35182 55987 36364 55994
rect 35182 55953 36958 55987
rect 35182 55901 35220 55953
rect 35272 55901 35430 55953
rect 35482 55901 35641 55953
rect 35693 55901 35853 55953
rect 35905 55901 36064 55953
rect 36116 55901 36274 55953
rect 36326 55950 36958 55953
rect 36326 55904 36489 55950
rect 36723 55904 36958 55950
rect 36326 55901 36958 55904
rect 35182 55867 36958 55901
rect 37946 55953 38842 55994
rect 37946 55950 38330 55953
rect 38382 55950 38541 55953
rect 37946 55904 37957 55950
rect 38473 55904 38541 55950
rect 37946 55901 38330 55904
rect 38382 55901 38541 55904
rect 38593 55901 38752 55953
rect 38804 55901 38842 55953
rect 35182 55860 36364 55867
rect 37946 55860 38842 55901
rect 39014 55953 39323 56439
rect 39014 55901 39052 55953
rect 39104 55950 39232 55953
rect 39108 55904 39220 55950
rect 39104 55901 39232 55904
rect 39284 55901 39323 55953
rect 30683 55826 31040 55860
rect 30683 55820 30855 55826
rect 30583 55780 30855 55820
rect 30901 55780 31040 55826
rect 30583 55703 31040 55780
rect 33484 55784 33552 55795
rect 33019 55729 33327 55770
rect 33019 55726 33057 55729
rect 33109 55726 33237 55729
rect 33289 55726 33327 55729
rect 30583 55657 30637 55703
rect 30683 55662 31040 55703
rect 31336 55680 31349 55726
rect 33323 55680 33336 55726
rect 30683 55657 30855 55662
rect 30583 55616 30855 55657
rect 30901 55616 31040 55662
rect 33019 55677 33057 55680
rect 33109 55677 33237 55680
rect 33289 55677 33327 55680
rect 33019 55637 33327 55677
rect 30583 55540 31040 55616
rect 30583 55494 30637 55540
rect 30683 55524 31040 55540
rect 30683 55502 31493 55524
rect 30683 55499 31349 55502
rect 30683 55494 30855 55499
rect 30583 55453 30855 55494
rect 30901 55456 31349 55499
rect 33323 55456 33336 55502
rect 30901 55453 31493 55456
rect 30583 55405 31493 55453
rect 30583 55377 31040 55405
rect 30583 55331 30637 55377
rect 30683 55336 31040 55377
rect 30683 55331 30855 55336
rect 30583 55290 30855 55331
rect 30901 55290 31040 55336
rect 33484 55362 33495 55784
rect 33541 55362 33552 55784
rect 33781 55737 34089 55778
rect 33781 55726 33819 55737
rect 33871 55726 33999 55737
rect 34051 55726 34089 55737
rect 33671 55680 33684 55726
rect 33730 55680 33787 55726
rect 33871 55685 33890 55726
rect 33833 55680 33890 55685
rect 33936 55680 33993 55726
rect 34051 55685 34096 55726
rect 34039 55680 34096 55685
rect 34142 55680 34199 55726
rect 34245 55680 34302 55726
rect 34348 55680 34405 55726
rect 34451 55680 34508 55726
rect 34554 55680 34612 55726
rect 34658 55680 34671 55726
rect 33781 55645 34089 55680
rect 35294 55651 36266 55691
rect 37853 55688 38161 55704
rect 35294 55639 35332 55651
rect 35384 55639 35543 55651
rect 35595 55639 35754 55651
rect 35806 55639 35965 55651
rect 36017 55639 36176 55651
rect 36228 55639 36266 55651
rect 36438 55639 36953 55688
rect 37439 55663 38161 55688
rect 37439 55639 37891 55663
rect 37943 55639 38071 55663
rect 38123 55639 38161 55663
rect 35260 55593 35273 55639
rect 35523 55599 35543 55639
rect 35523 55593 35580 55599
rect 35626 55593 35683 55639
rect 35729 55599 35754 55639
rect 35729 55593 35786 55599
rect 35832 55593 35889 55639
rect 35935 55599 35965 55639
rect 35935 55593 35992 55599
rect 36038 55593 36095 55639
rect 36141 55599 36176 55639
rect 36141 55593 36198 55599
rect 36244 55593 36301 55639
rect 36347 55593 36360 55639
rect 36438 55593 36854 55639
rect 36900 55593 36971 55639
rect 37017 55593 37088 55639
rect 37134 55593 37206 55639
rect 37252 55593 37324 55639
rect 37370 55593 37442 55639
rect 37488 55611 37891 55639
rect 37488 55593 37909 55611
rect 37955 55593 38026 55639
rect 38123 55611 38143 55639
rect 38072 55593 38143 55611
rect 38189 55593 38261 55639
rect 38307 55593 38379 55639
rect 38425 55593 38497 55639
rect 38543 55593 38556 55639
rect 35294 55559 36266 55593
rect 36438 55568 36953 55593
rect 37439 55571 38161 55593
rect 37439 55568 37931 55571
rect 34228 55502 34718 55531
rect 33671 55456 33684 55502
rect 33730 55456 33787 55502
rect 33833 55456 33890 55502
rect 33936 55456 33993 55502
rect 34039 55456 34096 55502
rect 34142 55456 34199 55502
rect 34245 55491 34302 55502
rect 34245 55456 34267 55491
rect 34348 55456 34405 55502
rect 34451 55491 34508 55502
rect 34499 55456 34508 55491
rect 34554 55456 34612 55502
rect 34658 55491 34718 55502
rect 34228 55439 34267 55456
rect 34319 55439 34447 55456
rect 34499 55439 34627 55456
rect 34679 55439 34718 55491
rect 36438 55465 36554 55568
rect 34228 55398 34718 55439
rect 34964 55415 36360 55459
rect 30583 55213 31040 55290
rect 33019 55281 33327 55322
rect 33019 55278 33057 55281
rect 33109 55278 33237 55281
rect 33289 55278 33327 55281
rect 33484 55280 33552 55362
rect 34964 55369 35273 55415
rect 35523 55369 35580 55415
rect 35626 55369 35683 55415
rect 35729 55369 35786 55415
rect 35832 55369 35889 55415
rect 35935 55369 35992 55415
rect 36038 55369 36095 55415
rect 36141 55369 36198 55415
rect 36244 55369 36301 55415
rect 36347 55369 36360 55415
rect 34964 55337 36360 55369
rect 34964 55280 35082 55337
rect 31336 55232 31349 55278
rect 33323 55232 33336 55278
rect 33484 55243 35082 55280
rect 30583 55167 30637 55213
rect 30683 55173 31040 55213
rect 33019 55229 33057 55232
rect 33109 55229 33237 55232
rect 33289 55229 33327 55232
rect 33019 55189 33327 55229
rect 33484 55197 33816 55243
rect 33862 55197 34002 55243
rect 34048 55197 34189 55243
rect 34235 55197 34376 55243
rect 34422 55197 34562 55243
rect 34608 55197 35082 55243
rect 36438 55325 36475 55465
rect 36521 55325 36554 55465
rect 33484 55189 35082 55197
rect 35294 55191 36266 55231
rect 36438 55225 36554 55325
rect 36640 55465 36773 55488
rect 36640 55416 36697 55465
rect 36640 55364 36678 55416
rect 36640 55325 36697 55364
rect 36743 55325 36773 55465
rect 38658 55467 38726 55478
rect 36924 55457 37685 55463
rect 36923 55456 37685 55457
rect 36923 55423 37931 55456
rect 36923 55415 36961 55423
rect 37013 55415 37172 55423
rect 37224 55415 37384 55423
rect 36841 55369 36854 55415
rect 36900 55371 36961 55415
rect 36900 55369 36971 55371
rect 37017 55369 37088 55415
rect 37134 55371 37172 55415
rect 37134 55369 37206 55371
rect 37252 55369 37324 55415
rect 37370 55371 37384 55415
rect 37436 55415 37595 55423
rect 37436 55371 37442 55415
rect 37370 55369 37442 55371
rect 37488 55371 37595 55415
rect 37647 55415 37931 55423
rect 37647 55371 37909 55415
rect 37488 55369 37909 55371
rect 37955 55369 38026 55415
rect 38072 55369 38143 55415
rect 38189 55369 38261 55415
rect 38307 55369 38379 55415
rect 38425 55369 38497 55415
rect 38543 55369 38556 55415
rect 36923 55337 37931 55369
rect 36924 55330 37685 55337
rect 36640 55305 36773 55325
rect 38658 55327 38669 55467
rect 38715 55327 38726 55467
rect 39014 55415 39323 55901
rect 39492 55987 39608 56439
rect 39923 56406 40085 56537
rect 39923 56354 39994 56406
rect 40046 56354 40085 56406
rect 39923 56314 40085 56354
rect 39737 56218 39865 56231
rect 39737 56191 39866 56218
rect 39737 56174 39775 56191
rect 39827 56174 39866 56191
rect 39727 56128 39740 56174
rect 39827 56139 39862 56174
rect 39786 56128 39862 56139
rect 39908 56128 39985 56174
rect 40031 56128 40108 56174
rect 40154 56128 40167 56174
rect 40246 56163 40362 56561
rect 42229 56422 44509 56463
rect 42229 56370 42690 56422
rect 42742 56370 44509 56422
rect 42229 56330 44509 56370
rect 44341 56286 44509 56330
rect 44341 56240 44358 56286
rect 44498 56240 44509 56286
rect 39737 56099 39866 56128
rect 40246 56117 40281 56163
rect 40327 56117 40362 56163
rect 40246 56080 40362 56117
rect 40718 56191 43524 56232
rect 44341 56229 44509 56240
rect 40718 56139 41935 56191
rect 41987 56139 43524 56191
rect 40718 56098 43524 56139
rect 44605 56174 44721 56561
rect 45400 56531 48379 56572
rect 45400 56517 45975 56531
rect 45400 56471 45464 56517
rect 45604 56479 45975 56517
rect 46027 56479 48379 56531
rect 45604 56471 48379 56479
rect 44901 56415 45241 56456
rect 45400 56438 48379 56471
rect 48557 56525 48596 56577
rect 48648 56525 48687 56577
rect 48557 56502 48687 56525
rect 50044 56611 50516 56657
rect 50562 56611 50703 56657
rect 50749 56611 50890 56657
rect 50936 56611 51076 56657
rect 51122 56611 51263 56657
rect 51309 56611 51657 56657
rect 51797 56647 52105 56687
rect 51797 56622 51835 56647
rect 51887 56622 52015 56647
rect 52067 56622 52105 56647
rect 54085 56681 54223 56727
rect 54269 56687 54540 56727
rect 54269 56681 54440 56687
rect 54085 56641 54440 56681
rect 54486 56641 54540 56687
rect 50044 56574 51657 56611
rect 51789 56576 51802 56622
rect 53776 56576 53789 56622
rect 50044 56517 50160 56574
rect 44901 56398 44939 56415
rect 44991 56398 45151 56415
rect 45203 56398 45241 56415
rect 44799 56352 44812 56398
rect 44858 56352 44925 56398
rect 44991 56363 45038 56398
rect 44971 56352 45038 56363
rect 45084 56352 45151 56398
rect 45203 56363 45264 56398
rect 45197 56352 45264 56363
rect 45310 56352 45323 56398
rect 48557 56362 48622 56502
rect 48668 56362 48687 56502
rect 49820 56485 50160 56517
rect 48765 56439 48778 56485
rect 48824 56439 48881 56485
rect 48927 56439 48984 56485
rect 49030 56439 49087 56485
rect 49133 56439 49190 56485
rect 49236 56439 49293 56485
rect 49339 56439 49396 56485
rect 49442 56439 49499 56485
rect 49545 56439 49602 56485
rect 49852 56439 50160 56485
rect 51589 56522 51657 56574
rect 51797 56554 52105 56576
rect 49820 56398 50160 56439
rect 50262 56415 50812 56456
rect 48557 56359 48687 56362
rect 44901 56323 45241 56352
rect 48557 56307 48596 56359
rect 48648 56307 48687 56359
rect 50262 56363 50300 56415
rect 50352 56398 50511 56415
rect 50563 56398 50722 56415
rect 50352 56363 50467 56398
rect 50563 56363 50571 56398
rect 50262 56352 50467 56363
rect 50513 56352 50571 56363
rect 50617 56352 50674 56398
rect 50720 56363 50722 56398
rect 50774 56398 50812 56415
rect 50774 56363 50777 56398
rect 50720 56352 50777 56363
rect 50823 56352 50880 56398
rect 50926 56352 50983 56398
rect 51029 56352 51086 56398
rect 51132 56352 51189 56398
rect 51235 56352 51292 56398
rect 51338 56352 51395 56398
rect 51441 56352 51454 56398
rect 50262 56323 50812 56352
rect 48557 56266 48687 56307
rect 48905 56261 49877 56292
rect 48765 56215 48778 56261
rect 48824 56215 48881 56261
rect 48927 56252 48984 56261
rect 48927 56215 48943 56252
rect 49030 56215 49087 56261
rect 49133 56252 49190 56261
rect 49133 56215 49154 56252
rect 49236 56215 49293 56261
rect 49339 56252 49396 56261
rect 49339 56215 49365 56252
rect 49442 56215 49499 56261
rect 49545 56252 49602 56261
rect 49545 56215 49576 56252
rect 49852 56215 49877 56261
rect 48905 56200 48943 56215
rect 48995 56200 49154 56215
rect 49206 56200 49365 56215
rect 49417 56200 49576 56215
rect 49628 56200 49787 56215
rect 49839 56200 49877 56215
rect 44605 56128 44812 56174
rect 44858 56128 44925 56174
rect 44971 56128 45038 56174
rect 45084 56128 45151 56174
rect 45197 56128 45264 56174
rect 45310 56128 45323 56174
rect 48905 56160 49877 56200
rect 51035 56177 51343 56217
rect 51035 56174 51073 56177
rect 51125 56174 51253 56177
rect 51305 56174 51343 56177
rect 43362 56091 43524 56098
rect 43362 56045 43373 56091
rect 43513 56045 43524 56091
rect 43362 56034 43524 56045
rect 45584 56114 48546 56150
rect 50454 56128 50467 56174
rect 50513 56128 50571 56174
rect 50617 56128 50674 56174
rect 50720 56128 50777 56174
rect 50823 56128 50880 56174
rect 50926 56128 50983 56174
rect 51029 56128 51073 56174
rect 51132 56128 51189 56174
rect 51235 56128 51253 56174
rect 51338 56128 51395 56174
rect 51441 56128 51454 56174
rect 45584 56068 45619 56114
rect 45665 56068 45777 56114
rect 45823 56068 45935 56114
rect 45981 56068 46093 56114
rect 46139 56068 46251 56114
rect 46297 56068 46409 56114
rect 46455 56068 46568 56114
rect 46614 56068 46726 56114
rect 46772 56068 46884 56114
rect 46930 56068 47042 56114
rect 47088 56068 47200 56114
rect 47246 56068 47358 56114
rect 47404 56068 47516 56114
rect 47562 56068 47675 56114
rect 47721 56068 47833 56114
rect 47879 56068 47991 56114
rect 48037 56068 48149 56114
rect 48195 56068 48307 56114
rect 48353 56068 48465 56114
rect 48511 56068 48546 56114
rect 51035 56125 51073 56128
rect 51125 56125 51253 56128
rect 51305 56125 51343 56128
rect 51035 56084 51343 56125
rect 51589 56100 51600 56522
rect 51646 56100 51657 56522
rect 54085 56523 54540 56641
rect 54085 56477 54440 56523
rect 54486 56477 54540 56523
rect 54085 56449 54540 56477
rect 53585 56398 54540 56449
rect 51789 56352 51802 56398
rect 53776 56360 54540 56398
rect 53776 56352 54440 56360
rect 53585 56330 54440 56352
rect 54085 56314 54440 56330
rect 54486 56314 54540 56360
rect 54085 56238 54540 56314
rect 51797 56184 52105 56224
rect 51797 56174 51835 56184
rect 51887 56174 52015 56184
rect 52067 56174 52105 56184
rect 54085 56192 54223 56238
rect 54269 56197 54540 56238
rect 54269 56192 54440 56197
rect 51789 56128 51802 56174
rect 53776 56128 53789 56174
rect 54085 56151 54440 56192
rect 54486 56151 54540 56197
rect 51589 56089 51657 56100
rect 51797 56091 52105 56128
rect 40215 55987 40523 55994
rect 40788 55987 42986 56001
rect 43753 55987 44514 55994
rect 39492 55964 42986 55987
rect 43704 55964 44514 55987
rect 39492 55953 44514 55964
rect 39492 55950 40253 55953
rect 39492 55904 39740 55950
rect 39786 55904 39862 55950
rect 39908 55904 39985 55950
rect 40031 55904 40108 55950
rect 40154 55904 40253 55950
rect 39492 55901 40253 55904
rect 40305 55901 40433 55953
rect 40485 55950 43790 55953
rect 40485 55904 40836 55950
rect 40882 55904 40994 55950
rect 41040 55904 41152 55950
rect 41198 55904 41310 55950
rect 41356 55904 41469 55950
rect 41515 55904 41627 55950
rect 41673 55904 41785 55950
rect 41831 55904 41943 55950
rect 41989 55904 42101 55950
rect 42147 55904 42259 55950
rect 42305 55904 42418 55950
rect 42464 55904 42576 55950
rect 42622 55904 42734 55950
rect 42780 55904 42892 55950
rect 42938 55904 43739 55950
rect 43785 55904 43790 55950
rect 40485 55901 43790 55904
rect 43842 55950 44001 55953
rect 43842 55904 43906 55950
rect 43952 55904 44001 55950
rect 43842 55901 44001 55904
rect 44053 55950 44213 55953
rect 44265 55950 44424 55953
rect 44053 55904 44071 55950
rect 44117 55904 44213 55950
rect 44282 55904 44424 55950
rect 44053 55901 44213 55904
rect 44265 55901 44424 55904
rect 44476 55901 44514 55953
rect 39492 55890 44514 55901
rect 39492 55867 42986 55890
rect 43704 55867 44514 55890
rect 39492 55415 39608 55867
rect 40215 55860 40523 55867
rect 40788 55853 42986 55867
rect 43753 55860 44514 55867
rect 44796 55987 45346 55994
rect 45584 55987 48546 56068
rect 54085 56074 54540 56151
rect 54085 56028 54223 56074
rect 54269 56034 54540 56074
rect 54269 56028 54440 56034
rect 54085 55994 54440 56028
rect 48800 55987 49982 55994
rect 50308 55987 50859 55994
rect 44796 55953 49982 55987
rect 44796 55950 44834 55953
rect 44886 55950 45045 55953
rect 45097 55950 45256 55953
rect 45308 55950 48838 55953
rect 44796 55904 44812 55950
rect 44886 55904 44925 55950
rect 44971 55904 45038 55950
rect 45097 55904 45151 55950
rect 45197 55904 45256 55950
rect 45310 55904 45619 55950
rect 45665 55904 45777 55950
rect 45823 55904 45935 55950
rect 45981 55904 46093 55950
rect 46139 55904 46251 55950
rect 46297 55904 46409 55950
rect 46455 55904 46568 55950
rect 46614 55904 46726 55950
rect 46772 55904 46884 55950
rect 46930 55904 47042 55950
rect 47088 55904 47200 55950
rect 47246 55904 47358 55950
rect 47404 55904 47516 55950
rect 47562 55904 47675 55950
rect 47721 55904 47833 55950
rect 47879 55904 47991 55950
rect 48037 55904 48149 55950
rect 48195 55904 48307 55950
rect 48353 55904 48465 55950
rect 48511 55904 48838 55950
rect 44796 55901 44834 55904
rect 44886 55901 45045 55904
rect 45097 55901 45256 55904
rect 45308 55901 48838 55904
rect 48890 55901 49048 55953
rect 49100 55901 49259 55953
rect 49311 55901 49471 55953
rect 49523 55901 49682 55953
rect 49734 55901 49892 55953
rect 49944 55901 49982 55953
rect 44796 55867 49982 55901
rect 50307 55953 50859 55987
rect 50307 55901 50346 55953
rect 50398 55950 50557 55953
rect 50609 55950 50768 55953
rect 50820 55950 50859 55953
rect 52278 55988 54440 55994
rect 54486 55988 54540 56034
rect 55927 56687 57736 56801
rect 55927 56644 56267 56687
rect 55927 56598 55961 56644
rect 56007 56641 56267 56644
rect 56313 56641 57736 56687
rect 56007 56598 57736 56641
rect 55927 56523 57736 56598
rect 55927 56481 56267 56523
rect 55927 56435 55961 56481
rect 56007 56477 56267 56481
rect 56313 56477 57736 56523
rect 56007 56435 57736 56477
rect 55927 56360 57736 56435
rect 55927 56317 56267 56360
rect 55927 56271 55961 56317
rect 56007 56314 56267 56317
rect 56313 56314 57736 56360
rect 56007 56271 57736 56314
rect 55927 56197 57736 56271
rect 55927 56154 56267 56197
rect 55927 56108 55961 56154
rect 56007 56151 56267 56154
rect 56313 56151 57736 56197
rect 56007 56108 57736 56151
rect 55927 56034 57736 56108
rect 52278 55953 54540 55988
rect 52278 55950 52316 55953
rect 52368 55950 52527 55953
rect 52579 55950 52738 55953
rect 52790 55950 52948 55953
rect 53000 55950 53159 55953
rect 53211 55950 53371 55953
rect 53423 55950 53582 55953
rect 53634 55950 53792 55953
rect 50398 55904 50467 55950
rect 50513 55904 50557 55950
rect 50617 55904 50674 55950
rect 50720 55904 50768 55950
rect 50823 55904 50880 55950
rect 50926 55904 50983 55950
rect 51029 55904 51086 55950
rect 51132 55904 51189 55950
rect 51235 55904 51292 55950
rect 51338 55904 51395 55950
rect 51441 55904 51454 55950
rect 51789 55904 51802 55950
rect 53776 55904 53792 55950
rect 50398 55901 50557 55904
rect 50609 55901 50768 55904
rect 50820 55901 50859 55904
rect 50307 55867 50859 55901
rect 44796 55860 45346 55867
rect 43362 55809 43524 55820
rect 39737 55726 39866 55755
rect 40246 55737 40362 55774
rect 43362 55763 43373 55809
rect 43513 55763 43524 55809
rect 43362 55756 43524 55763
rect 39727 55680 39740 55726
rect 39786 55715 39862 55726
rect 39827 55680 39862 55715
rect 39908 55680 39985 55726
rect 40031 55680 40108 55726
rect 40154 55680 40167 55726
rect 40246 55691 40281 55737
rect 40327 55691 40362 55737
rect 39737 55663 39775 55680
rect 39827 55663 39866 55680
rect 39737 55636 39866 55663
rect 39737 55623 39865 55636
rect 39923 55500 40085 55540
rect 39923 55448 39994 55500
rect 40046 55448 40085 55500
rect 39008 55369 39021 55415
rect 39067 55369 39144 55415
rect 39190 55369 39267 55415
rect 39313 55369 39326 55415
rect 39492 55369 39641 55415
rect 39687 55369 39730 55415
rect 39014 55337 39323 55369
rect 39492 55337 39608 55369
rect 37853 55225 38161 55230
rect 36438 55191 36953 55225
rect 37439 55191 38161 55225
rect 38658 55205 38726 55327
rect 39923 55317 40085 55448
rect 39809 55314 40085 55317
rect 39809 55306 39994 55314
rect 39809 55260 39844 55306
rect 39890 55262 39994 55306
rect 40046 55293 40085 55314
rect 40246 55293 40362 55691
rect 40718 55715 43524 55756
rect 45584 55786 48546 55867
rect 48800 55860 49982 55867
rect 50308 55860 50859 55867
rect 52278 55901 52316 55904
rect 52368 55901 52527 55904
rect 52579 55901 52738 55904
rect 52790 55901 52948 55904
rect 53000 55901 53159 55904
rect 53211 55901 53371 55904
rect 53423 55901 53582 55904
rect 53634 55901 53792 55904
rect 53844 55901 54003 55953
rect 54055 55901 54214 55953
rect 54266 55901 54540 55953
rect 52278 55866 54540 55901
rect 52278 55860 54440 55866
rect 45584 55740 45619 55786
rect 45665 55740 45777 55786
rect 45823 55740 45935 55786
rect 45981 55740 46093 55786
rect 46139 55740 46251 55786
rect 46297 55740 46409 55786
rect 46455 55740 46568 55786
rect 46614 55740 46726 55786
rect 46772 55740 46884 55786
rect 46930 55740 47042 55786
rect 47088 55740 47200 55786
rect 47246 55740 47358 55786
rect 47404 55740 47516 55786
rect 47562 55740 47675 55786
rect 47721 55740 47833 55786
rect 47879 55740 47991 55786
rect 48037 55740 48149 55786
rect 48195 55740 48307 55786
rect 48353 55740 48465 55786
rect 48511 55740 48546 55786
rect 54085 55826 54440 55860
rect 54085 55780 54223 55826
rect 54269 55820 54440 55826
rect 54486 55820 54540 55866
rect 54758 55953 55840 55994
rect 54758 55950 54855 55953
rect 54758 55904 54793 55950
rect 54839 55904 54855 55950
rect 54758 55901 54855 55904
rect 54907 55950 55066 55953
rect 54907 55904 54956 55950
rect 55002 55904 55066 55950
rect 54907 55901 55066 55904
rect 55118 55950 55278 55953
rect 55330 55950 55489 55953
rect 55164 55904 55278 55950
rect 55330 55904 55439 55950
rect 55485 55904 55489 55950
rect 55118 55901 55278 55904
rect 55330 55901 55489 55904
rect 55541 55950 55840 55953
rect 55541 55904 55599 55950
rect 55645 55904 55760 55950
rect 55806 55904 55840 55950
rect 55541 55901 55840 55904
rect 54758 55861 55840 55901
rect 55927 55988 56267 56034
rect 56313 55988 57736 56034
rect 55927 55866 57736 55988
rect 54817 55860 55579 55861
rect 54269 55780 54540 55820
rect 40718 55663 41935 55715
rect 41987 55663 43524 55715
rect 40718 55622 43524 55663
rect 44605 55680 44812 55726
rect 44858 55680 44925 55726
rect 44971 55680 45038 55726
rect 45084 55680 45151 55726
rect 45197 55680 45264 55726
rect 45310 55680 45323 55726
rect 45584 55704 48546 55740
rect 51035 55729 51343 55770
rect 51035 55726 51073 55729
rect 51125 55726 51253 55729
rect 51305 55726 51343 55729
rect 51589 55754 51657 55765
rect 44341 55614 44509 55625
rect 44341 55568 44358 55614
rect 44498 55568 44509 55614
rect 44341 55524 44509 55568
rect 42229 55484 44509 55524
rect 42229 55432 42690 55484
rect 42742 55432 44509 55484
rect 42229 55391 44509 55432
rect 44605 55293 44721 55680
rect 48905 55654 49877 55694
rect 50454 55680 50467 55726
rect 50513 55680 50571 55726
rect 50617 55680 50674 55726
rect 50720 55680 50777 55726
rect 50823 55680 50880 55726
rect 50926 55680 50983 55726
rect 51029 55680 51073 55726
rect 51132 55680 51189 55726
rect 51235 55680 51253 55726
rect 51338 55680 51395 55726
rect 51441 55680 51454 55726
rect 48905 55639 48943 55654
rect 48995 55639 49154 55654
rect 49206 55639 49365 55654
rect 49417 55639 49576 55654
rect 49628 55639 49787 55654
rect 49839 55639 49877 55654
rect 48765 55593 48778 55639
rect 48824 55593 48881 55639
rect 48927 55602 48943 55639
rect 48927 55593 48984 55602
rect 49030 55593 49087 55639
rect 49133 55602 49154 55639
rect 49133 55593 49190 55602
rect 49236 55593 49293 55639
rect 49339 55602 49365 55639
rect 49339 55593 49396 55602
rect 49442 55593 49499 55639
rect 49545 55602 49576 55639
rect 49545 55593 49602 55602
rect 49852 55593 49877 55639
rect 51035 55677 51073 55680
rect 51125 55677 51253 55680
rect 51305 55677 51343 55680
rect 51035 55637 51343 55677
rect 48557 55547 48687 55588
rect 48905 55562 49877 55593
rect 44901 55502 45241 55531
rect 44799 55456 44812 55502
rect 44858 55456 44925 55502
rect 44971 55491 45038 55502
rect 44991 55456 45038 55491
rect 45084 55456 45151 55502
rect 45197 55491 45264 55502
rect 45203 55456 45264 55491
rect 45310 55456 45323 55502
rect 48557 55495 48596 55547
rect 48648 55495 48687 55547
rect 48557 55492 48687 55495
rect 44901 55439 44939 55456
rect 44991 55439 45151 55456
rect 45203 55439 45241 55456
rect 44901 55398 45241 55439
rect 45400 55383 48379 55416
rect 45400 55337 45464 55383
rect 45604 55375 48379 55383
rect 45604 55337 46353 55375
rect 45400 55323 46353 55337
rect 46405 55323 48379 55375
rect 40046 55278 44918 55293
rect 45400 55282 48379 55323
rect 48557 55352 48622 55492
rect 48668 55352 48687 55492
rect 50262 55502 50812 55531
rect 50262 55491 50467 55502
rect 50513 55491 50571 55502
rect 49820 55415 50160 55456
rect 48765 55369 48778 55415
rect 48824 55369 48881 55415
rect 48927 55369 48984 55415
rect 49030 55369 49087 55415
rect 49133 55369 49190 55415
rect 49236 55369 49293 55415
rect 49339 55369 49396 55415
rect 49442 55369 49499 55415
rect 49545 55369 49602 55415
rect 49852 55369 50160 55415
rect 50262 55439 50300 55491
rect 50352 55456 50467 55491
rect 50563 55456 50571 55491
rect 50617 55456 50674 55502
rect 50720 55491 50777 55502
rect 50720 55456 50722 55491
rect 50352 55439 50511 55456
rect 50563 55439 50722 55456
rect 50774 55456 50777 55491
rect 50823 55456 50880 55502
rect 50926 55456 50983 55502
rect 51029 55456 51086 55502
rect 51132 55456 51189 55502
rect 51235 55456 51292 55502
rect 51338 55456 51395 55502
rect 51441 55456 51454 55502
rect 50774 55439 50812 55456
rect 50262 55398 50812 55439
rect 48557 55329 48687 55352
rect 49820 55337 50160 55369
rect 40046 55262 44812 55278
rect 39890 55260 44812 55262
rect 39809 55257 44812 55260
rect 39809 55211 43739 55257
rect 43785 55211 43906 55257
rect 43952 55211 44071 55257
rect 44117 55211 44236 55257
rect 44282 55232 44812 55257
rect 44858 55232 44925 55278
rect 44971 55232 45038 55278
rect 45084 55232 45151 55278
rect 45197 55232 45264 55278
rect 45310 55232 45323 55278
rect 48557 55277 48596 55329
rect 48648 55277 48687 55329
rect 48557 55237 48687 55277
rect 50044 55280 50160 55337
rect 51589 55332 51600 55754
rect 51646 55332 51657 55754
rect 51797 55726 52105 55763
rect 51789 55680 51802 55726
rect 53776 55680 53789 55726
rect 54085 55703 54540 55780
rect 51797 55670 51835 55680
rect 51887 55670 52015 55680
rect 52067 55670 52105 55680
rect 51797 55630 52105 55670
rect 54085 55662 54440 55703
rect 54085 55616 54223 55662
rect 54269 55657 54440 55662
rect 54486 55657 54540 55703
rect 54269 55616 54540 55657
rect 54085 55540 54540 55616
rect 54085 55524 54440 55540
rect 53585 55502 54440 55524
rect 51789 55456 51802 55502
rect 53776 55494 54440 55502
rect 54486 55494 54540 55540
rect 53776 55456 54540 55494
rect 53585 55405 54540 55456
rect 51589 55280 51657 55332
rect 54085 55377 54540 55405
rect 54085 55331 54440 55377
rect 54486 55331 54540 55377
rect 50044 55243 51657 55280
rect 51797 55278 52105 55300
rect 44282 55211 44918 55232
rect 38658 55191 39723 55205
rect 30683 55167 30855 55173
rect 30583 55127 30855 55167
rect 30901 55127 31040 55173
rect 33484 55160 34643 55189
rect 35260 55145 35273 55191
rect 35523 55145 35543 55191
rect 35626 55145 35683 55191
rect 35729 55145 35754 55191
rect 35832 55145 35889 55191
rect 35935 55145 35965 55191
rect 36038 55145 36095 55191
rect 36141 55145 36176 55191
rect 36244 55145 36301 55191
rect 36347 55145 36360 55191
rect 36438 55145 36854 55191
rect 36900 55145 36971 55191
rect 37017 55145 37088 55191
rect 37134 55145 37206 55191
rect 37252 55145 37324 55191
rect 37370 55145 37442 55191
rect 37488 55189 37909 55191
rect 37488 55145 37891 55189
rect 37955 55145 38026 55191
rect 38072 55189 38143 55191
rect 38123 55145 38143 55189
rect 38189 55145 38261 55191
rect 38307 55145 38379 55191
rect 38425 55145 38497 55191
rect 38543 55145 38556 55191
rect 38658 55145 39021 55191
rect 39067 55145 39144 55191
rect 39190 55145 39267 55191
rect 39313 55145 39641 55191
rect 39687 55145 39730 55191
rect 39809 55173 44918 55211
rect 48905 55191 49877 55231
rect 48765 55145 48778 55191
rect 48824 55145 48881 55191
rect 48927 55145 48943 55191
rect 49030 55145 49087 55191
rect 49133 55145 49154 55191
rect 49236 55145 49293 55191
rect 49339 55145 49365 55191
rect 49442 55145 49499 55191
rect 49545 55145 49576 55191
rect 49852 55145 49877 55191
rect 50044 55197 50516 55243
rect 50562 55197 50703 55243
rect 50749 55197 50890 55243
rect 50936 55197 51076 55243
rect 51122 55197 51263 55243
rect 51309 55197 51657 55243
rect 51789 55232 51802 55278
rect 53776 55232 53789 55278
rect 50044 55187 51657 55197
rect 50481 55160 51657 55187
rect 51797 55207 51835 55232
rect 51887 55207 52015 55232
rect 52067 55207 52105 55232
rect 51797 55167 52105 55207
rect 54085 55213 54540 55331
rect 54085 55173 54440 55213
rect 30583 55094 31040 55127
rect 35294 55139 35332 55145
rect 35384 55139 35543 55145
rect 35595 55139 35754 55145
rect 35806 55139 35965 55145
rect 36017 55139 36176 55145
rect 36228 55139 36266 55145
rect 34870 55094 35025 55101
rect 35294 55099 36266 55139
rect 36438 55105 36953 55145
rect 37439 55137 37891 55145
rect 37943 55137 38071 55145
rect 38123 55137 38161 55145
rect 37439 55105 38161 55137
rect 37853 55097 38161 55105
rect 27387 55001 27790 55053
rect 27842 55001 28001 55053
rect 28053 55001 28212 55053
rect 28264 55001 28423 55053
rect 28475 55001 28634 55053
rect 28686 55050 28845 55053
rect 28686 55004 28810 55050
rect 28686 55001 28845 55004
rect 28897 55001 29056 55053
rect 29108 55001 29196 55053
rect 27387 54887 29196 55001
rect 29283 55053 30365 55094
rect 29283 55050 29582 55053
rect 29283 55004 29317 55050
rect 29363 55004 29478 55050
rect 29524 55004 29582 55050
rect 29283 55001 29582 55004
rect 29634 55050 29793 55053
rect 29845 55050 30005 55053
rect 29634 55004 29638 55050
rect 29684 55004 29793 55050
rect 29845 55004 29959 55050
rect 29634 55001 29793 55004
rect 29845 55001 30005 55004
rect 30057 55050 30216 55053
rect 30057 55004 30121 55050
rect 30167 55004 30216 55050
rect 30057 55001 30216 55004
rect 30268 55050 30365 55053
rect 30268 55004 30284 55050
rect 30330 55004 30365 55050
rect 30268 55001 30365 55004
rect 29283 54961 30365 55001
rect 30583 55053 32842 55094
rect 30583 55050 30854 55053
rect 30583 55004 30637 55050
rect 30683 55004 30854 55050
rect 30583 55001 30854 55004
rect 30906 55001 31065 55053
rect 31117 55001 31276 55053
rect 31328 55001 31486 55053
rect 31538 55001 31697 55053
rect 31749 55001 31909 55053
rect 31961 55001 32120 55053
rect 32172 55001 32330 55053
rect 32382 55001 32541 55053
rect 32593 55001 32752 55053
rect 32804 55001 32842 55053
rect 29544 54960 30306 54961
rect 30583 54960 32842 55001
rect 34717 55053 35025 55094
rect 38658 55085 39723 55145
rect 48905 55139 48943 55145
rect 48995 55139 49154 55145
rect 49206 55139 49365 55145
rect 49417 55139 49576 55145
rect 49628 55139 49787 55145
rect 49839 55139 49877 55145
rect 48905 55099 49877 55139
rect 54085 55127 54223 55173
rect 54269 55167 54440 55173
rect 54486 55167 54540 55213
rect 54269 55127 54540 55167
rect 50099 55094 50255 55101
rect 54085 55094 54540 55127
rect 55927 55820 56267 55866
rect 56313 55820 57736 55866
rect 55927 55744 57736 55820
rect 55927 55698 55961 55744
rect 56007 55703 57736 55744
rect 56007 55698 56267 55703
rect 55927 55657 56267 55698
rect 56313 55657 57736 55703
rect 55927 55581 57736 55657
rect 55927 55535 55961 55581
rect 56007 55540 57736 55581
rect 56007 55535 56267 55540
rect 55927 55494 56267 55535
rect 56313 55494 57736 55540
rect 55927 55417 57736 55494
rect 55927 55371 55961 55417
rect 56007 55377 57736 55417
rect 56007 55371 56267 55377
rect 55927 55331 56267 55371
rect 56313 55331 57736 55377
rect 55927 55254 57736 55331
rect 55927 55208 55961 55254
rect 56007 55213 57736 55254
rect 56007 55208 56267 55213
rect 55927 55167 56267 55208
rect 56313 55167 57736 55213
rect 34717 55001 34755 55053
rect 34807 55050 34935 55053
rect 34807 55004 34916 55050
rect 34807 55001 34935 55004
rect 34987 55001 35025 55053
rect 34717 54960 35025 55001
rect 50099 55053 50408 55094
rect 50099 55001 50138 55053
rect 50190 55050 50318 55053
rect 50206 55004 50318 55050
rect 50190 55001 50318 55004
rect 50370 55001 50408 55053
rect 27387 54841 28810 54887
rect 28856 54844 29196 54887
rect 28856 54841 29116 54844
rect 27387 54798 29116 54841
rect 29162 54798 29196 54844
rect 27387 54723 29196 54798
rect 27387 54677 28810 54723
rect 28856 54681 29196 54723
rect 28856 54677 29116 54681
rect 27387 54635 29116 54677
rect 29162 54635 29196 54681
rect 27387 54560 29196 54635
rect 27387 54514 28810 54560
rect 28856 54517 29196 54560
rect 28856 54514 29116 54517
rect 27387 54471 29116 54514
rect 29162 54471 29196 54517
rect 27387 54397 29196 54471
rect 27387 54351 28810 54397
rect 28856 54354 29196 54397
rect 28856 54351 29116 54354
rect 27387 54308 29116 54351
rect 29162 54308 29196 54354
rect 27387 54234 29196 54308
rect 27387 54188 28810 54234
rect 28856 54188 29196 54234
rect 30583 54927 31040 54960
rect 34870 54953 35025 54960
rect 30583 54887 30855 54927
rect 30583 54841 30637 54887
rect 30683 54881 30855 54887
rect 30901 54881 31040 54927
rect 35294 54915 36266 54955
rect 37853 54949 38161 54957
rect 35294 54909 35332 54915
rect 35384 54909 35543 54915
rect 35595 54909 35754 54915
rect 35806 54909 35965 54915
rect 36017 54909 36176 54915
rect 36228 54909 36266 54915
rect 36438 54909 36953 54949
rect 37439 54917 38161 54949
rect 37439 54909 37891 54917
rect 37943 54909 38071 54917
rect 38123 54909 38161 54917
rect 38658 54909 39723 54969
rect 50099 54960 50408 55001
rect 52278 55053 54540 55094
rect 52278 55001 52316 55053
rect 52368 55001 52527 55053
rect 52579 55001 52738 55053
rect 52790 55001 52948 55053
rect 53000 55001 53159 55053
rect 53211 55001 53371 55053
rect 53423 55001 53582 55053
rect 53634 55001 53792 55053
rect 53844 55001 54003 55053
rect 54055 55001 54214 55053
rect 54266 55050 54540 55053
rect 54266 55004 54440 55050
rect 54486 55004 54540 55050
rect 54266 55001 54540 55004
rect 52278 54960 54540 55001
rect 54758 55053 55840 55094
rect 54758 55050 54855 55053
rect 54758 55004 54793 55050
rect 54839 55004 54855 55050
rect 54758 55001 54855 55004
rect 54907 55050 55066 55053
rect 54907 55004 54956 55050
rect 55002 55004 55066 55050
rect 54907 55001 55066 55004
rect 55118 55050 55278 55053
rect 55330 55050 55489 55053
rect 55164 55004 55278 55050
rect 55330 55004 55439 55050
rect 55485 55004 55489 55050
rect 55118 55001 55278 55004
rect 55330 55001 55489 55004
rect 55541 55050 55840 55053
rect 55541 55004 55599 55050
rect 55645 55004 55760 55050
rect 55806 55004 55840 55050
rect 55541 55001 55840 55004
rect 54758 54961 55840 55001
rect 55927 55053 57736 55167
rect 55927 55001 56015 55053
rect 56067 55001 56226 55053
rect 56278 55050 56437 55053
rect 56313 55004 56437 55050
rect 56278 55001 56437 55004
rect 56489 55001 56648 55053
rect 56700 55001 56859 55053
rect 56911 55001 57070 55053
rect 57122 55001 57281 55053
rect 57333 55001 57736 55053
rect 54817 54960 55579 54961
rect 48905 54915 49877 54955
rect 50099 54953 50255 54960
rect 48905 54909 48943 54915
rect 48995 54909 49154 54915
rect 49206 54909 49365 54915
rect 49417 54909 49576 54915
rect 49628 54909 49787 54915
rect 49839 54909 49877 54915
rect 30683 54841 31040 54881
rect 33484 54865 34643 54894
rect 30583 54764 31040 54841
rect 33019 54825 33327 54865
rect 33019 54822 33057 54825
rect 33109 54822 33237 54825
rect 33289 54822 33327 54825
rect 33484 54857 35082 54865
rect 35260 54863 35273 54909
rect 35523 54863 35543 54909
rect 35626 54863 35683 54909
rect 35729 54863 35754 54909
rect 35832 54863 35889 54909
rect 35935 54863 35965 54909
rect 36038 54863 36095 54909
rect 36141 54863 36176 54909
rect 36244 54863 36301 54909
rect 36347 54863 36360 54909
rect 36438 54863 36854 54909
rect 36900 54863 36971 54909
rect 37017 54863 37088 54909
rect 37134 54863 37206 54909
rect 37252 54863 37324 54909
rect 37370 54863 37442 54909
rect 37488 54865 37891 54909
rect 37488 54863 37909 54865
rect 37955 54863 38026 54909
rect 38123 54865 38143 54909
rect 38072 54863 38143 54865
rect 38189 54863 38261 54909
rect 38307 54863 38379 54909
rect 38425 54863 38497 54909
rect 38543 54863 38556 54909
rect 38658 54863 39021 54909
rect 39067 54863 39144 54909
rect 39190 54863 39267 54909
rect 39313 54863 39641 54909
rect 39687 54863 39730 54909
rect 31336 54776 31349 54822
rect 33323 54776 33336 54822
rect 33484 54811 33816 54857
rect 33862 54811 34002 54857
rect 34048 54811 34189 54857
rect 34235 54811 34376 54857
rect 34422 54811 34562 54857
rect 34608 54811 35082 54857
rect 35294 54823 36266 54863
rect 36438 54829 36953 54863
rect 37439 54829 38161 54863
rect 30583 54723 30855 54764
rect 30583 54677 30637 54723
rect 30683 54718 30855 54723
rect 30901 54718 31040 54764
rect 33019 54773 33057 54776
rect 33109 54773 33237 54776
rect 33289 54773 33327 54776
rect 33019 54732 33327 54773
rect 33484 54774 35082 54811
rect 30683 54677 31040 54718
rect 30583 54649 31040 54677
rect 33484 54692 33552 54774
rect 30583 54601 31493 54649
rect 30583 54560 30855 54601
rect 30583 54514 30637 54560
rect 30683 54555 30855 54560
rect 30901 54598 31493 54601
rect 30901 54555 31349 54598
rect 30683 54552 31349 54555
rect 33323 54552 33336 54598
rect 30683 54530 31493 54552
rect 30683 54514 31040 54530
rect 30583 54438 31040 54514
rect 30583 54397 30855 54438
rect 30583 54351 30637 54397
rect 30683 54392 30855 54397
rect 30901 54392 31040 54438
rect 30683 54351 31040 54392
rect 33019 54377 33327 54417
rect 33019 54374 33057 54377
rect 33109 54374 33237 54377
rect 33289 54374 33327 54377
rect 30583 54274 31040 54351
rect 31336 54328 31349 54374
rect 33323 54328 33336 54374
rect 33019 54325 33057 54328
rect 33109 54325 33237 54328
rect 33289 54325 33327 54328
rect 33019 54284 33327 54325
rect 30583 54234 30855 54274
rect 27387 54066 29196 54188
rect 27387 54020 28810 54066
rect 28856 54020 29196 54066
rect 29283 54153 30365 54194
rect 29283 54150 29582 54153
rect 29283 54104 29317 54150
rect 29363 54104 29478 54150
rect 29524 54104 29582 54150
rect 29283 54101 29582 54104
rect 29634 54150 29793 54153
rect 29845 54150 30005 54153
rect 29634 54104 29638 54150
rect 29684 54104 29793 54150
rect 29845 54104 29959 54150
rect 29634 54101 29793 54104
rect 29845 54101 30005 54104
rect 30057 54150 30216 54153
rect 30057 54104 30121 54150
rect 30167 54104 30216 54150
rect 30057 54101 30216 54104
rect 30268 54150 30365 54153
rect 30268 54104 30284 54150
rect 30330 54104 30365 54150
rect 30268 54101 30365 54104
rect 29283 54061 30365 54101
rect 30583 54188 30637 54234
rect 30683 54228 30855 54234
rect 30901 54228 31040 54274
rect 33484 54270 33495 54692
rect 33541 54270 33552 54692
rect 34964 54717 35082 54774
rect 36438 54729 36554 54829
rect 37853 54824 38161 54829
rect 38658 54849 39723 54863
rect 34964 54685 36360 54717
rect 34228 54615 34718 54656
rect 34228 54598 34267 54615
rect 34319 54598 34447 54615
rect 34499 54598 34627 54615
rect 33671 54552 33684 54598
rect 33730 54552 33787 54598
rect 33833 54552 33890 54598
rect 33936 54552 33993 54598
rect 34039 54552 34096 54598
rect 34142 54552 34199 54598
rect 34245 54563 34267 54598
rect 34245 54552 34302 54563
rect 34348 54552 34405 54598
rect 34499 54563 34508 54598
rect 34451 54552 34508 54563
rect 34554 54552 34612 54598
rect 34679 54563 34718 54615
rect 34964 54639 35273 54685
rect 35523 54639 35580 54685
rect 35626 54639 35683 54685
rect 35729 54639 35786 54685
rect 35832 54639 35889 54685
rect 35935 54639 35992 54685
rect 36038 54639 36095 54685
rect 36141 54639 36198 54685
rect 36244 54639 36301 54685
rect 36347 54639 36360 54685
rect 34964 54595 36360 54639
rect 34658 54552 34718 54563
rect 34228 54523 34718 54552
rect 36438 54589 36475 54729
rect 36521 54589 36554 54729
rect 35294 54461 36266 54495
rect 36438 54486 36554 54589
rect 36640 54729 36773 54749
rect 36640 54690 36697 54729
rect 36640 54638 36678 54690
rect 36640 54589 36697 54638
rect 36743 54589 36773 54729
rect 38658 54727 38726 54849
rect 39809 54843 44918 54881
rect 48765 54863 48778 54909
rect 48824 54863 48881 54909
rect 48927 54863 48943 54909
rect 49030 54863 49087 54909
rect 49133 54863 49154 54909
rect 49236 54863 49293 54909
rect 49339 54863 49365 54909
rect 49442 54863 49499 54909
rect 49545 54863 49576 54909
rect 49852 54863 49877 54909
rect 54085 54927 54540 54960
rect 50481 54867 51657 54894
rect 39809 54797 43739 54843
rect 43785 54797 43906 54843
rect 43952 54797 44071 54843
rect 44117 54797 44236 54843
rect 44282 54822 44918 54843
rect 48905 54823 49877 54863
rect 50044 54857 51657 54867
rect 44282 54797 44812 54822
rect 39809 54794 44812 54797
rect 39809 54748 39844 54794
rect 39890 54792 44812 54794
rect 39890 54748 39994 54792
rect 39809 54740 39994 54748
rect 40046 54776 44812 54792
rect 44858 54776 44925 54822
rect 44971 54776 45038 54822
rect 45084 54776 45151 54822
rect 45197 54776 45264 54822
rect 45310 54776 45323 54822
rect 48557 54777 48687 54817
rect 40046 54761 44918 54776
rect 40046 54740 40085 54761
rect 39809 54737 40085 54740
rect 36924 54717 37685 54724
rect 36923 54685 37931 54717
rect 36841 54639 36854 54685
rect 36900 54683 36971 54685
rect 36900 54639 36961 54683
rect 37017 54639 37088 54685
rect 37134 54683 37206 54685
rect 37134 54639 37172 54683
rect 37252 54639 37324 54685
rect 37370 54683 37442 54685
rect 37370 54639 37384 54683
rect 36923 54631 36961 54639
rect 37013 54631 37172 54639
rect 37224 54631 37384 54639
rect 37436 54639 37442 54683
rect 37488 54683 37909 54685
rect 37488 54639 37595 54683
rect 37436 54631 37595 54639
rect 37647 54639 37909 54683
rect 37955 54639 38026 54685
rect 38072 54639 38143 54685
rect 38189 54639 38261 54685
rect 38307 54639 38379 54685
rect 38425 54639 38497 54685
rect 38543 54639 38556 54685
rect 37647 54631 37931 54639
rect 36923 54598 37931 54631
rect 36923 54597 37685 54598
rect 36924 54591 37685 54597
rect 36640 54566 36773 54589
rect 38658 54587 38669 54727
rect 38715 54587 38726 54727
rect 39014 54685 39323 54717
rect 39492 54685 39608 54717
rect 39008 54639 39021 54685
rect 39067 54639 39144 54685
rect 39190 54639 39267 54685
rect 39313 54639 39326 54685
rect 39492 54639 39641 54685
rect 39687 54639 39730 54685
rect 38658 54576 38726 54587
rect 36438 54461 36953 54486
rect 37439 54483 37931 54486
rect 37439 54461 38161 54483
rect 35260 54415 35273 54461
rect 35523 54455 35580 54461
rect 35523 54415 35543 54455
rect 35626 54415 35683 54461
rect 35729 54455 35786 54461
rect 35729 54415 35754 54455
rect 35832 54415 35889 54461
rect 35935 54455 35992 54461
rect 35935 54415 35965 54455
rect 36038 54415 36095 54461
rect 36141 54455 36198 54461
rect 36141 54415 36176 54455
rect 36244 54415 36301 54461
rect 36347 54415 36360 54461
rect 36438 54415 36854 54461
rect 36900 54415 36971 54461
rect 37017 54415 37088 54461
rect 37134 54415 37206 54461
rect 37252 54415 37324 54461
rect 37370 54415 37442 54461
rect 37488 54443 37909 54461
rect 37488 54415 37891 54443
rect 37955 54415 38026 54461
rect 38072 54443 38143 54461
rect 38123 54415 38143 54443
rect 38189 54415 38261 54461
rect 38307 54415 38379 54461
rect 38425 54415 38497 54461
rect 38543 54415 38556 54461
rect 33781 54374 34089 54409
rect 35294 54403 35332 54415
rect 35384 54403 35543 54415
rect 35595 54403 35754 54415
rect 35806 54403 35965 54415
rect 36017 54403 36176 54415
rect 36228 54403 36266 54415
rect 33671 54328 33684 54374
rect 33730 54328 33787 54374
rect 33833 54369 33890 54374
rect 33871 54328 33890 54369
rect 33936 54328 33993 54374
rect 34039 54369 34096 54374
rect 34051 54328 34096 54369
rect 34142 54328 34199 54374
rect 34245 54328 34302 54374
rect 34348 54328 34405 54374
rect 34451 54328 34508 54374
rect 34554 54328 34612 54374
rect 34658 54328 34671 54374
rect 35294 54363 36266 54403
rect 36438 54366 36953 54415
rect 37439 54391 37891 54415
rect 37943 54391 38071 54415
rect 38123 54391 38161 54415
rect 37439 54366 38161 54391
rect 37853 54350 38161 54366
rect 33781 54317 33819 54328
rect 33871 54317 33999 54328
rect 34051 54317 34089 54328
rect 33781 54276 34089 54317
rect 33484 54259 33552 54270
rect 30683 54194 31040 54228
rect 30683 54188 32842 54194
rect 30583 54153 32842 54188
rect 34247 54187 35008 54194
rect 30583 54101 30854 54153
rect 30906 54101 31065 54153
rect 31117 54101 31276 54153
rect 31328 54150 31486 54153
rect 31538 54150 31697 54153
rect 31749 54150 31909 54153
rect 31961 54150 32120 54153
rect 32172 54150 32330 54153
rect 32382 54150 32541 54153
rect 32593 54150 32752 54153
rect 32804 54150 32842 54153
rect 34246 54153 35008 54187
rect 34246 54150 34284 54153
rect 34336 54150 34495 54153
rect 34547 54150 34707 54153
rect 31328 54104 31349 54150
rect 33323 54104 33336 54150
rect 33671 54104 33684 54150
rect 33730 54104 33787 54150
rect 33833 54104 33890 54150
rect 33936 54104 33993 54150
rect 34039 54104 34096 54150
rect 34142 54104 34199 54150
rect 34245 54104 34284 54150
rect 34348 54104 34405 54150
rect 34451 54104 34495 54150
rect 34554 54104 34612 54150
rect 34658 54104 34707 54150
rect 31328 54101 31486 54104
rect 31538 54101 31697 54104
rect 31749 54101 31909 54104
rect 31961 54101 32120 54104
rect 32172 54101 32330 54104
rect 32382 54101 32541 54104
rect 32593 54101 32752 54104
rect 32804 54101 32842 54104
rect 30583 54066 32842 54101
rect 34246 54101 34284 54104
rect 34336 54101 34495 54104
rect 34547 54101 34707 54104
rect 34759 54101 34918 54153
rect 34970 54101 35008 54153
rect 34246 54067 35008 54101
rect 29544 54060 30306 54061
rect 27387 53944 29196 54020
rect 27387 53903 29116 53944
rect 27387 53857 28810 53903
rect 28856 53898 29116 53903
rect 29162 53898 29196 53944
rect 28856 53857 29196 53898
rect 27387 53781 29196 53857
rect 27387 53740 29116 53781
rect 27387 53694 28810 53740
rect 28856 53735 29116 53740
rect 29162 53735 29196 53781
rect 28856 53694 29196 53735
rect 27387 53617 29196 53694
rect 27387 53577 29116 53617
rect 27387 53531 28810 53577
rect 28856 53571 29116 53577
rect 29162 53571 29196 53617
rect 28856 53531 29196 53571
rect 27387 53454 29196 53531
rect 27387 53413 29116 53454
rect 27387 53367 28810 53413
rect 28856 53408 29116 53413
rect 29162 53408 29196 53454
rect 28856 53367 29196 53408
rect 27387 53253 29196 53367
rect 30583 54020 30637 54066
rect 30683 54060 32842 54066
rect 34247 54060 35008 54067
rect 35182 54187 36364 54194
rect 35182 54153 36958 54187
rect 35182 54101 35220 54153
rect 35272 54101 35430 54153
rect 35482 54101 35641 54153
rect 35693 54101 35853 54153
rect 35905 54101 36064 54153
rect 36116 54101 36274 54153
rect 36326 54150 36958 54153
rect 36326 54104 36489 54150
rect 36723 54104 36958 54150
rect 36326 54101 36958 54104
rect 35182 54067 36958 54101
rect 37946 54153 38842 54194
rect 37946 54150 38330 54153
rect 38382 54150 38541 54153
rect 37946 54104 37957 54150
rect 38473 54104 38541 54150
rect 37946 54101 38330 54104
rect 38382 54101 38541 54104
rect 38593 54101 38752 54153
rect 38804 54101 38842 54153
rect 35182 54060 36364 54067
rect 37946 54060 38842 54101
rect 39014 54153 39323 54639
rect 39014 54101 39052 54153
rect 39104 54150 39232 54153
rect 39108 54104 39220 54150
rect 39104 54101 39232 54104
rect 39284 54101 39323 54153
rect 30683 54026 31040 54060
rect 30683 54020 30855 54026
rect 30583 53980 30855 54020
rect 30901 53980 31040 54026
rect 30583 53903 31040 53980
rect 33484 53984 33552 53995
rect 33019 53929 33327 53970
rect 33019 53926 33057 53929
rect 33109 53926 33237 53929
rect 33289 53926 33327 53929
rect 30583 53857 30637 53903
rect 30683 53862 31040 53903
rect 31336 53880 31349 53926
rect 33323 53880 33336 53926
rect 30683 53857 30855 53862
rect 30583 53816 30855 53857
rect 30901 53816 31040 53862
rect 33019 53877 33057 53880
rect 33109 53877 33237 53880
rect 33289 53877 33327 53880
rect 33019 53837 33327 53877
rect 30583 53740 31040 53816
rect 30583 53694 30637 53740
rect 30683 53724 31040 53740
rect 30683 53702 31493 53724
rect 30683 53699 31349 53702
rect 30683 53694 30855 53699
rect 30583 53653 30855 53694
rect 30901 53656 31349 53699
rect 33323 53656 33336 53702
rect 30901 53653 31493 53656
rect 30583 53605 31493 53653
rect 30583 53577 31040 53605
rect 30583 53531 30637 53577
rect 30683 53536 31040 53577
rect 30683 53531 30855 53536
rect 30583 53490 30855 53531
rect 30901 53490 31040 53536
rect 33484 53562 33495 53984
rect 33541 53562 33552 53984
rect 33781 53937 34089 53978
rect 33781 53926 33819 53937
rect 33871 53926 33999 53937
rect 34051 53926 34089 53937
rect 33671 53880 33684 53926
rect 33730 53880 33787 53926
rect 33871 53885 33890 53926
rect 33833 53880 33890 53885
rect 33936 53880 33993 53926
rect 34051 53885 34096 53926
rect 34039 53880 34096 53885
rect 34142 53880 34199 53926
rect 34245 53880 34302 53926
rect 34348 53880 34405 53926
rect 34451 53880 34508 53926
rect 34554 53880 34612 53926
rect 34658 53880 34671 53926
rect 33781 53845 34089 53880
rect 35294 53851 36266 53891
rect 37853 53888 38161 53904
rect 35294 53839 35332 53851
rect 35384 53839 35543 53851
rect 35595 53839 35754 53851
rect 35806 53839 35965 53851
rect 36017 53839 36176 53851
rect 36228 53839 36266 53851
rect 36438 53839 36953 53888
rect 37439 53863 38161 53888
rect 37439 53839 37891 53863
rect 37943 53839 38071 53863
rect 38123 53839 38161 53863
rect 35260 53793 35273 53839
rect 35523 53799 35543 53839
rect 35523 53793 35580 53799
rect 35626 53793 35683 53839
rect 35729 53799 35754 53839
rect 35729 53793 35786 53799
rect 35832 53793 35889 53839
rect 35935 53799 35965 53839
rect 35935 53793 35992 53799
rect 36038 53793 36095 53839
rect 36141 53799 36176 53839
rect 36141 53793 36198 53799
rect 36244 53793 36301 53839
rect 36347 53793 36360 53839
rect 36438 53793 36854 53839
rect 36900 53793 36971 53839
rect 37017 53793 37088 53839
rect 37134 53793 37206 53839
rect 37252 53793 37324 53839
rect 37370 53793 37442 53839
rect 37488 53811 37891 53839
rect 37488 53793 37909 53811
rect 37955 53793 38026 53839
rect 38123 53811 38143 53839
rect 38072 53793 38143 53811
rect 38189 53793 38261 53839
rect 38307 53793 38379 53839
rect 38425 53793 38497 53839
rect 38543 53793 38556 53839
rect 35294 53759 36266 53793
rect 36438 53768 36953 53793
rect 37439 53771 38161 53793
rect 37439 53768 37931 53771
rect 34228 53702 34718 53731
rect 33671 53656 33684 53702
rect 33730 53656 33787 53702
rect 33833 53656 33890 53702
rect 33936 53656 33993 53702
rect 34039 53656 34096 53702
rect 34142 53656 34199 53702
rect 34245 53691 34302 53702
rect 34245 53656 34267 53691
rect 34348 53656 34405 53702
rect 34451 53691 34508 53702
rect 34499 53656 34508 53691
rect 34554 53656 34612 53702
rect 34658 53691 34718 53702
rect 34228 53639 34267 53656
rect 34319 53639 34447 53656
rect 34499 53639 34627 53656
rect 34679 53639 34718 53691
rect 36438 53665 36554 53768
rect 34228 53598 34718 53639
rect 34964 53615 36360 53659
rect 30583 53413 31040 53490
rect 33019 53481 33327 53522
rect 33019 53478 33057 53481
rect 33109 53478 33237 53481
rect 33289 53478 33327 53481
rect 33484 53480 33552 53562
rect 34964 53569 35273 53615
rect 35523 53569 35580 53615
rect 35626 53569 35683 53615
rect 35729 53569 35786 53615
rect 35832 53569 35889 53615
rect 35935 53569 35992 53615
rect 36038 53569 36095 53615
rect 36141 53569 36198 53615
rect 36244 53569 36301 53615
rect 36347 53569 36360 53615
rect 34964 53537 36360 53569
rect 34964 53480 35082 53537
rect 31336 53432 31349 53478
rect 33323 53432 33336 53478
rect 33484 53443 35082 53480
rect 30583 53367 30637 53413
rect 30683 53373 31040 53413
rect 33019 53429 33057 53432
rect 33109 53429 33237 53432
rect 33289 53429 33327 53432
rect 33019 53389 33327 53429
rect 33484 53397 33816 53443
rect 33862 53397 34002 53443
rect 34048 53397 34189 53443
rect 34235 53397 34376 53443
rect 34422 53397 34562 53443
rect 34608 53397 35082 53443
rect 36438 53525 36475 53665
rect 36521 53525 36554 53665
rect 33484 53389 35082 53397
rect 35294 53391 36266 53431
rect 36438 53425 36554 53525
rect 36640 53665 36773 53688
rect 36640 53616 36697 53665
rect 36640 53564 36678 53616
rect 36640 53525 36697 53564
rect 36743 53525 36773 53665
rect 38658 53667 38726 53678
rect 36924 53657 37685 53663
rect 36923 53656 37685 53657
rect 36923 53623 37931 53656
rect 36923 53615 36961 53623
rect 37013 53615 37172 53623
rect 37224 53615 37384 53623
rect 36841 53569 36854 53615
rect 36900 53571 36961 53615
rect 36900 53569 36971 53571
rect 37017 53569 37088 53615
rect 37134 53571 37172 53615
rect 37134 53569 37206 53571
rect 37252 53569 37324 53615
rect 37370 53571 37384 53615
rect 37436 53615 37595 53623
rect 37436 53571 37442 53615
rect 37370 53569 37442 53571
rect 37488 53571 37595 53615
rect 37647 53615 37931 53623
rect 37647 53571 37909 53615
rect 37488 53569 37909 53571
rect 37955 53569 38026 53615
rect 38072 53569 38143 53615
rect 38189 53569 38261 53615
rect 38307 53569 38379 53615
rect 38425 53569 38497 53615
rect 38543 53569 38556 53615
rect 36923 53537 37931 53569
rect 36924 53530 37685 53537
rect 36640 53505 36773 53525
rect 38658 53527 38669 53667
rect 38715 53527 38726 53667
rect 39014 53615 39323 54101
rect 39492 54187 39608 54639
rect 39923 54606 40085 54737
rect 39923 54554 39994 54606
rect 40046 54554 40085 54606
rect 39923 54514 40085 54554
rect 39737 54418 39865 54431
rect 39737 54391 39866 54418
rect 39737 54374 39775 54391
rect 39827 54374 39866 54391
rect 39727 54328 39740 54374
rect 39827 54339 39862 54374
rect 39786 54328 39862 54339
rect 39908 54328 39985 54374
rect 40031 54328 40108 54374
rect 40154 54328 40167 54374
rect 40246 54363 40362 54761
rect 42229 54622 44509 54663
rect 42229 54570 42690 54622
rect 42742 54570 44509 54622
rect 42229 54530 44509 54570
rect 44341 54486 44509 54530
rect 44341 54440 44358 54486
rect 44498 54440 44509 54486
rect 39737 54299 39866 54328
rect 40246 54317 40281 54363
rect 40327 54317 40362 54363
rect 40246 54280 40362 54317
rect 40718 54391 43524 54432
rect 44341 54429 44509 54440
rect 40718 54339 41935 54391
rect 41987 54339 43524 54391
rect 40718 54298 43524 54339
rect 44605 54374 44721 54761
rect 45400 54731 48379 54772
rect 45400 54717 46731 54731
rect 45400 54671 45464 54717
rect 45604 54679 46731 54717
rect 46783 54679 48379 54731
rect 45604 54671 48379 54679
rect 44901 54615 45241 54656
rect 45400 54638 48379 54671
rect 48557 54725 48596 54777
rect 48648 54725 48687 54777
rect 48557 54702 48687 54725
rect 50044 54811 50516 54857
rect 50562 54811 50703 54857
rect 50749 54811 50890 54857
rect 50936 54811 51076 54857
rect 51122 54811 51263 54857
rect 51309 54811 51657 54857
rect 51797 54847 52105 54887
rect 51797 54822 51835 54847
rect 51887 54822 52015 54847
rect 52067 54822 52105 54847
rect 54085 54881 54223 54927
rect 54269 54887 54540 54927
rect 54269 54881 54440 54887
rect 54085 54841 54440 54881
rect 54486 54841 54540 54887
rect 50044 54774 51657 54811
rect 51789 54776 51802 54822
rect 53776 54776 53789 54822
rect 50044 54717 50160 54774
rect 44901 54598 44939 54615
rect 44991 54598 45151 54615
rect 45203 54598 45241 54615
rect 44799 54552 44812 54598
rect 44858 54552 44925 54598
rect 44991 54563 45038 54598
rect 44971 54552 45038 54563
rect 45084 54552 45151 54598
rect 45203 54563 45264 54598
rect 45197 54552 45264 54563
rect 45310 54552 45323 54598
rect 48557 54562 48622 54702
rect 48668 54562 48687 54702
rect 49820 54685 50160 54717
rect 48765 54639 48778 54685
rect 48824 54639 48881 54685
rect 48927 54639 48984 54685
rect 49030 54639 49087 54685
rect 49133 54639 49190 54685
rect 49236 54639 49293 54685
rect 49339 54639 49396 54685
rect 49442 54639 49499 54685
rect 49545 54639 49602 54685
rect 49852 54639 50160 54685
rect 51589 54722 51657 54774
rect 51797 54754 52105 54776
rect 49820 54598 50160 54639
rect 50262 54615 50812 54656
rect 48557 54559 48687 54562
rect 44901 54523 45241 54552
rect 48557 54507 48596 54559
rect 48648 54507 48687 54559
rect 50262 54563 50300 54615
rect 50352 54598 50511 54615
rect 50563 54598 50722 54615
rect 50352 54563 50467 54598
rect 50563 54563 50571 54598
rect 50262 54552 50467 54563
rect 50513 54552 50571 54563
rect 50617 54552 50674 54598
rect 50720 54563 50722 54598
rect 50774 54598 50812 54615
rect 50774 54563 50777 54598
rect 50720 54552 50777 54563
rect 50823 54552 50880 54598
rect 50926 54552 50983 54598
rect 51029 54552 51086 54598
rect 51132 54552 51189 54598
rect 51235 54552 51292 54598
rect 51338 54552 51395 54598
rect 51441 54552 51454 54598
rect 50262 54523 50812 54552
rect 48557 54466 48687 54507
rect 48905 54461 49877 54492
rect 48765 54415 48778 54461
rect 48824 54415 48881 54461
rect 48927 54452 48984 54461
rect 48927 54415 48943 54452
rect 49030 54415 49087 54461
rect 49133 54452 49190 54461
rect 49133 54415 49154 54452
rect 49236 54415 49293 54461
rect 49339 54452 49396 54461
rect 49339 54415 49365 54452
rect 49442 54415 49499 54461
rect 49545 54452 49602 54461
rect 49545 54415 49576 54452
rect 49852 54415 49877 54461
rect 48905 54400 48943 54415
rect 48995 54400 49154 54415
rect 49206 54400 49365 54415
rect 49417 54400 49576 54415
rect 49628 54400 49787 54415
rect 49839 54400 49877 54415
rect 44605 54328 44812 54374
rect 44858 54328 44925 54374
rect 44971 54328 45038 54374
rect 45084 54328 45151 54374
rect 45197 54328 45264 54374
rect 45310 54328 45323 54374
rect 48905 54360 49877 54400
rect 51035 54377 51343 54417
rect 51035 54374 51073 54377
rect 51125 54374 51253 54377
rect 51305 54374 51343 54377
rect 43362 54291 43524 54298
rect 43362 54245 43373 54291
rect 43513 54245 43524 54291
rect 43362 54234 43524 54245
rect 45584 54314 48546 54350
rect 50454 54328 50467 54374
rect 50513 54328 50571 54374
rect 50617 54328 50674 54374
rect 50720 54328 50777 54374
rect 50823 54328 50880 54374
rect 50926 54328 50983 54374
rect 51029 54328 51073 54374
rect 51132 54328 51189 54374
rect 51235 54328 51253 54374
rect 51338 54328 51395 54374
rect 51441 54328 51454 54374
rect 45584 54268 45619 54314
rect 45665 54268 45777 54314
rect 45823 54268 45935 54314
rect 45981 54268 46093 54314
rect 46139 54268 46251 54314
rect 46297 54268 46409 54314
rect 46455 54268 46568 54314
rect 46614 54268 46726 54314
rect 46772 54268 46884 54314
rect 46930 54268 47042 54314
rect 47088 54268 47200 54314
rect 47246 54268 47358 54314
rect 47404 54268 47516 54314
rect 47562 54268 47675 54314
rect 47721 54268 47833 54314
rect 47879 54268 47991 54314
rect 48037 54268 48149 54314
rect 48195 54268 48307 54314
rect 48353 54268 48465 54314
rect 48511 54268 48546 54314
rect 51035 54325 51073 54328
rect 51125 54325 51253 54328
rect 51305 54325 51343 54328
rect 51035 54284 51343 54325
rect 51589 54300 51600 54722
rect 51646 54300 51657 54722
rect 54085 54723 54540 54841
rect 54085 54677 54440 54723
rect 54486 54677 54540 54723
rect 54085 54649 54540 54677
rect 53585 54598 54540 54649
rect 51789 54552 51802 54598
rect 53776 54560 54540 54598
rect 53776 54552 54440 54560
rect 53585 54530 54440 54552
rect 54085 54514 54440 54530
rect 54486 54514 54540 54560
rect 54085 54438 54540 54514
rect 51797 54384 52105 54424
rect 51797 54374 51835 54384
rect 51887 54374 52015 54384
rect 52067 54374 52105 54384
rect 54085 54392 54223 54438
rect 54269 54397 54540 54438
rect 54269 54392 54440 54397
rect 51789 54328 51802 54374
rect 53776 54328 53789 54374
rect 54085 54351 54440 54392
rect 54486 54351 54540 54397
rect 51589 54289 51657 54300
rect 51797 54291 52105 54328
rect 40215 54187 40523 54194
rect 40788 54187 42986 54201
rect 43753 54187 44514 54194
rect 39492 54164 42986 54187
rect 43704 54164 44514 54187
rect 39492 54153 44514 54164
rect 39492 54150 40253 54153
rect 39492 54104 39740 54150
rect 39786 54104 39862 54150
rect 39908 54104 39985 54150
rect 40031 54104 40108 54150
rect 40154 54104 40253 54150
rect 39492 54101 40253 54104
rect 40305 54101 40433 54153
rect 40485 54150 43790 54153
rect 40485 54104 40836 54150
rect 40882 54104 40994 54150
rect 41040 54104 41152 54150
rect 41198 54104 41310 54150
rect 41356 54104 41469 54150
rect 41515 54104 41627 54150
rect 41673 54104 41785 54150
rect 41831 54104 41943 54150
rect 41989 54104 42101 54150
rect 42147 54104 42259 54150
rect 42305 54104 42418 54150
rect 42464 54104 42576 54150
rect 42622 54104 42734 54150
rect 42780 54104 42892 54150
rect 42938 54104 43739 54150
rect 43785 54104 43790 54150
rect 40485 54101 43790 54104
rect 43842 54150 44001 54153
rect 43842 54104 43906 54150
rect 43952 54104 44001 54150
rect 43842 54101 44001 54104
rect 44053 54150 44213 54153
rect 44265 54150 44424 54153
rect 44053 54104 44071 54150
rect 44117 54104 44213 54150
rect 44282 54104 44424 54150
rect 44053 54101 44213 54104
rect 44265 54101 44424 54104
rect 44476 54101 44514 54153
rect 39492 54090 44514 54101
rect 39492 54067 42986 54090
rect 43704 54067 44514 54090
rect 39492 53615 39608 54067
rect 40215 54060 40523 54067
rect 40788 54053 42986 54067
rect 43753 54060 44514 54067
rect 44796 54187 45346 54194
rect 45584 54187 48546 54268
rect 54085 54274 54540 54351
rect 54085 54228 54223 54274
rect 54269 54234 54540 54274
rect 54269 54228 54440 54234
rect 54085 54194 54440 54228
rect 48800 54187 49982 54194
rect 50308 54187 50859 54194
rect 44796 54153 49982 54187
rect 44796 54150 44834 54153
rect 44886 54150 45045 54153
rect 45097 54150 45256 54153
rect 45308 54150 48838 54153
rect 44796 54104 44812 54150
rect 44886 54104 44925 54150
rect 44971 54104 45038 54150
rect 45097 54104 45151 54150
rect 45197 54104 45256 54150
rect 45310 54104 45619 54150
rect 45665 54104 45777 54150
rect 45823 54104 45935 54150
rect 45981 54104 46093 54150
rect 46139 54104 46251 54150
rect 46297 54104 46409 54150
rect 46455 54104 46568 54150
rect 46614 54104 46726 54150
rect 46772 54104 46884 54150
rect 46930 54104 47042 54150
rect 47088 54104 47200 54150
rect 47246 54104 47358 54150
rect 47404 54104 47516 54150
rect 47562 54104 47675 54150
rect 47721 54104 47833 54150
rect 47879 54104 47991 54150
rect 48037 54104 48149 54150
rect 48195 54104 48307 54150
rect 48353 54104 48465 54150
rect 48511 54104 48838 54150
rect 44796 54101 44834 54104
rect 44886 54101 45045 54104
rect 45097 54101 45256 54104
rect 45308 54101 48838 54104
rect 48890 54101 49048 54153
rect 49100 54101 49259 54153
rect 49311 54101 49471 54153
rect 49523 54101 49682 54153
rect 49734 54101 49892 54153
rect 49944 54101 49982 54153
rect 44796 54067 49982 54101
rect 50307 54153 50859 54187
rect 50307 54101 50346 54153
rect 50398 54150 50557 54153
rect 50609 54150 50768 54153
rect 50820 54150 50859 54153
rect 52278 54188 54440 54194
rect 54486 54188 54540 54234
rect 55927 54887 57736 55001
rect 55927 54844 56267 54887
rect 55927 54798 55961 54844
rect 56007 54841 56267 54844
rect 56313 54841 57736 54887
rect 56007 54798 57736 54841
rect 55927 54723 57736 54798
rect 55927 54681 56267 54723
rect 55927 54635 55961 54681
rect 56007 54677 56267 54681
rect 56313 54677 57736 54723
rect 56007 54635 57736 54677
rect 55927 54560 57736 54635
rect 55927 54517 56267 54560
rect 55927 54471 55961 54517
rect 56007 54514 56267 54517
rect 56313 54514 57736 54560
rect 56007 54471 57736 54514
rect 55927 54397 57736 54471
rect 55927 54354 56267 54397
rect 55927 54308 55961 54354
rect 56007 54351 56267 54354
rect 56313 54351 57736 54397
rect 56007 54308 57736 54351
rect 55927 54234 57736 54308
rect 52278 54153 54540 54188
rect 52278 54150 52316 54153
rect 52368 54150 52527 54153
rect 52579 54150 52738 54153
rect 52790 54150 52948 54153
rect 53000 54150 53159 54153
rect 53211 54150 53371 54153
rect 53423 54150 53582 54153
rect 53634 54150 53792 54153
rect 50398 54104 50467 54150
rect 50513 54104 50557 54150
rect 50617 54104 50674 54150
rect 50720 54104 50768 54150
rect 50823 54104 50880 54150
rect 50926 54104 50983 54150
rect 51029 54104 51086 54150
rect 51132 54104 51189 54150
rect 51235 54104 51292 54150
rect 51338 54104 51395 54150
rect 51441 54104 51454 54150
rect 51789 54104 51802 54150
rect 53776 54104 53792 54150
rect 50398 54101 50557 54104
rect 50609 54101 50768 54104
rect 50820 54101 50859 54104
rect 50307 54067 50859 54101
rect 44796 54060 45346 54067
rect 43362 54009 43524 54020
rect 39737 53926 39866 53955
rect 40246 53937 40362 53974
rect 43362 53963 43373 54009
rect 43513 53963 43524 54009
rect 43362 53956 43524 53963
rect 39727 53880 39740 53926
rect 39786 53915 39862 53926
rect 39827 53880 39862 53915
rect 39908 53880 39985 53926
rect 40031 53880 40108 53926
rect 40154 53880 40167 53926
rect 40246 53891 40281 53937
rect 40327 53891 40362 53937
rect 39737 53863 39775 53880
rect 39827 53863 39866 53880
rect 39737 53836 39866 53863
rect 39737 53823 39865 53836
rect 39923 53700 40085 53740
rect 39923 53648 39994 53700
rect 40046 53648 40085 53700
rect 39008 53569 39021 53615
rect 39067 53569 39144 53615
rect 39190 53569 39267 53615
rect 39313 53569 39326 53615
rect 39492 53569 39641 53615
rect 39687 53569 39730 53615
rect 39014 53537 39323 53569
rect 39492 53537 39608 53569
rect 37853 53425 38161 53430
rect 36438 53391 36953 53425
rect 37439 53391 38161 53425
rect 38658 53405 38726 53527
rect 39923 53517 40085 53648
rect 39809 53514 40085 53517
rect 39809 53506 39994 53514
rect 39809 53460 39844 53506
rect 39890 53462 39994 53506
rect 40046 53493 40085 53514
rect 40246 53493 40362 53891
rect 40718 53915 43524 53956
rect 45584 53986 48546 54067
rect 48800 54060 49982 54067
rect 50308 54060 50859 54067
rect 52278 54101 52316 54104
rect 52368 54101 52527 54104
rect 52579 54101 52738 54104
rect 52790 54101 52948 54104
rect 53000 54101 53159 54104
rect 53211 54101 53371 54104
rect 53423 54101 53582 54104
rect 53634 54101 53792 54104
rect 53844 54101 54003 54153
rect 54055 54101 54214 54153
rect 54266 54101 54540 54153
rect 52278 54066 54540 54101
rect 52278 54060 54440 54066
rect 45584 53940 45619 53986
rect 45665 53940 45777 53986
rect 45823 53940 45935 53986
rect 45981 53940 46093 53986
rect 46139 53940 46251 53986
rect 46297 53940 46409 53986
rect 46455 53940 46568 53986
rect 46614 53940 46726 53986
rect 46772 53940 46884 53986
rect 46930 53940 47042 53986
rect 47088 53940 47200 53986
rect 47246 53940 47358 53986
rect 47404 53940 47516 53986
rect 47562 53940 47675 53986
rect 47721 53940 47833 53986
rect 47879 53940 47991 53986
rect 48037 53940 48149 53986
rect 48195 53940 48307 53986
rect 48353 53940 48465 53986
rect 48511 53940 48546 53986
rect 54085 54026 54440 54060
rect 54085 53980 54223 54026
rect 54269 54020 54440 54026
rect 54486 54020 54540 54066
rect 54758 54153 55840 54194
rect 54758 54150 54855 54153
rect 54758 54104 54793 54150
rect 54839 54104 54855 54150
rect 54758 54101 54855 54104
rect 54907 54150 55066 54153
rect 54907 54104 54956 54150
rect 55002 54104 55066 54150
rect 54907 54101 55066 54104
rect 55118 54150 55278 54153
rect 55330 54150 55489 54153
rect 55164 54104 55278 54150
rect 55330 54104 55439 54150
rect 55485 54104 55489 54150
rect 55118 54101 55278 54104
rect 55330 54101 55489 54104
rect 55541 54150 55840 54153
rect 55541 54104 55599 54150
rect 55645 54104 55760 54150
rect 55806 54104 55840 54150
rect 55541 54101 55840 54104
rect 54758 54061 55840 54101
rect 55927 54188 56267 54234
rect 56313 54188 57736 54234
rect 55927 54066 57736 54188
rect 54817 54060 55579 54061
rect 54269 53980 54540 54020
rect 40718 53863 41935 53915
rect 41987 53863 43524 53915
rect 40718 53822 43524 53863
rect 44605 53880 44812 53926
rect 44858 53880 44925 53926
rect 44971 53880 45038 53926
rect 45084 53880 45151 53926
rect 45197 53880 45264 53926
rect 45310 53880 45323 53926
rect 45584 53904 48546 53940
rect 51035 53929 51343 53970
rect 51035 53926 51073 53929
rect 51125 53926 51253 53929
rect 51305 53926 51343 53929
rect 51589 53954 51657 53965
rect 44341 53814 44509 53825
rect 44341 53768 44358 53814
rect 44498 53768 44509 53814
rect 44341 53724 44509 53768
rect 42229 53684 44509 53724
rect 42229 53632 42690 53684
rect 42742 53632 44509 53684
rect 42229 53591 44509 53632
rect 44605 53493 44721 53880
rect 48905 53854 49877 53894
rect 50454 53880 50467 53926
rect 50513 53880 50571 53926
rect 50617 53880 50674 53926
rect 50720 53880 50777 53926
rect 50823 53880 50880 53926
rect 50926 53880 50983 53926
rect 51029 53880 51073 53926
rect 51132 53880 51189 53926
rect 51235 53880 51253 53926
rect 51338 53880 51395 53926
rect 51441 53880 51454 53926
rect 48905 53839 48943 53854
rect 48995 53839 49154 53854
rect 49206 53839 49365 53854
rect 49417 53839 49576 53854
rect 49628 53839 49787 53854
rect 49839 53839 49877 53854
rect 48765 53793 48778 53839
rect 48824 53793 48881 53839
rect 48927 53802 48943 53839
rect 48927 53793 48984 53802
rect 49030 53793 49087 53839
rect 49133 53802 49154 53839
rect 49133 53793 49190 53802
rect 49236 53793 49293 53839
rect 49339 53802 49365 53839
rect 49339 53793 49396 53802
rect 49442 53793 49499 53839
rect 49545 53802 49576 53839
rect 49545 53793 49602 53802
rect 49852 53793 49877 53839
rect 51035 53877 51073 53880
rect 51125 53877 51253 53880
rect 51305 53877 51343 53880
rect 51035 53837 51343 53877
rect 48557 53747 48687 53788
rect 48905 53762 49877 53793
rect 44901 53702 45241 53731
rect 44799 53656 44812 53702
rect 44858 53656 44925 53702
rect 44971 53691 45038 53702
rect 44991 53656 45038 53691
rect 45084 53656 45151 53702
rect 45197 53691 45264 53702
rect 45203 53656 45264 53691
rect 45310 53656 45323 53702
rect 48557 53695 48596 53747
rect 48648 53695 48687 53747
rect 48557 53692 48687 53695
rect 44901 53639 44939 53656
rect 44991 53639 45151 53656
rect 45203 53639 45241 53656
rect 44901 53598 45241 53639
rect 45400 53583 48379 53616
rect 45400 53537 45464 53583
rect 45604 53575 48379 53583
rect 45604 53537 47108 53575
rect 45400 53523 47108 53537
rect 47160 53523 48379 53575
rect 40046 53478 44918 53493
rect 45400 53482 48379 53523
rect 48557 53552 48622 53692
rect 48668 53552 48687 53692
rect 50262 53702 50812 53731
rect 50262 53691 50467 53702
rect 50513 53691 50571 53702
rect 49820 53615 50160 53656
rect 48765 53569 48778 53615
rect 48824 53569 48881 53615
rect 48927 53569 48984 53615
rect 49030 53569 49087 53615
rect 49133 53569 49190 53615
rect 49236 53569 49293 53615
rect 49339 53569 49396 53615
rect 49442 53569 49499 53615
rect 49545 53569 49602 53615
rect 49852 53569 50160 53615
rect 50262 53639 50300 53691
rect 50352 53656 50467 53691
rect 50563 53656 50571 53691
rect 50617 53656 50674 53702
rect 50720 53691 50777 53702
rect 50720 53656 50722 53691
rect 50352 53639 50511 53656
rect 50563 53639 50722 53656
rect 50774 53656 50777 53691
rect 50823 53656 50880 53702
rect 50926 53656 50983 53702
rect 51029 53656 51086 53702
rect 51132 53656 51189 53702
rect 51235 53656 51292 53702
rect 51338 53656 51395 53702
rect 51441 53656 51454 53702
rect 50774 53639 50812 53656
rect 50262 53598 50812 53639
rect 48557 53529 48687 53552
rect 49820 53537 50160 53569
rect 40046 53462 44812 53478
rect 39890 53460 44812 53462
rect 39809 53457 44812 53460
rect 39809 53411 43739 53457
rect 43785 53411 43906 53457
rect 43952 53411 44071 53457
rect 44117 53411 44236 53457
rect 44282 53432 44812 53457
rect 44858 53432 44925 53478
rect 44971 53432 45038 53478
rect 45084 53432 45151 53478
rect 45197 53432 45264 53478
rect 45310 53432 45323 53478
rect 48557 53477 48596 53529
rect 48648 53477 48687 53529
rect 48557 53437 48687 53477
rect 50044 53480 50160 53537
rect 51589 53532 51600 53954
rect 51646 53532 51657 53954
rect 51797 53926 52105 53963
rect 51789 53880 51802 53926
rect 53776 53880 53789 53926
rect 54085 53903 54540 53980
rect 51797 53870 51835 53880
rect 51887 53870 52015 53880
rect 52067 53870 52105 53880
rect 51797 53830 52105 53870
rect 54085 53862 54440 53903
rect 54085 53816 54223 53862
rect 54269 53857 54440 53862
rect 54486 53857 54540 53903
rect 54269 53816 54540 53857
rect 54085 53740 54540 53816
rect 54085 53724 54440 53740
rect 53585 53702 54440 53724
rect 51789 53656 51802 53702
rect 53776 53694 54440 53702
rect 54486 53694 54540 53740
rect 53776 53656 54540 53694
rect 53585 53605 54540 53656
rect 51589 53480 51657 53532
rect 54085 53577 54540 53605
rect 54085 53531 54440 53577
rect 54486 53531 54540 53577
rect 50044 53443 51657 53480
rect 51797 53478 52105 53500
rect 44282 53411 44918 53432
rect 38658 53391 39723 53405
rect 30683 53367 30855 53373
rect 30583 53327 30855 53367
rect 30901 53327 31040 53373
rect 33484 53360 34643 53389
rect 35260 53345 35273 53391
rect 35523 53345 35543 53391
rect 35626 53345 35683 53391
rect 35729 53345 35754 53391
rect 35832 53345 35889 53391
rect 35935 53345 35965 53391
rect 36038 53345 36095 53391
rect 36141 53345 36176 53391
rect 36244 53345 36301 53391
rect 36347 53345 36360 53391
rect 36438 53345 36854 53391
rect 36900 53345 36971 53391
rect 37017 53345 37088 53391
rect 37134 53345 37206 53391
rect 37252 53345 37324 53391
rect 37370 53345 37442 53391
rect 37488 53389 37909 53391
rect 37488 53345 37891 53389
rect 37955 53345 38026 53391
rect 38072 53389 38143 53391
rect 38123 53345 38143 53389
rect 38189 53345 38261 53391
rect 38307 53345 38379 53391
rect 38425 53345 38497 53391
rect 38543 53345 38556 53391
rect 38658 53345 39021 53391
rect 39067 53345 39144 53391
rect 39190 53345 39267 53391
rect 39313 53345 39641 53391
rect 39687 53345 39730 53391
rect 39809 53373 44918 53411
rect 48905 53391 49877 53431
rect 48765 53345 48778 53391
rect 48824 53345 48881 53391
rect 48927 53345 48943 53391
rect 49030 53345 49087 53391
rect 49133 53345 49154 53391
rect 49236 53345 49293 53391
rect 49339 53345 49365 53391
rect 49442 53345 49499 53391
rect 49545 53345 49576 53391
rect 49852 53345 49877 53391
rect 50044 53397 50516 53443
rect 50562 53397 50703 53443
rect 50749 53397 50890 53443
rect 50936 53397 51076 53443
rect 51122 53397 51263 53443
rect 51309 53397 51657 53443
rect 51789 53432 51802 53478
rect 53776 53432 53789 53478
rect 50044 53387 51657 53397
rect 50481 53360 51657 53387
rect 51797 53407 51835 53432
rect 51887 53407 52015 53432
rect 52067 53407 52105 53432
rect 51797 53367 52105 53407
rect 54085 53413 54540 53531
rect 54085 53373 54440 53413
rect 30583 53294 31040 53327
rect 35294 53339 35332 53345
rect 35384 53339 35543 53345
rect 35595 53339 35754 53345
rect 35806 53339 35965 53345
rect 36017 53339 36176 53345
rect 36228 53339 36266 53345
rect 34870 53294 35025 53301
rect 35294 53299 36266 53339
rect 36438 53305 36953 53345
rect 37439 53337 37891 53345
rect 37943 53337 38071 53345
rect 38123 53337 38161 53345
rect 37439 53305 38161 53337
rect 37853 53297 38161 53305
rect 27387 53201 27790 53253
rect 27842 53201 28001 53253
rect 28053 53201 28212 53253
rect 28264 53201 28423 53253
rect 28475 53201 28634 53253
rect 28686 53250 28845 53253
rect 28686 53204 28810 53250
rect 28686 53201 28845 53204
rect 28897 53201 29056 53253
rect 29108 53201 29196 53253
rect 27387 53087 29196 53201
rect 29283 53253 30365 53294
rect 29283 53250 29582 53253
rect 29283 53204 29317 53250
rect 29363 53204 29478 53250
rect 29524 53204 29582 53250
rect 29283 53201 29582 53204
rect 29634 53250 29793 53253
rect 29845 53250 30005 53253
rect 29634 53204 29638 53250
rect 29684 53204 29793 53250
rect 29845 53204 29959 53250
rect 29634 53201 29793 53204
rect 29845 53201 30005 53204
rect 30057 53250 30216 53253
rect 30057 53204 30121 53250
rect 30167 53204 30216 53250
rect 30057 53201 30216 53204
rect 30268 53250 30365 53253
rect 30268 53204 30284 53250
rect 30330 53204 30365 53250
rect 30268 53201 30365 53204
rect 29283 53161 30365 53201
rect 30583 53253 32842 53294
rect 30583 53250 30854 53253
rect 30583 53204 30637 53250
rect 30683 53204 30854 53250
rect 30583 53201 30854 53204
rect 30906 53201 31065 53253
rect 31117 53201 31276 53253
rect 31328 53201 31486 53253
rect 31538 53201 31697 53253
rect 31749 53201 31909 53253
rect 31961 53201 32120 53253
rect 32172 53201 32330 53253
rect 32382 53201 32541 53253
rect 32593 53201 32752 53253
rect 32804 53201 32842 53253
rect 29544 53160 30306 53161
rect 30583 53160 32842 53201
rect 34717 53253 35025 53294
rect 38658 53285 39723 53345
rect 48905 53339 48943 53345
rect 48995 53339 49154 53345
rect 49206 53339 49365 53345
rect 49417 53339 49576 53345
rect 49628 53339 49787 53345
rect 49839 53339 49877 53345
rect 48905 53299 49877 53339
rect 54085 53327 54223 53373
rect 54269 53367 54440 53373
rect 54486 53367 54540 53413
rect 54269 53327 54540 53367
rect 50099 53294 50255 53301
rect 54085 53294 54540 53327
rect 55927 54020 56267 54066
rect 56313 54020 57736 54066
rect 55927 53944 57736 54020
rect 55927 53898 55961 53944
rect 56007 53903 57736 53944
rect 56007 53898 56267 53903
rect 55927 53857 56267 53898
rect 56313 53857 57736 53903
rect 55927 53781 57736 53857
rect 55927 53735 55961 53781
rect 56007 53740 57736 53781
rect 56007 53735 56267 53740
rect 55927 53694 56267 53735
rect 56313 53694 57736 53740
rect 55927 53617 57736 53694
rect 55927 53571 55961 53617
rect 56007 53577 57736 53617
rect 56007 53571 56267 53577
rect 55927 53531 56267 53571
rect 56313 53531 57736 53577
rect 55927 53454 57736 53531
rect 55927 53408 55961 53454
rect 56007 53413 57736 53454
rect 56007 53408 56267 53413
rect 55927 53367 56267 53408
rect 56313 53367 57736 53413
rect 34717 53201 34755 53253
rect 34807 53250 34935 53253
rect 34807 53204 34916 53250
rect 34807 53201 34935 53204
rect 34987 53201 35025 53253
rect 34717 53160 35025 53201
rect 50099 53253 50408 53294
rect 50099 53201 50138 53253
rect 50190 53250 50318 53253
rect 50206 53204 50318 53250
rect 50190 53201 50318 53204
rect 50370 53201 50408 53253
rect 27387 53041 28810 53087
rect 28856 53044 29196 53087
rect 28856 53041 29116 53044
rect 27387 52998 29116 53041
rect 29162 52998 29196 53044
rect 27387 52923 29196 52998
rect 27387 52877 28810 52923
rect 28856 52881 29196 52923
rect 28856 52877 29116 52881
rect 27387 52835 29116 52877
rect 29162 52835 29196 52881
rect 27387 52760 29196 52835
rect 27387 52714 28810 52760
rect 28856 52717 29196 52760
rect 28856 52714 29116 52717
rect 27387 52671 29116 52714
rect 29162 52671 29196 52717
rect 27387 52597 29196 52671
rect 27387 52551 28810 52597
rect 28856 52554 29196 52597
rect 28856 52551 29116 52554
rect 27387 52508 29116 52551
rect 29162 52508 29196 52554
rect 27387 52434 29196 52508
rect 27387 52388 28810 52434
rect 28856 52388 29196 52434
rect 30583 53127 31040 53160
rect 34870 53153 35025 53160
rect 30583 53087 30855 53127
rect 30583 53041 30637 53087
rect 30683 53081 30855 53087
rect 30901 53081 31040 53127
rect 35294 53115 36266 53155
rect 37853 53149 38161 53157
rect 35294 53109 35332 53115
rect 35384 53109 35543 53115
rect 35595 53109 35754 53115
rect 35806 53109 35965 53115
rect 36017 53109 36176 53115
rect 36228 53109 36266 53115
rect 36438 53109 36953 53149
rect 37439 53117 38161 53149
rect 37439 53109 37891 53117
rect 37943 53109 38071 53117
rect 38123 53109 38161 53117
rect 38658 53109 39723 53169
rect 50099 53160 50408 53201
rect 52278 53253 54540 53294
rect 52278 53201 52316 53253
rect 52368 53201 52527 53253
rect 52579 53201 52738 53253
rect 52790 53201 52948 53253
rect 53000 53201 53159 53253
rect 53211 53201 53371 53253
rect 53423 53201 53582 53253
rect 53634 53201 53792 53253
rect 53844 53201 54003 53253
rect 54055 53201 54214 53253
rect 54266 53250 54540 53253
rect 54266 53204 54440 53250
rect 54486 53204 54540 53250
rect 54266 53201 54540 53204
rect 52278 53160 54540 53201
rect 54758 53253 55840 53294
rect 54758 53250 54855 53253
rect 54758 53204 54793 53250
rect 54839 53204 54855 53250
rect 54758 53201 54855 53204
rect 54907 53250 55066 53253
rect 54907 53204 54956 53250
rect 55002 53204 55066 53250
rect 54907 53201 55066 53204
rect 55118 53250 55278 53253
rect 55330 53250 55489 53253
rect 55164 53204 55278 53250
rect 55330 53204 55439 53250
rect 55485 53204 55489 53250
rect 55118 53201 55278 53204
rect 55330 53201 55489 53204
rect 55541 53250 55840 53253
rect 55541 53204 55599 53250
rect 55645 53204 55760 53250
rect 55806 53204 55840 53250
rect 55541 53201 55840 53204
rect 54758 53161 55840 53201
rect 55927 53253 57736 53367
rect 55927 53201 56015 53253
rect 56067 53201 56226 53253
rect 56278 53250 56437 53253
rect 56313 53204 56437 53250
rect 56278 53201 56437 53204
rect 56489 53201 56648 53253
rect 56700 53201 56859 53253
rect 56911 53201 57070 53253
rect 57122 53201 57281 53253
rect 57333 53201 57736 53253
rect 54817 53160 55579 53161
rect 48905 53115 49877 53155
rect 50099 53153 50255 53160
rect 48905 53109 48943 53115
rect 48995 53109 49154 53115
rect 49206 53109 49365 53115
rect 49417 53109 49576 53115
rect 49628 53109 49787 53115
rect 49839 53109 49877 53115
rect 30683 53041 31040 53081
rect 33484 53065 34643 53094
rect 30583 52964 31040 53041
rect 33019 53025 33327 53065
rect 33019 53022 33057 53025
rect 33109 53022 33237 53025
rect 33289 53022 33327 53025
rect 33484 53057 35082 53065
rect 35260 53063 35273 53109
rect 35523 53063 35543 53109
rect 35626 53063 35683 53109
rect 35729 53063 35754 53109
rect 35832 53063 35889 53109
rect 35935 53063 35965 53109
rect 36038 53063 36095 53109
rect 36141 53063 36176 53109
rect 36244 53063 36301 53109
rect 36347 53063 36360 53109
rect 36438 53063 36854 53109
rect 36900 53063 36971 53109
rect 37017 53063 37088 53109
rect 37134 53063 37206 53109
rect 37252 53063 37324 53109
rect 37370 53063 37442 53109
rect 37488 53065 37891 53109
rect 37488 53063 37909 53065
rect 37955 53063 38026 53109
rect 38123 53065 38143 53109
rect 38072 53063 38143 53065
rect 38189 53063 38261 53109
rect 38307 53063 38379 53109
rect 38425 53063 38497 53109
rect 38543 53063 38556 53109
rect 38658 53063 39021 53109
rect 39067 53063 39144 53109
rect 39190 53063 39267 53109
rect 39313 53063 39641 53109
rect 39687 53063 39730 53109
rect 31336 52976 31349 53022
rect 33323 52976 33336 53022
rect 33484 53011 33816 53057
rect 33862 53011 34002 53057
rect 34048 53011 34189 53057
rect 34235 53011 34376 53057
rect 34422 53011 34562 53057
rect 34608 53011 35082 53057
rect 35294 53023 36266 53063
rect 36438 53029 36953 53063
rect 37439 53029 38161 53063
rect 30583 52923 30855 52964
rect 30583 52877 30637 52923
rect 30683 52918 30855 52923
rect 30901 52918 31040 52964
rect 33019 52973 33057 52976
rect 33109 52973 33237 52976
rect 33289 52973 33327 52976
rect 33019 52932 33327 52973
rect 33484 52974 35082 53011
rect 30683 52877 31040 52918
rect 30583 52849 31040 52877
rect 33484 52892 33552 52974
rect 30583 52801 31493 52849
rect 30583 52760 30855 52801
rect 30583 52714 30637 52760
rect 30683 52755 30855 52760
rect 30901 52798 31493 52801
rect 30901 52755 31349 52798
rect 30683 52752 31349 52755
rect 33323 52752 33336 52798
rect 30683 52730 31493 52752
rect 30683 52714 31040 52730
rect 30583 52638 31040 52714
rect 30583 52597 30855 52638
rect 30583 52551 30637 52597
rect 30683 52592 30855 52597
rect 30901 52592 31040 52638
rect 30683 52551 31040 52592
rect 33019 52577 33327 52617
rect 33019 52574 33057 52577
rect 33109 52574 33237 52577
rect 33289 52574 33327 52577
rect 30583 52474 31040 52551
rect 31336 52528 31349 52574
rect 33323 52528 33336 52574
rect 33019 52525 33057 52528
rect 33109 52525 33237 52528
rect 33289 52525 33327 52528
rect 33019 52484 33327 52525
rect 30583 52434 30855 52474
rect 27387 52266 29196 52388
rect 27387 52220 28810 52266
rect 28856 52220 29196 52266
rect 29283 52353 30365 52394
rect 29283 52350 29582 52353
rect 29283 52304 29317 52350
rect 29363 52304 29478 52350
rect 29524 52304 29582 52350
rect 29283 52301 29582 52304
rect 29634 52350 29793 52353
rect 29845 52350 30005 52353
rect 29634 52304 29638 52350
rect 29684 52304 29793 52350
rect 29845 52304 29959 52350
rect 29634 52301 29793 52304
rect 29845 52301 30005 52304
rect 30057 52350 30216 52353
rect 30057 52304 30121 52350
rect 30167 52304 30216 52350
rect 30057 52301 30216 52304
rect 30268 52350 30365 52353
rect 30268 52304 30284 52350
rect 30330 52304 30365 52350
rect 30268 52301 30365 52304
rect 29283 52261 30365 52301
rect 30583 52388 30637 52434
rect 30683 52428 30855 52434
rect 30901 52428 31040 52474
rect 33484 52470 33495 52892
rect 33541 52470 33552 52892
rect 34964 52917 35082 52974
rect 36438 52929 36554 53029
rect 37853 53024 38161 53029
rect 38658 53049 39723 53063
rect 34964 52885 36360 52917
rect 34228 52815 34718 52856
rect 34228 52798 34267 52815
rect 34319 52798 34447 52815
rect 34499 52798 34627 52815
rect 33671 52752 33684 52798
rect 33730 52752 33787 52798
rect 33833 52752 33890 52798
rect 33936 52752 33993 52798
rect 34039 52752 34096 52798
rect 34142 52752 34199 52798
rect 34245 52763 34267 52798
rect 34245 52752 34302 52763
rect 34348 52752 34405 52798
rect 34499 52763 34508 52798
rect 34451 52752 34508 52763
rect 34554 52752 34612 52798
rect 34679 52763 34718 52815
rect 34964 52839 35273 52885
rect 35523 52839 35580 52885
rect 35626 52839 35683 52885
rect 35729 52839 35786 52885
rect 35832 52839 35889 52885
rect 35935 52839 35992 52885
rect 36038 52839 36095 52885
rect 36141 52839 36198 52885
rect 36244 52839 36301 52885
rect 36347 52839 36360 52885
rect 34964 52795 36360 52839
rect 34658 52752 34718 52763
rect 34228 52723 34718 52752
rect 36438 52789 36475 52929
rect 36521 52789 36554 52929
rect 35294 52661 36266 52695
rect 36438 52686 36554 52789
rect 36640 52929 36773 52949
rect 36640 52890 36697 52929
rect 36640 52838 36678 52890
rect 36640 52789 36697 52838
rect 36743 52789 36773 52929
rect 38658 52927 38726 53049
rect 39809 53043 44918 53081
rect 48765 53063 48778 53109
rect 48824 53063 48881 53109
rect 48927 53063 48943 53109
rect 49030 53063 49087 53109
rect 49133 53063 49154 53109
rect 49236 53063 49293 53109
rect 49339 53063 49365 53109
rect 49442 53063 49499 53109
rect 49545 53063 49576 53109
rect 49852 53063 49877 53109
rect 54085 53127 54540 53160
rect 50481 53067 51657 53094
rect 39809 52997 43739 53043
rect 43785 52997 43906 53043
rect 43952 52997 44071 53043
rect 44117 52997 44236 53043
rect 44282 53022 44918 53043
rect 48905 53023 49877 53063
rect 50044 53057 51657 53067
rect 44282 52997 44812 53022
rect 39809 52994 44812 52997
rect 39809 52948 39844 52994
rect 39890 52992 44812 52994
rect 39890 52948 39994 52992
rect 39809 52940 39994 52948
rect 40046 52976 44812 52992
rect 44858 52976 44925 53022
rect 44971 52976 45038 53022
rect 45084 52976 45151 53022
rect 45197 52976 45264 53022
rect 45310 52976 45323 53022
rect 48557 52977 48687 53017
rect 40046 52961 44918 52976
rect 40046 52940 40085 52961
rect 39809 52937 40085 52940
rect 36924 52917 37685 52924
rect 36923 52885 37931 52917
rect 36841 52839 36854 52885
rect 36900 52883 36971 52885
rect 36900 52839 36961 52883
rect 37017 52839 37088 52885
rect 37134 52883 37206 52885
rect 37134 52839 37172 52883
rect 37252 52839 37324 52885
rect 37370 52883 37442 52885
rect 37370 52839 37384 52883
rect 36923 52831 36961 52839
rect 37013 52831 37172 52839
rect 37224 52831 37384 52839
rect 37436 52839 37442 52883
rect 37488 52883 37909 52885
rect 37488 52839 37595 52883
rect 37436 52831 37595 52839
rect 37647 52839 37909 52883
rect 37955 52839 38026 52885
rect 38072 52839 38143 52885
rect 38189 52839 38261 52885
rect 38307 52839 38379 52885
rect 38425 52839 38497 52885
rect 38543 52839 38556 52885
rect 37647 52831 37931 52839
rect 36923 52798 37931 52831
rect 36923 52797 37685 52798
rect 36924 52791 37685 52797
rect 36640 52766 36773 52789
rect 38658 52787 38669 52927
rect 38715 52787 38726 52927
rect 39014 52885 39323 52917
rect 39492 52885 39608 52917
rect 39008 52839 39021 52885
rect 39067 52839 39144 52885
rect 39190 52839 39267 52885
rect 39313 52839 39326 52885
rect 39492 52839 39641 52885
rect 39687 52839 39730 52885
rect 38658 52776 38726 52787
rect 36438 52661 36953 52686
rect 37439 52683 37931 52686
rect 37439 52661 38161 52683
rect 35260 52615 35273 52661
rect 35523 52655 35580 52661
rect 35523 52615 35543 52655
rect 35626 52615 35683 52661
rect 35729 52655 35786 52661
rect 35729 52615 35754 52655
rect 35832 52615 35889 52661
rect 35935 52655 35992 52661
rect 35935 52615 35965 52655
rect 36038 52615 36095 52661
rect 36141 52655 36198 52661
rect 36141 52615 36176 52655
rect 36244 52615 36301 52661
rect 36347 52615 36360 52661
rect 36438 52615 36854 52661
rect 36900 52615 36971 52661
rect 37017 52615 37088 52661
rect 37134 52615 37206 52661
rect 37252 52615 37324 52661
rect 37370 52615 37442 52661
rect 37488 52643 37909 52661
rect 37488 52615 37891 52643
rect 37955 52615 38026 52661
rect 38072 52643 38143 52661
rect 38123 52615 38143 52643
rect 38189 52615 38261 52661
rect 38307 52615 38379 52661
rect 38425 52615 38497 52661
rect 38543 52615 38556 52661
rect 33781 52574 34089 52609
rect 35294 52603 35332 52615
rect 35384 52603 35543 52615
rect 35595 52603 35754 52615
rect 35806 52603 35965 52615
rect 36017 52603 36176 52615
rect 36228 52603 36266 52615
rect 33671 52528 33684 52574
rect 33730 52528 33787 52574
rect 33833 52569 33890 52574
rect 33871 52528 33890 52569
rect 33936 52528 33993 52574
rect 34039 52569 34096 52574
rect 34051 52528 34096 52569
rect 34142 52528 34199 52574
rect 34245 52528 34302 52574
rect 34348 52528 34405 52574
rect 34451 52528 34508 52574
rect 34554 52528 34612 52574
rect 34658 52528 34671 52574
rect 35294 52563 36266 52603
rect 36438 52566 36953 52615
rect 37439 52591 37891 52615
rect 37943 52591 38071 52615
rect 38123 52591 38161 52615
rect 37439 52566 38161 52591
rect 37853 52550 38161 52566
rect 33781 52517 33819 52528
rect 33871 52517 33999 52528
rect 34051 52517 34089 52528
rect 33781 52476 34089 52517
rect 33484 52459 33552 52470
rect 30683 52394 31040 52428
rect 30683 52388 32842 52394
rect 30583 52353 32842 52388
rect 34247 52387 35008 52394
rect 30583 52301 30854 52353
rect 30906 52301 31065 52353
rect 31117 52301 31276 52353
rect 31328 52350 31486 52353
rect 31538 52350 31697 52353
rect 31749 52350 31909 52353
rect 31961 52350 32120 52353
rect 32172 52350 32330 52353
rect 32382 52350 32541 52353
rect 32593 52350 32752 52353
rect 32804 52350 32842 52353
rect 34246 52353 35008 52387
rect 34246 52350 34284 52353
rect 34336 52350 34495 52353
rect 34547 52350 34707 52353
rect 31328 52304 31349 52350
rect 33323 52304 33336 52350
rect 33671 52304 33684 52350
rect 33730 52304 33787 52350
rect 33833 52304 33890 52350
rect 33936 52304 33993 52350
rect 34039 52304 34096 52350
rect 34142 52304 34199 52350
rect 34245 52304 34284 52350
rect 34348 52304 34405 52350
rect 34451 52304 34495 52350
rect 34554 52304 34612 52350
rect 34658 52304 34707 52350
rect 31328 52301 31486 52304
rect 31538 52301 31697 52304
rect 31749 52301 31909 52304
rect 31961 52301 32120 52304
rect 32172 52301 32330 52304
rect 32382 52301 32541 52304
rect 32593 52301 32752 52304
rect 32804 52301 32842 52304
rect 30583 52266 32842 52301
rect 34246 52301 34284 52304
rect 34336 52301 34495 52304
rect 34547 52301 34707 52304
rect 34759 52301 34918 52353
rect 34970 52301 35008 52353
rect 34246 52267 35008 52301
rect 29544 52260 30306 52261
rect 27387 52144 29196 52220
rect 27387 52103 29116 52144
rect 27387 52057 28810 52103
rect 28856 52098 29116 52103
rect 29162 52098 29196 52144
rect 28856 52057 29196 52098
rect 27387 51981 29196 52057
rect 27387 51940 29116 51981
rect 27387 51894 28810 51940
rect 28856 51935 29116 51940
rect 29162 51935 29196 51981
rect 28856 51894 29196 51935
rect 27387 51817 29196 51894
rect 27387 51777 29116 51817
rect 27387 51731 28810 51777
rect 28856 51771 29116 51777
rect 29162 51771 29196 51817
rect 28856 51731 29196 51771
rect 27387 51654 29196 51731
rect 27387 51613 29116 51654
rect 27387 51567 28810 51613
rect 28856 51608 29116 51613
rect 29162 51608 29196 51654
rect 28856 51567 29196 51608
rect 27387 51453 29196 51567
rect 30583 52220 30637 52266
rect 30683 52260 32842 52266
rect 34247 52260 35008 52267
rect 35182 52387 36364 52394
rect 35182 52353 36958 52387
rect 35182 52301 35220 52353
rect 35272 52301 35430 52353
rect 35482 52301 35641 52353
rect 35693 52301 35853 52353
rect 35905 52301 36064 52353
rect 36116 52301 36274 52353
rect 36326 52350 36958 52353
rect 36326 52304 36489 52350
rect 36723 52304 36958 52350
rect 36326 52301 36958 52304
rect 35182 52267 36958 52301
rect 37946 52353 38842 52394
rect 37946 52350 38330 52353
rect 38382 52350 38541 52353
rect 37946 52304 37957 52350
rect 38473 52304 38541 52350
rect 37946 52301 38330 52304
rect 38382 52301 38541 52304
rect 38593 52301 38752 52353
rect 38804 52301 38842 52353
rect 35182 52260 36364 52267
rect 37946 52260 38842 52301
rect 39014 52353 39323 52839
rect 39014 52301 39052 52353
rect 39104 52350 39232 52353
rect 39108 52304 39220 52350
rect 39104 52301 39232 52304
rect 39284 52301 39323 52353
rect 30683 52226 31040 52260
rect 30683 52220 30855 52226
rect 30583 52180 30855 52220
rect 30901 52180 31040 52226
rect 30583 52103 31040 52180
rect 33484 52184 33552 52195
rect 33019 52129 33327 52170
rect 33019 52126 33057 52129
rect 33109 52126 33237 52129
rect 33289 52126 33327 52129
rect 30583 52057 30637 52103
rect 30683 52062 31040 52103
rect 31336 52080 31349 52126
rect 33323 52080 33336 52126
rect 30683 52057 30855 52062
rect 30583 52016 30855 52057
rect 30901 52016 31040 52062
rect 33019 52077 33057 52080
rect 33109 52077 33237 52080
rect 33289 52077 33327 52080
rect 33019 52037 33327 52077
rect 30583 51940 31040 52016
rect 30583 51894 30637 51940
rect 30683 51924 31040 51940
rect 30683 51902 31493 51924
rect 30683 51899 31349 51902
rect 30683 51894 30855 51899
rect 30583 51853 30855 51894
rect 30901 51856 31349 51899
rect 33323 51856 33336 51902
rect 30901 51853 31493 51856
rect 30583 51805 31493 51853
rect 30583 51777 31040 51805
rect 30583 51731 30637 51777
rect 30683 51736 31040 51777
rect 30683 51731 30855 51736
rect 30583 51690 30855 51731
rect 30901 51690 31040 51736
rect 33484 51762 33495 52184
rect 33541 51762 33552 52184
rect 33781 52137 34089 52178
rect 33781 52126 33819 52137
rect 33871 52126 33999 52137
rect 34051 52126 34089 52137
rect 33671 52080 33684 52126
rect 33730 52080 33787 52126
rect 33871 52085 33890 52126
rect 33833 52080 33890 52085
rect 33936 52080 33993 52126
rect 34051 52085 34096 52126
rect 34039 52080 34096 52085
rect 34142 52080 34199 52126
rect 34245 52080 34302 52126
rect 34348 52080 34405 52126
rect 34451 52080 34508 52126
rect 34554 52080 34612 52126
rect 34658 52080 34671 52126
rect 33781 52045 34089 52080
rect 35294 52051 36266 52091
rect 37853 52088 38161 52104
rect 35294 52039 35332 52051
rect 35384 52039 35543 52051
rect 35595 52039 35754 52051
rect 35806 52039 35965 52051
rect 36017 52039 36176 52051
rect 36228 52039 36266 52051
rect 36438 52039 36953 52088
rect 37439 52063 38161 52088
rect 37439 52039 37891 52063
rect 37943 52039 38071 52063
rect 38123 52039 38161 52063
rect 35260 51993 35273 52039
rect 35523 51999 35543 52039
rect 35523 51993 35580 51999
rect 35626 51993 35683 52039
rect 35729 51999 35754 52039
rect 35729 51993 35786 51999
rect 35832 51993 35889 52039
rect 35935 51999 35965 52039
rect 35935 51993 35992 51999
rect 36038 51993 36095 52039
rect 36141 51999 36176 52039
rect 36141 51993 36198 51999
rect 36244 51993 36301 52039
rect 36347 51993 36360 52039
rect 36438 51993 36854 52039
rect 36900 51993 36971 52039
rect 37017 51993 37088 52039
rect 37134 51993 37206 52039
rect 37252 51993 37324 52039
rect 37370 51993 37442 52039
rect 37488 52011 37891 52039
rect 37488 51993 37909 52011
rect 37955 51993 38026 52039
rect 38123 52011 38143 52039
rect 38072 51993 38143 52011
rect 38189 51993 38261 52039
rect 38307 51993 38379 52039
rect 38425 51993 38497 52039
rect 38543 51993 38556 52039
rect 35294 51959 36266 51993
rect 36438 51968 36953 51993
rect 37439 51971 38161 51993
rect 37439 51968 37931 51971
rect 34228 51902 34718 51931
rect 33671 51856 33684 51902
rect 33730 51856 33787 51902
rect 33833 51856 33890 51902
rect 33936 51856 33993 51902
rect 34039 51856 34096 51902
rect 34142 51856 34199 51902
rect 34245 51891 34302 51902
rect 34245 51856 34267 51891
rect 34348 51856 34405 51902
rect 34451 51891 34508 51902
rect 34499 51856 34508 51891
rect 34554 51856 34612 51902
rect 34658 51891 34718 51902
rect 34228 51839 34267 51856
rect 34319 51839 34447 51856
rect 34499 51839 34627 51856
rect 34679 51839 34718 51891
rect 36438 51865 36554 51968
rect 34228 51798 34718 51839
rect 34964 51815 36360 51859
rect 30583 51613 31040 51690
rect 33019 51681 33327 51722
rect 33019 51678 33057 51681
rect 33109 51678 33237 51681
rect 33289 51678 33327 51681
rect 33484 51680 33552 51762
rect 34964 51769 35273 51815
rect 35523 51769 35580 51815
rect 35626 51769 35683 51815
rect 35729 51769 35786 51815
rect 35832 51769 35889 51815
rect 35935 51769 35992 51815
rect 36038 51769 36095 51815
rect 36141 51769 36198 51815
rect 36244 51769 36301 51815
rect 36347 51769 36360 51815
rect 34964 51737 36360 51769
rect 34964 51680 35082 51737
rect 31336 51632 31349 51678
rect 33323 51632 33336 51678
rect 33484 51643 35082 51680
rect 30583 51567 30637 51613
rect 30683 51573 31040 51613
rect 33019 51629 33057 51632
rect 33109 51629 33237 51632
rect 33289 51629 33327 51632
rect 33019 51589 33327 51629
rect 33484 51597 33816 51643
rect 33862 51597 34002 51643
rect 34048 51597 34189 51643
rect 34235 51597 34376 51643
rect 34422 51597 34562 51643
rect 34608 51597 35082 51643
rect 36438 51725 36475 51865
rect 36521 51725 36554 51865
rect 33484 51589 35082 51597
rect 35294 51591 36266 51631
rect 36438 51625 36554 51725
rect 36640 51865 36773 51888
rect 36640 51816 36697 51865
rect 36640 51764 36678 51816
rect 36640 51725 36697 51764
rect 36743 51725 36773 51865
rect 38658 51867 38726 51878
rect 36924 51857 37685 51863
rect 36923 51856 37685 51857
rect 36923 51823 37931 51856
rect 36923 51815 36961 51823
rect 37013 51815 37172 51823
rect 37224 51815 37384 51823
rect 36841 51769 36854 51815
rect 36900 51771 36961 51815
rect 36900 51769 36971 51771
rect 37017 51769 37088 51815
rect 37134 51771 37172 51815
rect 37134 51769 37206 51771
rect 37252 51769 37324 51815
rect 37370 51771 37384 51815
rect 37436 51815 37595 51823
rect 37436 51771 37442 51815
rect 37370 51769 37442 51771
rect 37488 51771 37595 51815
rect 37647 51815 37931 51823
rect 37647 51771 37909 51815
rect 37488 51769 37909 51771
rect 37955 51769 38026 51815
rect 38072 51769 38143 51815
rect 38189 51769 38261 51815
rect 38307 51769 38379 51815
rect 38425 51769 38497 51815
rect 38543 51769 38556 51815
rect 36923 51737 37931 51769
rect 36924 51730 37685 51737
rect 36640 51705 36773 51725
rect 38658 51727 38669 51867
rect 38715 51727 38726 51867
rect 39014 51815 39323 52301
rect 39492 52387 39608 52839
rect 39923 52806 40085 52937
rect 39923 52754 39994 52806
rect 40046 52754 40085 52806
rect 39923 52714 40085 52754
rect 39737 52618 39865 52631
rect 39737 52591 39866 52618
rect 39737 52574 39775 52591
rect 39827 52574 39866 52591
rect 39727 52528 39740 52574
rect 39827 52539 39862 52574
rect 39786 52528 39862 52539
rect 39908 52528 39985 52574
rect 40031 52528 40108 52574
rect 40154 52528 40167 52574
rect 40246 52563 40362 52961
rect 42229 52822 44509 52863
rect 42229 52770 42690 52822
rect 42742 52770 44509 52822
rect 42229 52730 44509 52770
rect 44341 52686 44509 52730
rect 44341 52640 44358 52686
rect 44498 52640 44509 52686
rect 39737 52499 39866 52528
rect 40246 52517 40281 52563
rect 40327 52517 40362 52563
rect 40246 52480 40362 52517
rect 40718 52591 43524 52632
rect 44341 52629 44509 52640
rect 40718 52539 41935 52591
rect 41987 52539 43524 52591
rect 40718 52498 43524 52539
rect 44605 52574 44721 52961
rect 45400 52931 48379 52972
rect 45400 52917 47486 52931
rect 45400 52871 45464 52917
rect 45604 52879 47486 52917
rect 47538 52879 48379 52931
rect 45604 52871 48379 52879
rect 44901 52815 45241 52856
rect 45400 52838 48379 52871
rect 48557 52925 48596 52977
rect 48648 52925 48687 52977
rect 48557 52902 48687 52925
rect 50044 53011 50516 53057
rect 50562 53011 50703 53057
rect 50749 53011 50890 53057
rect 50936 53011 51076 53057
rect 51122 53011 51263 53057
rect 51309 53011 51657 53057
rect 51797 53047 52105 53087
rect 51797 53022 51835 53047
rect 51887 53022 52015 53047
rect 52067 53022 52105 53047
rect 54085 53081 54223 53127
rect 54269 53087 54540 53127
rect 54269 53081 54440 53087
rect 54085 53041 54440 53081
rect 54486 53041 54540 53087
rect 50044 52974 51657 53011
rect 51789 52976 51802 53022
rect 53776 52976 53789 53022
rect 50044 52917 50160 52974
rect 44901 52798 44939 52815
rect 44991 52798 45151 52815
rect 45203 52798 45241 52815
rect 44799 52752 44812 52798
rect 44858 52752 44925 52798
rect 44991 52763 45038 52798
rect 44971 52752 45038 52763
rect 45084 52752 45151 52798
rect 45203 52763 45264 52798
rect 45197 52752 45264 52763
rect 45310 52752 45323 52798
rect 48557 52762 48622 52902
rect 48668 52762 48687 52902
rect 49820 52885 50160 52917
rect 48765 52839 48778 52885
rect 48824 52839 48881 52885
rect 48927 52839 48984 52885
rect 49030 52839 49087 52885
rect 49133 52839 49190 52885
rect 49236 52839 49293 52885
rect 49339 52839 49396 52885
rect 49442 52839 49499 52885
rect 49545 52839 49602 52885
rect 49852 52839 50160 52885
rect 51589 52922 51657 52974
rect 51797 52954 52105 52976
rect 49820 52798 50160 52839
rect 50262 52815 50812 52856
rect 48557 52759 48687 52762
rect 44901 52723 45241 52752
rect 48557 52707 48596 52759
rect 48648 52707 48687 52759
rect 50262 52763 50300 52815
rect 50352 52798 50511 52815
rect 50563 52798 50722 52815
rect 50352 52763 50467 52798
rect 50563 52763 50571 52798
rect 50262 52752 50467 52763
rect 50513 52752 50571 52763
rect 50617 52752 50674 52798
rect 50720 52763 50722 52798
rect 50774 52798 50812 52815
rect 50774 52763 50777 52798
rect 50720 52752 50777 52763
rect 50823 52752 50880 52798
rect 50926 52752 50983 52798
rect 51029 52752 51086 52798
rect 51132 52752 51189 52798
rect 51235 52752 51292 52798
rect 51338 52752 51395 52798
rect 51441 52752 51454 52798
rect 50262 52723 50812 52752
rect 48557 52666 48687 52707
rect 48905 52661 49877 52692
rect 48765 52615 48778 52661
rect 48824 52615 48881 52661
rect 48927 52652 48984 52661
rect 48927 52615 48943 52652
rect 49030 52615 49087 52661
rect 49133 52652 49190 52661
rect 49133 52615 49154 52652
rect 49236 52615 49293 52661
rect 49339 52652 49396 52661
rect 49339 52615 49365 52652
rect 49442 52615 49499 52661
rect 49545 52652 49602 52661
rect 49545 52615 49576 52652
rect 49852 52615 49877 52661
rect 48905 52600 48943 52615
rect 48995 52600 49154 52615
rect 49206 52600 49365 52615
rect 49417 52600 49576 52615
rect 49628 52600 49787 52615
rect 49839 52600 49877 52615
rect 44605 52528 44812 52574
rect 44858 52528 44925 52574
rect 44971 52528 45038 52574
rect 45084 52528 45151 52574
rect 45197 52528 45264 52574
rect 45310 52528 45323 52574
rect 48905 52560 49877 52600
rect 51035 52577 51343 52617
rect 51035 52574 51073 52577
rect 51125 52574 51253 52577
rect 51305 52574 51343 52577
rect 43362 52491 43524 52498
rect 43362 52445 43373 52491
rect 43513 52445 43524 52491
rect 43362 52434 43524 52445
rect 45584 52514 48546 52550
rect 50454 52528 50467 52574
rect 50513 52528 50571 52574
rect 50617 52528 50674 52574
rect 50720 52528 50777 52574
rect 50823 52528 50880 52574
rect 50926 52528 50983 52574
rect 51029 52528 51073 52574
rect 51132 52528 51189 52574
rect 51235 52528 51253 52574
rect 51338 52528 51395 52574
rect 51441 52528 51454 52574
rect 45584 52468 45619 52514
rect 45665 52468 45777 52514
rect 45823 52468 45935 52514
rect 45981 52468 46093 52514
rect 46139 52468 46251 52514
rect 46297 52468 46409 52514
rect 46455 52468 46568 52514
rect 46614 52468 46726 52514
rect 46772 52468 46884 52514
rect 46930 52468 47042 52514
rect 47088 52468 47200 52514
rect 47246 52468 47358 52514
rect 47404 52468 47516 52514
rect 47562 52468 47675 52514
rect 47721 52468 47833 52514
rect 47879 52468 47991 52514
rect 48037 52468 48149 52514
rect 48195 52468 48307 52514
rect 48353 52468 48465 52514
rect 48511 52468 48546 52514
rect 51035 52525 51073 52528
rect 51125 52525 51253 52528
rect 51305 52525 51343 52528
rect 51035 52484 51343 52525
rect 51589 52500 51600 52922
rect 51646 52500 51657 52922
rect 54085 52923 54540 53041
rect 54085 52877 54440 52923
rect 54486 52877 54540 52923
rect 54085 52849 54540 52877
rect 53585 52798 54540 52849
rect 51789 52752 51802 52798
rect 53776 52760 54540 52798
rect 53776 52752 54440 52760
rect 53585 52730 54440 52752
rect 54085 52714 54440 52730
rect 54486 52714 54540 52760
rect 54085 52638 54540 52714
rect 51797 52584 52105 52624
rect 51797 52574 51835 52584
rect 51887 52574 52015 52584
rect 52067 52574 52105 52584
rect 54085 52592 54223 52638
rect 54269 52597 54540 52638
rect 54269 52592 54440 52597
rect 51789 52528 51802 52574
rect 53776 52528 53789 52574
rect 54085 52551 54440 52592
rect 54486 52551 54540 52597
rect 51589 52489 51657 52500
rect 51797 52491 52105 52528
rect 40215 52387 40523 52394
rect 40788 52387 42986 52401
rect 43753 52387 44514 52394
rect 39492 52364 42986 52387
rect 43704 52364 44514 52387
rect 39492 52353 44514 52364
rect 39492 52350 40253 52353
rect 39492 52304 39740 52350
rect 39786 52304 39862 52350
rect 39908 52304 39985 52350
rect 40031 52304 40108 52350
rect 40154 52304 40253 52350
rect 39492 52301 40253 52304
rect 40305 52301 40433 52353
rect 40485 52350 43790 52353
rect 40485 52304 40836 52350
rect 40882 52304 40994 52350
rect 41040 52304 41152 52350
rect 41198 52304 41310 52350
rect 41356 52304 41469 52350
rect 41515 52304 41627 52350
rect 41673 52304 41785 52350
rect 41831 52304 41943 52350
rect 41989 52304 42101 52350
rect 42147 52304 42259 52350
rect 42305 52304 42418 52350
rect 42464 52304 42576 52350
rect 42622 52304 42734 52350
rect 42780 52304 42892 52350
rect 42938 52304 43739 52350
rect 43785 52304 43790 52350
rect 40485 52301 43790 52304
rect 43842 52350 44001 52353
rect 43842 52304 43906 52350
rect 43952 52304 44001 52350
rect 43842 52301 44001 52304
rect 44053 52350 44213 52353
rect 44265 52350 44424 52353
rect 44053 52304 44071 52350
rect 44117 52304 44213 52350
rect 44282 52304 44424 52350
rect 44053 52301 44213 52304
rect 44265 52301 44424 52304
rect 44476 52301 44514 52353
rect 39492 52290 44514 52301
rect 39492 52267 42986 52290
rect 43704 52267 44514 52290
rect 39492 51815 39608 52267
rect 40215 52260 40523 52267
rect 40788 52253 42986 52267
rect 43753 52260 44514 52267
rect 44796 52387 45346 52394
rect 45584 52387 48546 52468
rect 54085 52474 54540 52551
rect 54085 52428 54223 52474
rect 54269 52434 54540 52474
rect 54269 52428 54440 52434
rect 54085 52394 54440 52428
rect 48800 52387 49982 52394
rect 50308 52387 50859 52394
rect 44796 52353 49982 52387
rect 44796 52350 44834 52353
rect 44886 52350 45045 52353
rect 45097 52350 45256 52353
rect 45308 52350 48838 52353
rect 44796 52304 44812 52350
rect 44886 52304 44925 52350
rect 44971 52304 45038 52350
rect 45097 52304 45151 52350
rect 45197 52304 45256 52350
rect 45310 52304 45619 52350
rect 45665 52304 45777 52350
rect 45823 52304 45935 52350
rect 45981 52304 46093 52350
rect 46139 52304 46251 52350
rect 46297 52304 46409 52350
rect 46455 52304 46568 52350
rect 46614 52304 46726 52350
rect 46772 52304 46884 52350
rect 46930 52304 47042 52350
rect 47088 52304 47200 52350
rect 47246 52304 47358 52350
rect 47404 52304 47516 52350
rect 47562 52304 47675 52350
rect 47721 52304 47833 52350
rect 47879 52304 47991 52350
rect 48037 52304 48149 52350
rect 48195 52304 48307 52350
rect 48353 52304 48465 52350
rect 48511 52304 48838 52350
rect 44796 52301 44834 52304
rect 44886 52301 45045 52304
rect 45097 52301 45256 52304
rect 45308 52301 48838 52304
rect 48890 52301 49048 52353
rect 49100 52301 49259 52353
rect 49311 52301 49471 52353
rect 49523 52301 49682 52353
rect 49734 52301 49892 52353
rect 49944 52301 49982 52353
rect 44796 52267 49982 52301
rect 50307 52353 50859 52387
rect 50307 52301 50346 52353
rect 50398 52350 50557 52353
rect 50609 52350 50768 52353
rect 50820 52350 50859 52353
rect 52278 52388 54440 52394
rect 54486 52388 54540 52434
rect 55927 53087 57736 53201
rect 55927 53044 56267 53087
rect 55927 52998 55961 53044
rect 56007 53041 56267 53044
rect 56313 53041 57736 53087
rect 56007 52998 57736 53041
rect 55927 52923 57736 52998
rect 55927 52881 56267 52923
rect 55927 52835 55961 52881
rect 56007 52877 56267 52881
rect 56313 52877 57736 52923
rect 56007 52835 57736 52877
rect 55927 52760 57736 52835
rect 55927 52717 56267 52760
rect 55927 52671 55961 52717
rect 56007 52714 56267 52717
rect 56313 52714 57736 52760
rect 56007 52671 57736 52714
rect 55927 52597 57736 52671
rect 55927 52554 56267 52597
rect 55927 52508 55961 52554
rect 56007 52551 56267 52554
rect 56313 52551 57736 52597
rect 56007 52508 57736 52551
rect 55927 52434 57736 52508
rect 52278 52353 54540 52388
rect 52278 52350 52316 52353
rect 52368 52350 52527 52353
rect 52579 52350 52738 52353
rect 52790 52350 52948 52353
rect 53000 52350 53159 52353
rect 53211 52350 53371 52353
rect 53423 52350 53582 52353
rect 53634 52350 53792 52353
rect 50398 52304 50467 52350
rect 50513 52304 50557 52350
rect 50617 52304 50674 52350
rect 50720 52304 50768 52350
rect 50823 52304 50880 52350
rect 50926 52304 50983 52350
rect 51029 52304 51086 52350
rect 51132 52304 51189 52350
rect 51235 52304 51292 52350
rect 51338 52304 51395 52350
rect 51441 52304 51454 52350
rect 51789 52304 51802 52350
rect 53776 52304 53792 52350
rect 50398 52301 50557 52304
rect 50609 52301 50768 52304
rect 50820 52301 50859 52304
rect 50307 52267 50859 52301
rect 44796 52260 45346 52267
rect 43362 52209 43524 52220
rect 39737 52126 39866 52155
rect 40246 52137 40362 52174
rect 43362 52163 43373 52209
rect 43513 52163 43524 52209
rect 43362 52156 43524 52163
rect 39727 52080 39740 52126
rect 39786 52115 39862 52126
rect 39827 52080 39862 52115
rect 39908 52080 39985 52126
rect 40031 52080 40108 52126
rect 40154 52080 40167 52126
rect 40246 52091 40281 52137
rect 40327 52091 40362 52137
rect 39737 52063 39775 52080
rect 39827 52063 39866 52080
rect 39737 52036 39866 52063
rect 39737 52023 39865 52036
rect 39923 51900 40085 51940
rect 39923 51848 39994 51900
rect 40046 51848 40085 51900
rect 39008 51769 39021 51815
rect 39067 51769 39144 51815
rect 39190 51769 39267 51815
rect 39313 51769 39326 51815
rect 39492 51769 39641 51815
rect 39687 51769 39730 51815
rect 39014 51737 39323 51769
rect 39492 51737 39608 51769
rect 37853 51625 38161 51630
rect 36438 51591 36953 51625
rect 37439 51591 38161 51625
rect 38658 51605 38726 51727
rect 39923 51717 40085 51848
rect 39809 51714 40085 51717
rect 39809 51706 39994 51714
rect 39809 51660 39844 51706
rect 39890 51662 39994 51706
rect 40046 51693 40085 51714
rect 40246 51693 40362 52091
rect 40718 52115 43524 52156
rect 45584 52186 48546 52267
rect 48800 52260 49982 52267
rect 50308 52260 50859 52267
rect 52278 52301 52316 52304
rect 52368 52301 52527 52304
rect 52579 52301 52738 52304
rect 52790 52301 52948 52304
rect 53000 52301 53159 52304
rect 53211 52301 53371 52304
rect 53423 52301 53582 52304
rect 53634 52301 53792 52304
rect 53844 52301 54003 52353
rect 54055 52301 54214 52353
rect 54266 52301 54540 52353
rect 52278 52266 54540 52301
rect 52278 52260 54440 52266
rect 45584 52140 45619 52186
rect 45665 52140 45777 52186
rect 45823 52140 45935 52186
rect 45981 52140 46093 52186
rect 46139 52140 46251 52186
rect 46297 52140 46409 52186
rect 46455 52140 46568 52186
rect 46614 52140 46726 52186
rect 46772 52140 46884 52186
rect 46930 52140 47042 52186
rect 47088 52140 47200 52186
rect 47246 52140 47358 52186
rect 47404 52140 47516 52186
rect 47562 52140 47675 52186
rect 47721 52140 47833 52186
rect 47879 52140 47991 52186
rect 48037 52140 48149 52186
rect 48195 52140 48307 52186
rect 48353 52140 48465 52186
rect 48511 52140 48546 52186
rect 54085 52226 54440 52260
rect 54085 52180 54223 52226
rect 54269 52220 54440 52226
rect 54486 52220 54540 52266
rect 54758 52353 55840 52394
rect 54758 52350 54855 52353
rect 54758 52304 54793 52350
rect 54839 52304 54855 52350
rect 54758 52301 54855 52304
rect 54907 52350 55066 52353
rect 54907 52304 54956 52350
rect 55002 52304 55066 52350
rect 54907 52301 55066 52304
rect 55118 52350 55278 52353
rect 55330 52350 55489 52353
rect 55164 52304 55278 52350
rect 55330 52304 55439 52350
rect 55485 52304 55489 52350
rect 55118 52301 55278 52304
rect 55330 52301 55489 52304
rect 55541 52350 55840 52353
rect 55541 52304 55599 52350
rect 55645 52304 55760 52350
rect 55806 52304 55840 52350
rect 55541 52301 55840 52304
rect 54758 52261 55840 52301
rect 55927 52388 56267 52434
rect 56313 52388 57736 52434
rect 55927 52266 57736 52388
rect 54817 52260 55579 52261
rect 54269 52180 54540 52220
rect 40718 52063 41935 52115
rect 41987 52063 43524 52115
rect 40718 52022 43524 52063
rect 44605 52080 44812 52126
rect 44858 52080 44925 52126
rect 44971 52080 45038 52126
rect 45084 52080 45151 52126
rect 45197 52080 45264 52126
rect 45310 52080 45323 52126
rect 45584 52104 48546 52140
rect 51035 52129 51343 52170
rect 51035 52126 51073 52129
rect 51125 52126 51253 52129
rect 51305 52126 51343 52129
rect 51589 52154 51657 52165
rect 44341 52014 44509 52025
rect 44341 51968 44358 52014
rect 44498 51968 44509 52014
rect 44341 51924 44509 51968
rect 42229 51884 44509 51924
rect 42229 51832 42690 51884
rect 42742 51832 44509 51884
rect 42229 51791 44509 51832
rect 44605 51693 44721 52080
rect 48905 52054 49877 52094
rect 50454 52080 50467 52126
rect 50513 52080 50571 52126
rect 50617 52080 50674 52126
rect 50720 52080 50777 52126
rect 50823 52080 50880 52126
rect 50926 52080 50983 52126
rect 51029 52080 51073 52126
rect 51132 52080 51189 52126
rect 51235 52080 51253 52126
rect 51338 52080 51395 52126
rect 51441 52080 51454 52126
rect 48905 52039 48943 52054
rect 48995 52039 49154 52054
rect 49206 52039 49365 52054
rect 49417 52039 49576 52054
rect 49628 52039 49787 52054
rect 49839 52039 49877 52054
rect 48765 51993 48778 52039
rect 48824 51993 48881 52039
rect 48927 52002 48943 52039
rect 48927 51993 48984 52002
rect 49030 51993 49087 52039
rect 49133 52002 49154 52039
rect 49133 51993 49190 52002
rect 49236 51993 49293 52039
rect 49339 52002 49365 52039
rect 49339 51993 49396 52002
rect 49442 51993 49499 52039
rect 49545 52002 49576 52039
rect 49545 51993 49602 52002
rect 49852 51993 49877 52039
rect 51035 52077 51073 52080
rect 51125 52077 51253 52080
rect 51305 52077 51343 52080
rect 51035 52037 51343 52077
rect 48557 51947 48687 51988
rect 48905 51962 49877 51993
rect 44901 51902 45241 51931
rect 44799 51856 44812 51902
rect 44858 51856 44925 51902
rect 44971 51891 45038 51902
rect 44991 51856 45038 51891
rect 45084 51856 45151 51902
rect 45197 51891 45264 51902
rect 45203 51856 45264 51891
rect 45310 51856 45323 51902
rect 48557 51895 48596 51947
rect 48648 51895 48687 51947
rect 48557 51892 48687 51895
rect 44901 51839 44939 51856
rect 44991 51839 45151 51856
rect 45203 51839 45241 51856
rect 44901 51798 45241 51839
rect 45400 51783 48379 51816
rect 45400 51737 45464 51783
rect 45604 51775 48379 51783
rect 45604 51737 47864 51775
rect 45400 51723 47864 51737
rect 47916 51723 48379 51775
rect 40046 51678 44918 51693
rect 45400 51682 48379 51723
rect 48557 51752 48622 51892
rect 48668 51752 48687 51892
rect 50262 51902 50812 51931
rect 50262 51891 50467 51902
rect 50513 51891 50571 51902
rect 49820 51815 50160 51856
rect 48765 51769 48778 51815
rect 48824 51769 48881 51815
rect 48927 51769 48984 51815
rect 49030 51769 49087 51815
rect 49133 51769 49190 51815
rect 49236 51769 49293 51815
rect 49339 51769 49396 51815
rect 49442 51769 49499 51815
rect 49545 51769 49602 51815
rect 49852 51769 50160 51815
rect 50262 51839 50300 51891
rect 50352 51856 50467 51891
rect 50563 51856 50571 51891
rect 50617 51856 50674 51902
rect 50720 51891 50777 51902
rect 50720 51856 50722 51891
rect 50352 51839 50511 51856
rect 50563 51839 50722 51856
rect 50774 51856 50777 51891
rect 50823 51856 50880 51902
rect 50926 51856 50983 51902
rect 51029 51856 51086 51902
rect 51132 51856 51189 51902
rect 51235 51856 51292 51902
rect 51338 51856 51395 51902
rect 51441 51856 51454 51902
rect 50774 51839 50812 51856
rect 50262 51798 50812 51839
rect 48557 51729 48687 51752
rect 49820 51737 50160 51769
rect 40046 51662 44812 51678
rect 39890 51660 44812 51662
rect 39809 51657 44812 51660
rect 39809 51611 43739 51657
rect 43785 51611 43906 51657
rect 43952 51611 44071 51657
rect 44117 51611 44236 51657
rect 44282 51632 44812 51657
rect 44858 51632 44925 51678
rect 44971 51632 45038 51678
rect 45084 51632 45151 51678
rect 45197 51632 45264 51678
rect 45310 51632 45323 51678
rect 48557 51677 48596 51729
rect 48648 51677 48687 51729
rect 48557 51637 48687 51677
rect 50044 51680 50160 51737
rect 51589 51732 51600 52154
rect 51646 51732 51657 52154
rect 51797 52126 52105 52163
rect 51789 52080 51802 52126
rect 53776 52080 53789 52126
rect 54085 52103 54540 52180
rect 51797 52070 51835 52080
rect 51887 52070 52015 52080
rect 52067 52070 52105 52080
rect 51797 52030 52105 52070
rect 54085 52062 54440 52103
rect 54085 52016 54223 52062
rect 54269 52057 54440 52062
rect 54486 52057 54540 52103
rect 54269 52016 54540 52057
rect 54085 51940 54540 52016
rect 54085 51924 54440 51940
rect 53585 51902 54440 51924
rect 51789 51856 51802 51902
rect 53776 51894 54440 51902
rect 54486 51894 54540 51940
rect 53776 51856 54540 51894
rect 53585 51805 54540 51856
rect 51589 51680 51657 51732
rect 54085 51777 54540 51805
rect 54085 51731 54440 51777
rect 54486 51731 54540 51777
rect 50044 51643 51657 51680
rect 51797 51678 52105 51700
rect 44282 51611 44918 51632
rect 38658 51591 39723 51605
rect 30683 51567 30855 51573
rect 30583 51527 30855 51567
rect 30901 51527 31040 51573
rect 33484 51560 34643 51589
rect 35260 51545 35273 51591
rect 35523 51545 35543 51591
rect 35626 51545 35683 51591
rect 35729 51545 35754 51591
rect 35832 51545 35889 51591
rect 35935 51545 35965 51591
rect 36038 51545 36095 51591
rect 36141 51545 36176 51591
rect 36244 51545 36301 51591
rect 36347 51545 36360 51591
rect 36438 51545 36854 51591
rect 36900 51545 36971 51591
rect 37017 51545 37088 51591
rect 37134 51545 37206 51591
rect 37252 51545 37324 51591
rect 37370 51545 37442 51591
rect 37488 51589 37909 51591
rect 37488 51545 37891 51589
rect 37955 51545 38026 51591
rect 38072 51589 38143 51591
rect 38123 51545 38143 51589
rect 38189 51545 38261 51591
rect 38307 51545 38379 51591
rect 38425 51545 38497 51591
rect 38543 51545 38556 51591
rect 38658 51545 39021 51591
rect 39067 51545 39144 51591
rect 39190 51545 39267 51591
rect 39313 51545 39641 51591
rect 39687 51545 39730 51591
rect 39809 51573 44918 51611
rect 48905 51591 49877 51631
rect 48765 51545 48778 51591
rect 48824 51545 48881 51591
rect 48927 51545 48943 51591
rect 49030 51545 49087 51591
rect 49133 51545 49154 51591
rect 49236 51545 49293 51591
rect 49339 51545 49365 51591
rect 49442 51545 49499 51591
rect 49545 51545 49576 51591
rect 49852 51545 49877 51591
rect 50044 51597 50516 51643
rect 50562 51597 50703 51643
rect 50749 51597 50890 51643
rect 50936 51597 51076 51643
rect 51122 51597 51263 51643
rect 51309 51597 51657 51643
rect 51789 51632 51802 51678
rect 53776 51632 53789 51678
rect 50044 51587 51657 51597
rect 50481 51560 51657 51587
rect 51797 51607 51835 51632
rect 51887 51607 52015 51632
rect 52067 51607 52105 51632
rect 51797 51567 52105 51607
rect 54085 51613 54540 51731
rect 54085 51573 54440 51613
rect 30583 51494 31040 51527
rect 35294 51539 35332 51545
rect 35384 51539 35543 51545
rect 35595 51539 35754 51545
rect 35806 51539 35965 51545
rect 36017 51539 36176 51545
rect 36228 51539 36266 51545
rect 34870 51494 35025 51501
rect 35294 51499 36266 51539
rect 36438 51505 36953 51545
rect 37439 51537 37891 51545
rect 37943 51537 38071 51545
rect 38123 51537 38161 51545
rect 37439 51505 38161 51537
rect 37853 51497 38161 51505
rect 27387 51401 27790 51453
rect 27842 51401 28001 51453
rect 28053 51401 28212 51453
rect 28264 51401 28423 51453
rect 28475 51401 28634 51453
rect 28686 51450 28845 51453
rect 28686 51404 28810 51450
rect 28686 51401 28845 51404
rect 28897 51401 29056 51453
rect 29108 51401 29196 51453
rect 27387 51287 29196 51401
rect 29283 51453 30365 51494
rect 29283 51450 29582 51453
rect 29283 51404 29317 51450
rect 29363 51404 29478 51450
rect 29524 51404 29582 51450
rect 29283 51401 29582 51404
rect 29634 51450 29793 51453
rect 29845 51450 30005 51453
rect 29634 51404 29638 51450
rect 29684 51404 29793 51450
rect 29845 51404 29959 51450
rect 29634 51401 29793 51404
rect 29845 51401 30005 51404
rect 30057 51450 30216 51453
rect 30057 51404 30121 51450
rect 30167 51404 30216 51450
rect 30057 51401 30216 51404
rect 30268 51450 30365 51453
rect 30268 51404 30284 51450
rect 30330 51404 30365 51450
rect 30268 51401 30365 51404
rect 29283 51361 30365 51401
rect 30583 51453 32842 51494
rect 30583 51450 30854 51453
rect 30583 51404 30637 51450
rect 30683 51404 30854 51450
rect 30583 51401 30854 51404
rect 30906 51401 31065 51453
rect 31117 51401 31276 51453
rect 31328 51401 31486 51453
rect 31538 51401 31697 51453
rect 31749 51401 31909 51453
rect 31961 51401 32120 51453
rect 32172 51401 32330 51453
rect 32382 51401 32541 51453
rect 32593 51401 32752 51453
rect 32804 51401 32842 51453
rect 29544 51360 30306 51361
rect 30583 51360 32842 51401
rect 34717 51453 35025 51494
rect 38658 51485 39723 51545
rect 48905 51539 48943 51545
rect 48995 51539 49154 51545
rect 49206 51539 49365 51545
rect 49417 51539 49576 51545
rect 49628 51539 49787 51545
rect 49839 51539 49877 51545
rect 48905 51499 49877 51539
rect 54085 51527 54223 51573
rect 54269 51567 54440 51573
rect 54486 51567 54540 51613
rect 54269 51527 54540 51567
rect 50099 51494 50255 51501
rect 54085 51494 54540 51527
rect 55927 52220 56267 52266
rect 56313 52220 57736 52266
rect 55927 52144 57736 52220
rect 55927 52098 55961 52144
rect 56007 52103 57736 52144
rect 56007 52098 56267 52103
rect 55927 52057 56267 52098
rect 56313 52057 57736 52103
rect 55927 51981 57736 52057
rect 55927 51935 55961 51981
rect 56007 51940 57736 51981
rect 56007 51935 56267 51940
rect 55927 51894 56267 51935
rect 56313 51894 57736 51940
rect 55927 51817 57736 51894
rect 55927 51771 55961 51817
rect 56007 51777 57736 51817
rect 56007 51771 56267 51777
rect 55927 51731 56267 51771
rect 56313 51731 57736 51777
rect 55927 51654 57736 51731
rect 55927 51608 55961 51654
rect 56007 51613 57736 51654
rect 56007 51608 56267 51613
rect 55927 51567 56267 51608
rect 56313 51567 57736 51613
rect 34717 51401 34755 51453
rect 34807 51450 34935 51453
rect 34807 51404 34916 51450
rect 34807 51401 34935 51404
rect 34987 51401 35025 51453
rect 34717 51360 35025 51401
rect 50099 51453 50408 51494
rect 50099 51401 50138 51453
rect 50190 51450 50318 51453
rect 50206 51404 50318 51450
rect 50190 51401 50318 51404
rect 50370 51401 50408 51453
rect 27387 51241 28810 51287
rect 28856 51244 29196 51287
rect 28856 51241 29116 51244
rect 27387 51198 29116 51241
rect 29162 51198 29196 51244
rect 27387 51123 29196 51198
rect 27387 51077 28810 51123
rect 28856 51081 29196 51123
rect 28856 51077 29116 51081
rect 27387 51035 29116 51077
rect 29162 51035 29196 51081
rect 27387 50960 29196 51035
rect 27387 50914 28810 50960
rect 28856 50917 29196 50960
rect 28856 50914 29116 50917
rect 27387 50871 29116 50914
rect 29162 50871 29196 50917
rect 27387 50797 29196 50871
rect 27387 50751 28810 50797
rect 28856 50754 29196 50797
rect 28856 50751 29116 50754
rect 27387 50708 29116 50751
rect 29162 50708 29196 50754
rect 27387 50634 29196 50708
rect 27387 50588 28810 50634
rect 28856 50588 29196 50634
rect 30583 51327 31040 51360
rect 34870 51353 35025 51360
rect 30583 51287 30855 51327
rect 30583 51241 30637 51287
rect 30683 51281 30855 51287
rect 30901 51281 31040 51327
rect 35294 51315 36266 51355
rect 37853 51349 38161 51357
rect 35294 51309 35332 51315
rect 35384 51309 35543 51315
rect 35595 51309 35754 51315
rect 35806 51309 35965 51315
rect 36017 51309 36176 51315
rect 36228 51309 36266 51315
rect 36438 51309 36953 51349
rect 37439 51317 38161 51349
rect 37439 51309 37891 51317
rect 37943 51309 38071 51317
rect 38123 51309 38161 51317
rect 38658 51309 39723 51369
rect 50099 51360 50408 51401
rect 52278 51453 54540 51494
rect 52278 51401 52316 51453
rect 52368 51401 52527 51453
rect 52579 51401 52738 51453
rect 52790 51401 52948 51453
rect 53000 51401 53159 51453
rect 53211 51401 53371 51453
rect 53423 51401 53582 51453
rect 53634 51401 53792 51453
rect 53844 51401 54003 51453
rect 54055 51401 54214 51453
rect 54266 51450 54540 51453
rect 54266 51404 54440 51450
rect 54486 51404 54540 51450
rect 54266 51401 54540 51404
rect 52278 51360 54540 51401
rect 54758 51453 55840 51494
rect 54758 51450 54855 51453
rect 54758 51404 54793 51450
rect 54839 51404 54855 51450
rect 54758 51401 54855 51404
rect 54907 51450 55066 51453
rect 54907 51404 54956 51450
rect 55002 51404 55066 51450
rect 54907 51401 55066 51404
rect 55118 51450 55278 51453
rect 55330 51450 55489 51453
rect 55164 51404 55278 51450
rect 55330 51404 55439 51450
rect 55485 51404 55489 51450
rect 55118 51401 55278 51404
rect 55330 51401 55489 51404
rect 55541 51450 55840 51453
rect 55541 51404 55599 51450
rect 55645 51404 55760 51450
rect 55806 51404 55840 51450
rect 55541 51401 55840 51404
rect 54758 51361 55840 51401
rect 55927 51453 57736 51567
rect 55927 51401 56015 51453
rect 56067 51401 56226 51453
rect 56278 51450 56437 51453
rect 56313 51404 56437 51450
rect 56278 51401 56437 51404
rect 56489 51401 56648 51453
rect 56700 51401 56859 51453
rect 56911 51401 57070 51453
rect 57122 51401 57281 51453
rect 57333 51401 57736 51453
rect 54817 51360 55579 51361
rect 48905 51315 49877 51355
rect 50099 51353 50255 51360
rect 48905 51309 48943 51315
rect 48995 51309 49154 51315
rect 49206 51309 49365 51315
rect 49417 51309 49576 51315
rect 49628 51309 49787 51315
rect 49839 51309 49877 51315
rect 30683 51241 31040 51281
rect 33484 51265 34643 51294
rect 30583 51164 31040 51241
rect 33019 51225 33327 51265
rect 33019 51222 33057 51225
rect 33109 51222 33237 51225
rect 33289 51222 33327 51225
rect 33484 51257 35082 51265
rect 35260 51263 35273 51309
rect 35523 51263 35543 51309
rect 35626 51263 35683 51309
rect 35729 51263 35754 51309
rect 35832 51263 35889 51309
rect 35935 51263 35965 51309
rect 36038 51263 36095 51309
rect 36141 51263 36176 51309
rect 36244 51263 36301 51309
rect 36347 51263 36360 51309
rect 36438 51263 36854 51309
rect 36900 51263 36971 51309
rect 37017 51263 37088 51309
rect 37134 51263 37206 51309
rect 37252 51263 37324 51309
rect 37370 51263 37442 51309
rect 37488 51265 37891 51309
rect 37488 51263 37909 51265
rect 37955 51263 38026 51309
rect 38123 51265 38143 51309
rect 38072 51263 38143 51265
rect 38189 51263 38261 51309
rect 38307 51263 38379 51309
rect 38425 51263 38497 51309
rect 38543 51263 38556 51309
rect 38658 51263 39021 51309
rect 39067 51263 39144 51309
rect 39190 51263 39267 51309
rect 39313 51263 39641 51309
rect 39687 51263 39730 51309
rect 31336 51176 31349 51222
rect 33323 51176 33336 51222
rect 33484 51211 33816 51257
rect 33862 51211 34002 51257
rect 34048 51211 34189 51257
rect 34235 51211 34376 51257
rect 34422 51211 34562 51257
rect 34608 51211 35082 51257
rect 35294 51223 36266 51263
rect 36438 51229 36953 51263
rect 37439 51229 38161 51263
rect 30583 51123 30855 51164
rect 30583 51077 30637 51123
rect 30683 51118 30855 51123
rect 30901 51118 31040 51164
rect 33019 51173 33057 51176
rect 33109 51173 33237 51176
rect 33289 51173 33327 51176
rect 33019 51132 33327 51173
rect 33484 51174 35082 51211
rect 30683 51077 31040 51118
rect 30583 51049 31040 51077
rect 33484 51092 33552 51174
rect 30583 51001 31493 51049
rect 30583 50960 30855 51001
rect 30583 50914 30637 50960
rect 30683 50955 30855 50960
rect 30901 50998 31493 51001
rect 30901 50955 31349 50998
rect 30683 50952 31349 50955
rect 33323 50952 33336 50998
rect 30683 50930 31493 50952
rect 30683 50914 31040 50930
rect 30583 50838 31040 50914
rect 30583 50797 30855 50838
rect 30583 50751 30637 50797
rect 30683 50792 30855 50797
rect 30901 50792 31040 50838
rect 30683 50751 31040 50792
rect 33019 50777 33327 50817
rect 33019 50774 33057 50777
rect 33109 50774 33237 50777
rect 33289 50774 33327 50777
rect 30583 50674 31040 50751
rect 31336 50728 31349 50774
rect 33323 50728 33336 50774
rect 33019 50725 33057 50728
rect 33109 50725 33237 50728
rect 33289 50725 33327 50728
rect 33019 50684 33327 50725
rect 30583 50634 30855 50674
rect 27387 50466 29196 50588
rect 27387 50420 28810 50466
rect 28856 50420 29196 50466
rect 29283 50553 30365 50594
rect 29283 50550 29582 50553
rect 29283 50504 29317 50550
rect 29363 50504 29478 50550
rect 29524 50504 29582 50550
rect 29283 50501 29582 50504
rect 29634 50550 29793 50553
rect 29845 50550 30005 50553
rect 29634 50504 29638 50550
rect 29684 50504 29793 50550
rect 29845 50504 29959 50550
rect 29634 50501 29793 50504
rect 29845 50501 30005 50504
rect 30057 50550 30216 50553
rect 30057 50504 30121 50550
rect 30167 50504 30216 50550
rect 30057 50501 30216 50504
rect 30268 50550 30365 50553
rect 30268 50504 30284 50550
rect 30330 50504 30365 50550
rect 30268 50501 30365 50504
rect 29283 50461 30365 50501
rect 30583 50588 30637 50634
rect 30683 50628 30855 50634
rect 30901 50628 31040 50674
rect 33484 50670 33495 51092
rect 33541 50670 33552 51092
rect 34964 51117 35082 51174
rect 36438 51129 36554 51229
rect 37853 51224 38161 51229
rect 38658 51249 39723 51263
rect 34964 51085 36360 51117
rect 34228 51015 34718 51056
rect 34228 50998 34267 51015
rect 34319 50998 34447 51015
rect 34499 50998 34627 51015
rect 33671 50952 33684 50998
rect 33730 50952 33787 50998
rect 33833 50952 33890 50998
rect 33936 50952 33993 50998
rect 34039 50952 34096 50998
rect 34142 50952 34199 50998
rect 34245 50963 34267 50998
rect 34245 50952 34302 50963
rect 34348 50952 34405 50998
rect 34499 50963 34508 50998
rect 34451 50952 34508 50963
rect 34554 50952 34612 50998
rect 34679 50963 34718 51015
rect 34964 51039 35273 51085
rect 35523 51039 35580 51085
rect 35626 51039 35683 51085
rect 35729 51039 35786 51085
rect 35832 51039 35889 51085
rect 35935 51039 35992 51085
rect 36038 51039 36095 51085
rect 36141 51039 36198 51085
rect 36244 51039 36301 51085
rect 36347 51039 36360 51085
rect 34964 50995 36360 51039
rect 34658 50952 34718 50963
rect 34228 50923 34718 50952
rect 36438 50989 36475 51129
rect 36521 50989 36554 51129
rect 35294 50861 36266 50895
rect 36438 50886 36554 50989
rect 36640 51129 36773 51149
rect 36640 51090 36697 51129
rect 36640 51038 36678 51090
rect 36640 50989 36697 51038
rect 36743 50989 36773 51129
rect 38658 51127 38726 51249
rect 39809 51243 44918 51281
rect 48765 51263 48778 51309
rect 48824 51263 48881 51309
rect 48927 51263 48943 51309
rect 49030 51263 49087 51309
rect 49133 51263 49154 51309
rect 49236 51263 49293 51309
rect 49339 51263 49365 51309
rect 49442 51263 49499 51309
rect 49545 51263 49576 51309
rect 49852 51263 49877 51309
rect 54085 51327 54540 51360
rect 50481 51267 51657 51294
rect 39809 51197 43739 51243
rect 43785 51197 43906 51243
rect 43952 51197 44071 51243
rect 44117 51197 44236 51243
rect 44282 51222 44918 51243
rect 48905 51223 49877 51263
rect 50044 51257 51657 51267
rect 44282 51197 44812 51222
rect 39809 51194 44812 51197
rect 39809 51148 39844 51194
rect 39890 51192 44812 51194
rect 39890 51148 39994 51192
rect 39809 51140 39994 51148
rect 40046 51176 44812 51192
rect 44858 51176 44925 51222
rect 44971 51176 45038 51222
rect 45084 51176 45151 51222
rect 45197 51176 45264 51222
rect 45310 51176 45323 51222
rect 48557 51177 48687 51217
rect 40046 51161 44918 51176
rect 40046 51140 40085 51161
rect 39809 51137 40085 51140
rect 36924 51117 37685 51124
rect 36923 51085 37931 51117
rect 36841 51039 36854 51085
rect 36900 51083 36971 51085
rect 36900 51039 36961 51083
rect 37017 51039 37088 51085
rect 37134 51083 37206 51085
rect 37134 51039 37172 51083
rect 37252 51039 37324 51085
rect 37370 51083 37442 51085
rect 37370 51039 37384 51083
rect 36923 51031 36961 51039
rect 37013 51031 37172 51039
rect 37224 51031 37384 51039
rect 37436 51039 37442 51083
rect 37488 51083 37909 51085
rect 37488 51039 37595 51083
rect 37436 51031 37595 51039
rect 37647 51039 37909 51083
rect 37955 51039 38026 51085
rect 38072 51039 38143 51085
rect 38189 51039 38261 51085
rect 38307 51039 38379 51085
rect 38425 51039 38497 51085
rect 38543 51039 38556 51085
rect 37647 51031 37931 51039
rect 36923 50998 37931 51031
rect 36923 50997 37685 50998
rect 36924 50991 37685 50997
rect 36640 50966 36773 50989
rect 38658 50987 38669 51127
rect 38715 50987 38726 51127
rect 39014 51085 39323 51117
rect 39492 51085 39608 51117
rect 39008 51039 39021 51085
rect 39067 51039 39144 51085
rect 39190 51039 39267 51085
rect 39313 51039 39326 51085
rect 39492 51039 39641 51085
rect 39687 51039 39730 51085
rect 38658 50976 38726 50987
rect 36438 50861 36953 50886
rect 37439 50883 37931 50886
rect 37439 50861 38161 50883
rect 35260 50815 35273 50861
rect 35523 50855 35580 50861
rect 35523 50815 35543 50855
rect 35626 50815 35683 50861
rect 35729 50855 35786 50861
rect 35729 50815 35754 50855
rect 35832 50815 35889 50861
rect 35935 50855 35992 50861
rect 35935 50815 35965 50855
rect 36038 50815 36095 50861
rect 36141 50855 36198 50861
rect 36141 50815 36176 50855
rect 36244 50815 36301 50861
rect 36347 50815 36360 50861
rect 36438 50815 36854 50861
rect 36900 50815 36971 50861
rect 37017 50815 37088 50861
rect 37134 50815 37206 50861
rect 37252 50815 37324 50861
rect 37370 50815 37442 50861
rect 37488 50843 37909 50861
rect 37488 50815 37891 50843
rect 37955 50815 38026 50861
rect 38072 50843 38143 50861
rect 38123 50815 38143 50843
rect 38189 50815 38261 50861
rect 38307 50815 38379 50861
rect 38425 50815 38497 50861
rect 38543 50815 38556 50861
rect 33781 50774 34089 50809
rect 35294 50803 35332 50815
rect 35384 50803 35543 50815
rect 35595 50803 35754 50815
rect 35806 50803 35965 50815
rect 36017 50803 36176 50815
rect 36228 50803 36266 50815
rect 33671 50728 33684 50774
rect 33730 50728 33787 50774
rect 33833 50769 33890 50774
rect 33871 50728 33890 50769
rect 33936 50728 33993 50774
rect 34039 50769 34096 50774
rect 34051 50728 34096 50769
rect 34142 50728 34199 50774
rect 34245 50728 34302 50774
rect 34348 50728 34405 50774
rect 34451 50728 34508 50774
rect 34554 50728 34612 50774
rect 34658 50728 34671 50774
rect 35294 50763 36266 50803
rect 36438 50766 36953 50815
rect 37439 50791 37891 50815
rect 37943 50791 38071 50815
rect 38123 50791 38161 50815
rect 37439 50766 38161 50791
rect 37853 50750 38161 50766
rect 33781 50717 33819 50728
rect 33871 50717 33999 50728
rect 34051 50717 34089 50728
rect 33781 50676 34089 50717
rect 33484 50659 33552 50670
rect 30683 50594 31040 50628
rect 30683 50588 32842 50594
rect 30583 50553 32842 50588
rect 34247 50587 35008 50594
rect 30583 50501 30854 50553
rect 30906 50501 31065 50553
rect 31117 50501 31276 50553
rect 31328 50550 31486 50553
rect 31538 50550 31697 50553
rect 31749 50550 31909 50553
rect 31961 50550 32120 50553
rect 32172 50550 32330 50553
rect 32382 50550 32541 50553
rect 32593 50550 32752 50553
rect 32804 50550 32842 50553
rect 34246 50553 35008 50587
rect 34246 50550 34284 50553
rect 34336 50550 34495 50553
rect 34547 50550 34707 50553
rect 31328 50504 31349 50550
rect 33323 50504 33336 50550
rect 33671 50504 33684 50550
rect 33730 50504 33787 50550
rect 33833 50504 33890 50550
rect 33936 50504 33993 50550
rect 34039 50504 34096 50550
rect 34142 50504 34199 50550
rect 34245 50504 34284 50550
rect 34348 50504 34405 50550
rect 34451 50504 34495 50550
rect 34554 50504 34612 50550
rect 34658 50504 34707 50550
rect 31328 50501 31486 50504
rect 31538 50501 31697 50504
rect 31749 50501 31909 50504
rect 31961 50501 32120 50504
rect 32172 50501 32330 50504
rect 32382 50501 32541 50504
rect 32593 50501 32752 50504
rect 32804 50501 32842 50504
rect 30583 50466 32842 50501
rect 34246 50501 34284 50504
rect 34336 50501 34495 50504
rect 34547 50501 34707 50504
rect 34759 50501 34918 50553
rect 34970 50501 35008 50553
rect 34246 50467 35008 50501
rect 29544 50460 30306 50461
rect 27387 50344 29196 50420
rect 27387 50303 29116 50344
rect 27387 50257 28810 50303
rect 28856 50298 29116 50303
rect 29162 50298 29196 50344
rect 28856 50257 29196 50298
rect 27387 50181 29196 50257
rect 27387 50140 29116 50181
rect 27387 50094 28810 50140
rect 28856 50135 29116 50140
rect 29162 50135 29196 50181
rect 28856 50094 29196 50135
rect 27387 50017 29196 50094
rect 27387 49977 29116 50017
rect 27387 49931 28810 49977
rect 28856 49971 29116 49977
rect 29162 49971 29196 50017
rect 28856 49931 29196 49971
rect 27387 49854 29196 49931
rect 27387 49813 29116 49854
rect 27387 49767 28810 49813
rect 28856 49808 29116 49813
rect 29162 49808 29196 49854
rect 28856 49767 29196 49808
rect 27387 49653 29196 49767
rect 30583 50420 30637 50466
rect 30683 50460 32842 50466
rect 34247 50460 35008 50467
rect 35182 50587 36364 50594
rect 35182 50553 36958 50587
rect 35182 50501 35220 50553
rect 35272 50501 35430 50553
rect 35482 50501 35641 50553
rect 35693 50501 35853 50553
rect 35905 50501 36064 50553
rect 36116 50501 36274 50553
rect 36326 50550 36958 50553
rect 36326 50504 36489 50550
rect 36723 50504 36958 50550
rect 36326 50501 36958 50504
rect 35182 50467 36958 50501
rect 37946 50553 38842 50594
rect 37946 50550 38330 50553
rect 38382 50550 38541 50553
rect 37946 50504 37957 50550
rect 38473 50504 38541 50550
rect 37946 50501 38330 50504
rect 38382 50501 38541 50504
rect 38593 50501 38752 50553
rect 38804 50501 38842 50553
rect 35182 50460 36364 50467
rect 37946 50460 38842 50501
rect 39014 50553 39323 51039
rect 39014 50501 39052 50553
rect 39104 50550 39232 50553
rect 39108 50504 39220 50550
rect 39104 50501 39232 50504
rect 39284 50501 39323 50553
rect 30683 50426 31040 50460
rect 30683 50420 30855 50426
rect 30583 50380 30855 50420
rect 30901 50380 31040 50426
rect 30583 50303 31040 50380
rect 33484 50384 33552 50395
rect 33019 50329 33327 50370
rect 33019 50326 33057 50329
rect 33109 50326 33237 50329
rect 33289 50326 33327 50329
rect 30583 50257 30637 50303
rect 30683 50262 31040 50303
rect 31336 50280 31349 50326
rect 33323 50280 33336 50326
rect 30683 50257 30855 50262
rect 30583 50216 30855 50257
rect 30901 50216 31040 50262
rect 33019 50277 33057 50280
rect 33109 50277 33237 50280
rect 33289 50277 33327 50280
rect 33019 50237 33327 50277
rect 30583 50140 31040 50216
rect 30583 50094 30637 50140
rect 30683 50124 31040 50140
rect 30683 50102 31493 50124
rect 30683 50099 31349 50102
rect 30683 50094 30855 50099
rect 30583 50053 30855 50094
rect 30901 50056 31349 50099
rect 33323 50056 33336 50102
rect 30901 50053 31493 50056
rect 30583 50005 31493 50053
rect 30583 49977 31040 50005
rect 30583 49931 30637 49977
rect 30683 49936 31040 49977
rect 30683 49931 30855 49936
rect 30583 49890 30855 49931
rect 30901 49890 31040 49936
rect 33484 49962 33495 50384
rect 33541 49962 33552 50384
rect 33781 50337 34089 50378
rect 33781 50326 33819 50337
rect 33871 50326 33999 50337
rect 34051 50326 34089 50337
rect 33671 50280 33684 50326
rect 33730 50280 33787 50326
rect 33871 50285 33890 50326
rect 33833 50280 33890 50285
rect 33936 50280 33993 50326
rect 34051 50285 34096 50326
rect 34039 50280 34096 50285
rect 34142 50280 34199 50326
rect 34245 50280 34302 50326
rect 34348 50280 34405 50326
rect 34451 50280 34508 50326
rect 34554 50280 34612 50326
rect 34658 50280 34671 50326
rect 33781 50245 34089 50280
rect 35294 50251 36266 50291
rect 37853 50288 38161 50304
rect 35294 50239 35332 50251
rect 35384 50239 35543 50251
rect 35595 50239 35754 50251
rect 35806 50239 35965 50251
rect 36017 50239 36176 50251
rect 36228 50239 36266 50251
rect 36438 50239 36953 50288
rect 37439 50263 38161 50288
rect 37439 50239 37891 50263
rect 37943 50239 38071 50263
rect 38123 50239 38161 50263
rect 35260 50193 35273 50239
rect 35523 50199 35543 50239
rect 35523 50193 35580 50199
rect 35626 50193 35683 50239
rect 35729 50199 35754 50239
rect 35729 50193 35786 50199
rect 35832 50193 35889 50239
rect 35935 50199 35965 50239
rect 35935 50193 35992 50199
rect 36038 50193 36095 50239
rect 36141 50199 36176 50239
rect 36141 50193 36198 50199
rect 36244 50193 36301 50239
rect 36347 50193 36360 50239
rect 36438 50193 36854 50239
rect 36900 50193 36971 50239
rect 37017 50193 37088 50239
rect 37134 50193 37206 50239
rect 37252 50193 37324 50239
rect 37370 50193 37442 50239
rect 37488 50211 37891 50239
rect 37488 50193 37909 50211
rect 37955 50193 38026 50239
rect 38123 50211 38143 50239
rect 38072 50193 38143 50211
rect 38189 50193 38261 50239
rect 38307 50193 38379 50239
rect 38425 50193 38497 50239
rect 38543 50193 38556 50239
rect 35294 50159 36266 50193
rect 36438 50168 36953 50193
rect 37439 50171 38161 50193
rect 37439 50168 37931 50171
rect 34228 50102 34718 50131
rect 33671 50056 33684 50102
rect 33730 50056 33787 50102
rect 33833 50056 33890 50102
rect 33936 50056 33993 50102
rect 34039 50056 34096 50102
rect 34142 50056 34199 50102
rect 34245 50091 34302 50102
rect 34245 50056 34267 50091
rect 34348 50056 34405 50102
rect 34451 50091 34508 50102
rect 34499 50056 34508 50091
rect 34554 50056 34612 50102
rect 34658 50091 34718 50102
rect 34228 50039 34267 50056
rect 34319 50039 34447 50056
rect 34499 50039 34627 50056
rect 34679 50039 34718 50091
rect 36438 50065 36554 50168
rect 34228 49998 34718 50039
rect 34964 50015 36360 50059
rect 30583 49813 31040 49890
rect 33019 49881 33327 49922
rect 33019 49878 33057 49881
rect 33109 49878 33237 49881
rect 33289 49878 33327 49881
rect 33484 49880 33552 49962
rect 34964 49969 35273 50015
rect 35523 49969 35580 50015
rect 35626 49969 35683 50015
rect 35729 49969 35786 50015
rect 35832 49969 35889 50015
rect 35935 49969 35992 50015
rect 36038 49969 36095 50015
rect 36141 49969 36198 50015
rect 36244 49969 36301 50015
rect 36347 49969 36360 50015
rect 34964 49937 36360 49969
rect 34964 49880 35082 49937
rect 31336 49832 31349 49878
rect 33323 49832 33336 49878
rect 33484 49843 35082 49880
rect 30583 49767 30637 49813
rect 30683 49773 31040 49813
rect 33019 49829 33057 49832
rect 33109 49829 33237 49832
rect 33289 49829 33327 49832
rect 33019 49789 33327 49829
rect 33484 49797 33816 49843
rect 33862 49797 34002 49843
rect 34048 49797 34189 49843
rect 34235 49797 34376 49843
rect 34422 49797 34562 49843
rect 34608 49797 35082 49843
rect 36438 49925 36475 50065
rect 36521 49925 36554 50065
rect 33484 49789 35082 49797
rect 35294 49791 36266 49831
rect 36438 49825 36554 49925
rect 36640 50065 36773 50088
rect 36640 50016 36697 50065
rect 36640 49964 36678 50016
rect 36640 49925 36697 49964
rect 36743 49925 36773 50065
rect 38658 50067 38726 50078
rect 36924 50057 37685 50063
rect 36923 50056 37685 50057
rect 36923 50023 37931 50056
rect 36923 50015 36961 50023
rect 37013 50015 37172 50023
rect 37224 50015 37384 50023
rect 36841 49969 36854 50015
rect 36900 49971 36961 50015
rect 36900 49969 36971 49971
rect 37017 49969 37088 50015
rect 37134 49971 37172 50015
rect 37134 49969 37206 49971
rect 37252 49969 37324 50015
rect 37370 49971 37384 50015
rect 37436 50015 37595 50023
rect 37436 49971 37442 50015
rect 37370 49969 37442 49971
rect 37488 49971 37595 50015
rect 37647 50015 37931 50023
rect 37647 49971 37909 50015
rect 37488 49969 37909 49971
rect 37955 49969 38026 50015
rect 38072 49969 38143 50015
rect 38189 49969 38261 50015
rect 38307 49969 38379 50015
rect 38425 49969 38497 50015
rect 38543 49969 38556 50015
rect 36923 49937 37931 49969
rect 36924 49930 37685 49937
rect 36640 49905 36773 49925
rect 38658 49927 38669 50067
rect 38715 49927 38726 50067
rect 39014 50015 39323 50501
rect 39492 50587 39608 51039
rect 39923 51006 40085 51137
rect 39923 50954 39994 51006
rect 40046 50954 40085 51006
rect 39923 50914 40085 50954
rect 39737 50818 39865 50831
rect 39737 50791 39866 50818
rect 39737 50774 39775 50791
rect 39827 50774 39866 50791
rect 39727 50728 39740 50774
rect 39827 50739 39862 50774
rect 39786 50728 39862 50739
rect 39908 50728 39985 50774
rect 40031 50728 40108 50774
rect 40154 50728 40167 50774
rect 40246 50763 40362 51161
rect 42229 51022 44509 51063
rect 42229 50970 42690 51022
rect 42742 50970 44509 51022
rect 42229 50930 44509 50970
rect 44341 50886 44509 50930
rect 44341 50840 44358 50886
rect 44498 50840 44509 50886
rect 39737 50699 39866 50728
rect 40246 50717 40281 50763
rect 40327 50717 40362 50763
rect 40246 50680 40362 50717
rect 40718 50791 43524 50832
rect 44341 50829 44509 50840
rect 40718 50739 41935 50791
rect 41987 50739 43524 50791
rect 40718 50698 43524 50739
rect 44605 50774 44721 51161
rect 45400 51131 48379 51172
rect 45400 51117 48241 51131
rect 45400 51071 45464 51117
rect 45604 51079 48241 51117
rect 48293 51079 48379 51131
rect 45604 51071 48379 51079
rect 44901 51015 45241 51056
rect 45400 51038 48379 51071
rect 48557 51125 48596 51177
rect 48648 51125 48687 51177
rect 48557 51102 48687 51125
rect 50044 51211 50516 51257
rect 50562 51211 50703 51257
rect 50749 51211 50890 51257
rect 50936 51211 51076 51257
rect 51122 51211 51263 51257
rect 51309 51211 51657 51257
rect 51797 51247 52105 51287
rect 51797 51222 51835 51247
rect 51887 51222 52015 51247
rect 52067 51222 52105 51247
rect 54085 51281 54223 51327
rect 54269 51287 54540 51327
rect 54269 51281 54440 51287
rect 54085 51241 54440 51281
rect 54486 51241 54540 51287
rect 50044 51174 51657 51211
rect 51789 51176 51802 51222
rect 53776 51176 53789 51222
rect 50044 51117 50160 51174
rect 44901 50998 44939 51015
rect 44991 50998 45151 51015
rect 45203 50998 45241 51015
rect 44799 50952 44812 50998
rect 44858 50952 44925 50998
rect 44991 50963 45038 50998
rect 44971 50952 45038 50963
rect 45084 50952 45151 50998
rect 45203 50963 45264 50998
rect 45197 50952 45264 50963
rect 45310 50952 45323 50998
rect 48557 50962 48622 51102
rect 48668 50962 48687 51102
rect 49820 51085 50160 51117
rect 48765 51039 48778 51085
rect 48824 51039 48881 51085
rect 48927 51039 48984 51085
rect 49030 51039 49087 51085
rect 49133 51039 49190 51085
rect 49236 51039 49293 51085
rect 49339 51039 49396 51085
rect 49442 51039 49499 51085
rect 49545 51039 49602 51085
rect 49852 51039 50160 51085
rect 51589 51122 51657 51174
rect 51797 51154 52105 51176
rect 49820 50998 50160 51039
rect 50262 51015 50812 51056
rect 48557 50959 48687 50962
rect 44901 50923 45241 50952
rect 48557 50907 48596 50959
rect 48648 50907 48687 50959
rect 50262 50963 50300 51015
rect 50352 50998 50511 51015
rect 50563 50998 50722 51015
rect 50352 50963 50467 50998
rect 50563 50963 50571 50998
rect 50262 50952 50467 50963
rect 50513 50952 50571 50963
rect 50617 50952 50674 50998
rect 50720 50963 50722 50998
rect 50774 50998 50812 51015
rect 50774 50963 50777 50998
rect 50720 50952 50777 50963
rect 50823 50952 50880 50998
rect 50926 50952 50983 50998
rect 51029 50952 51086 50998
rect 51132 50952 51189 50998
rect 51235 50952 51292 50998
rect 51338 50952 51395 50998
rect 51441 50952 51454 50998
rect 50262 50923 50812 50952
rect 48557 50866 48687 50907
rect 48905 50861 49877 50892
rect 48765 50815 48778 50861
rect 48824 50815 48881 50861
rect 48927 50852 48984 50861
rect 48927 50815 48943 50852
rect 49030 50815 49087 50861
rect 49133 50852 49190 50861
rect 49133 50815 49154 50852
rect 49236 50815 49293 50861
rect 49339 50852 49396 50861
rect 49339 50815 49365 50852
rect 49442 50815 49499 50861
rect 49545 50852 49602 50861
rect 49545 50815 49576 50852
rect 49852 50815 49877 50861
rect 48905 50800 48943 50815
rect 48995 50800 49154 50815
rect 49206 50800 49365 50815
rect 49417 50800 49576 50815
rect 49628 50800 49787 50815
rect 49839 50800 49877 50815
rect 44605 50728 44812 50774
rect 44858 50728 44925 50774
rect 44971 50728 45038 50774
rect 45084 50728 45151 50774
rect 45197 50728 45264 50774
rect 45310 50728 45323 50774
rect 48905 50760 49877 50800
rect 51035 50777 51343 50817
rect 51035 50774 51073 50777
rect 51125 50774 51253 50777
rect 51305 50774 51343 50777
rect 43362 50691 43524 50698
rect 43362 50645 43373 50691
rect 43513 50645 43524 50691
rect 43362 50634 43524 50645
rect 45584 50714 48546 50750
rect 50454 50728 50467 50774
rect 50513 50728 50571 50774
rect 50617 50728 50674 50774
rect 50720 50728 50777 50774
rect 50823 50728 50880 50774
rect 50926 50728 50983 50774
rect 51029 50728 51073 50774
rect 51132 50728 51189 50774
rect 51235 50728 51253 50774
rect 51338 50728 51395 50774
rect 51441 50728 51454 50774
rect 45584 50668 45619 50714
rect 45665 50668 45777 50714
rect 45823 50668 45935 50714
rect 45981 50668 46093 50714
rect 46139 50668 46251 50714
rect 46297 50668 46409 50714
rect 46455 50668 46568 50714
rect 46614 50668 46726 50714
rect 46772 50668 46884 50714
rect 46930 50668 47042 50714
rect 47088 50668 47200 50714
rect 47246 50668 47358 50714
rect 47404 50668 47516 50714
rect 47562 50668 47675 50714
rect 47721 50668 47833 50714
rect 47879 50668 47991 50714
rect 48037 50668 48149 50714
rect 48195 50668 48307 50714
rect 48353 50668 48465 50714
rect 48511 50668 48546 50714
rect 51035 50725 51073 50728
rect 51125 50725 51253 50728
rect 51305 50725 51343 50728
rect 51035 50684 51343 50725
rect 51589 50700 51600 51122
rect 51646 50700 51657 51122
rect 54085 51123 54540 51241
rect 54085 51077 54440 51123
rect 54486 51077 54540 51123
rect 54085 51049 54540 51077
rect 53585 50998 54540 51049
rect 51789 50952 51802 50998
rect 53776 50960 54540 50998
rect 53776 50952 54440 50960
rect 53585 50930 54440 50952
rect 54085 50914 54440 50930
rect 54486 50914 54540 50960
rect 54085 50838 54540 50914
rect 51797 50784 52105 50824
rect 51797 50774 51835 50784
rect 51887 50774 52015 50784
rect 52067 50774 52105 50784
rect 54085 50792 54223 50838
rect 54269 50797 54540 50838
rect 54269 50792 54440 50797
rect 51789 50728 51802 50774
rect 53776 50728 53789 50774
rect 54085 50751 54440 50792
rect 54486 50751 54540 50797
rect 51589 50689 51657 50700
rect 51797 50691 52105 50728
rect 40215 50587 40523 50594
rect 40788 50587 42986 50601
rect 43753 50587 44514 50594
rect 39492 50564 42986 50587
rect 43704 50564 44514 50587
rect 39492 50553 44514 50564
rect 39492 50550 40253 50553
rect 39492 50504 39740 50550
rect 39786 50504 39862 50550
rect 39908 50504 39985 50550
rect 40031 50504 40108 50550
rect 40154 50504 40253 50550
rect 39492 50501 40253 50504
rect 40305 50501 40433 50553
rect 40485 50550 43790 50553
rect 40485 50504 40836 50550
rect 40882 50504 40994 50550
rect 41040 50504 41152 50550
rect 41198 50504 41310 50550
rect 41356 50504 41469 50550
rect 41515 50504 41627 50550
rect 41673 50504 41785 50550
rect 41831 50504 41943 50550
rect 41989 50504 42101 50550
rect 42147 50504 42259 50550
rect 42305 50504 42418 50550
rect 42464 50504 42576 50550
rect 42622 50504 42734 50550
rect 42780 50504 42892 50550
rect 42938 50504 43739 50550
rect 43785 50504 43790 50550
rect 40485 50501 43790 50504
rect 43842 50550 44001 50553
rect 43842 50504 43906 50550
rect 43952 50504 44001 50550
rect 43842 50501 44001 50504
rect 44053 50550 44213 50553
rect 44265 50550 44424 50553
rect 44053 50504 44071 50550
rect 44117 50504 44213 50550
rect 44282 50504 44424 50550
rect 44053 50501 44213 50504
rect 44265 50501 44424 50504
rect 44476 50501 44514 50553
rect 39492 50490 44514 50501
rect 39492 50467 42986 50490
rect 43704 50467 44514 50490
rect 39492 50015 39608 50467
rect 40215 50460 40523 50467
rect 40788 50453 42986 50467
rect 43753 50460 44514 50467
rect 44796 50587 45346 50594
rect 45584 50587 48546 50668
rect 54085 50674 54540 50751
rect 54085 50628 54223 50674
rect 54269 50634 54540 50674
rect 54269 50628 54440 50634
rect 54085 50594 54440 50628
rect 48800 50587 49982 50594
rect 50308 50587 50859 50594
rect 44796 50553 49982 50587
rect 44796 50550 44834 50553
rect 44886 50550 45045 50553
rect 45097 50550 45256 50553
rect 45308 50550 48838 50553
rect 44796 50504 44812 50550
rect 44886 50504 44925 50550
rect 44971 50504 45038 50550
rect 45097 50504 45151 50550
rect 45197 50504 45256 50550
rect 45310 50504 45619 50550
rect 45665 50504 45777 50550
rect 45823 50504 45935 50550
rect 45981 50504 46093 50550
rect 46139 50504 46251 50550
rect 46297 50504 46409 50550
rect 46455 50504 46568 50550
rect 46614 50504 46726 50550
rect 46772 50504 46884 50550
rect 46930 50504 47042 50550
rect 47088 50504 47200 50550
rect 47246 50504 47358 50550
rect 47404 50504 47516 50550
rect 47562 50504 47675 50550
rect 47721 50504 47833 50550
rect 47879 50504 47991 50550
rect 48037 50504 48149 50550
rect 48195 50504 48307 50550
rect 48353 50504 48465 50550
rect 48511 50504 48838 50550
rect 44796 50501 44834 50504
rect 44886 50501 45045 50504
rect 45097 50501 45256 50504
rect 45308 50501 48838 50504
rect 48890 50501 49048 50553
rect 49100 50501 49259 50553
rect 49311 50501 49471 50553
rect 49523 50501 49682 50553
rect 49734 50501 49892 50553
rect 49944 50501 49982 50553
rect 44796 50467 49982 50501
rect 50307 50553 50859 50587
rect 50307 50501 50346 50553
rect 50398 50550 50557 50553
rect 50609 50550 50768 50553
rect 50820 50550 50859 50553
rect 52278 50588 54440 50594
rect 54486 50588 54540 50634
rect 55927 51287 57736 51401
rect 55927 51244 56267 51287
rect 55927 51198 55961 51244
rect 56007 51241 56267 51244
rect 56313 51241 57736 51287
rect 56007 51198 57736 51241
rect 55927 51123 57736 51198
rect 55927 51081 56267 51123
rect 55927 51035 55961 51081
rect 56007 51077 56267 51081
rect 56313 51077 57736 51123
rect 56007 51035 57736 51077
rect 55927 50960 57736 51035
rect 55927 50917 56267 50960
rect 55927 50871 55961 50917
rect 56007 50914 56267 50917
rect 56313 50914 57736 50960
rect 56007 50871 57736 50914
rect 55927 50797 57736 50871
rect 55927 50754 56267 50797
rect 55927 50708 55961 50754
rect 56007 50751 56267 50754
rect 56313 50751 57736 50797
rect 56007 50708 57736 50751
rect 55927 50634 57736 50708
rect 52278 50553 54540 50588
rect 52278 50550 52316 50553
rect 52368 50550 52527 50553
rect 52579 50550 52738 50553
rect 52790 50550 52948 50553
rect 53000 50550 53159 50553
rect 53211 50550 53371 50553
rect 53423 50550 53582 50553
rect 53634 50550 53792 50553
rect 50398 50504 50467 50550
rect 50513 50504 50557 50550
rect 50617 50504 50674 50550
rect 50720 50504 50768 50550
rect 50823 50504 50880 50550
rect 50926 50504 50983 50550
rect 51029 50504 51086 50550
rect 51132 50504 51189 50550
rect 51235 50504 51292 50550
rect 51338 50504 51395 50550
rect 51441 50504 51454 50550
rect 51789 50504 51802 50550
rect 53776 50504 53792 50550
rect 50398 50501 50557 50504
rect 50609 50501 50768 50504
rect 50820 50501 50859 50504
rect 50307 50467 50859 50501
rect 44796 50460 45346 50467
rect 43362 50409 43524 50420
rect 39737 50326 39866 50355
rect 40246 50337 40362 50374
rect 43362 50363 43373 50409
rect 43513 50363 43524 50409
rect 43362 50356 43524 50363
rect 39727 50280 39740 50326
rect 39786 50315 39862 50326
rect 39827 50280 39862 50315
rect 39908 50280 39985 50326
rect 40031 50280 40108 50326
rect 40154 50280 40167 50326
rect 40246 50291 40281 50337
rect 40327 50291 40362 50337
rect 39737 50263 39775 50280
rect 39827 50263 39866 50280
rect 39737 50236 39866 50263
rect 39737 50223 39865 50236
rect 39923 50100 40085 50140
rect 39923 50048 39994 50100
rect 40046 50048 40085 50100
rect 39008 49969 39021 50015
rect 39067 49969 39144 50015
rect 39190 49969 39267 50015
rect 39313 49969 39326 50015
rect 39492 49969 39641 50015
rect 39687 49969 39730 50015
rect 39014 49937 39323 49969
rect 39492 49937 39608 49969
rect 37853 49825 38161 49830
rect 36438 49791 36953 49825
rect 37439 49791 38161 49825
rect 38658 49805 38726 49927
rect 39923 49917 40085 50048
rect 39809 49914 40085 49917
rect 39809 49906 39994 49914
rect 39809 49860 39844 49906
rect 39890 49862 39994 49906
rect 40046 49893 40085 49914
rect 40246 49893 40362 50291
rect 40718 50315 43524 50356
rect 45584 50386 48546 50467
rect 48800 50460 49982 50467
rect 50308 50460 50859 50467
rect 52278 50501 52316 50504
rect 52368 50501 52527 50504
rect 52579 50501 52738 50504
rect 52790 50501 52948 50504
rect 53000 50501 53159 50504
rect 53211 50501 53371 50504
rect 53423 50501 53582 50504
rect 53634 50501 53792 50504
rect 53844 50501 54003 50553
rect 54055 50501 54214 50553
rect 54266 50501 54540 50553
rect 52278 50466 54540 50501
rect 52278 50460 54440 50466
rect 45584 50340 45619 50386
rect 45665 50340 45777 50386
rect 45823 50340 45935 50386
rect 45981 50340 46093 50386
rect 46139 50340 46251 50386
rect 46297 50340 46409 50386
rect 46455 50340 46568 50386
rect 46614 50340 46726 50386
rect 46772 50340 46884 50386
rect 46930 50340 47042 50386
rect 47088 50340 47200 50386
rect 47246 50340 47358 50386
rect 47404 50340 47516 50386
rect 47562 50340 47675 50386
rect 47721 50340 47833 50386
rect 47879 50340 47991 50386
rect 48037 50340 48149 50386
rect 48195 50340 48307 50386
rect 48353 50340 48465 50386
rect 48511 50340 48546 50386
rect 54085 50426 54440 50460
rect 54085 50380 54223 50426
rect 54269 50420 54440 50426
rect 54486 50420 54540 50466
rect 54758 50553 55840 50594
rect 54758 50550 54855 50553
rect 54758 50504 54793 50550
rect 54839 50504 54855 50550
rect 54758 50501 54855 50504
rect 54907 50550 55066 50553
rect 54907 50504 54956 50550
rect 55002 50504 55066 50550
rect 54907 50501 55066 50504
rect 55118 50550 55278 50553
rect 55330 50550 55489 50553
rect 55164 50504 55278 50550
rect 55330 50504 55439 50550
rect 55485 50504 55489 50550
rect 55118 50501 55278 50504
rect 55330 50501 55489 50504
rect 55541 50550 55840 50553
rect 55541 50504 55599 50550
rect 55645 50504 55760 50550
rect 55806 50504 55840 50550
rect 55541 50501 55840 50504
rect 54758 50461 55840 50501
rect 55927 50588 56267 50634
rect 56313 50588 57736 50634
rect 55927 50466 57736 50588
rect 54817 50460 55579 50461
rect 54269 50380 54540 50420
rect 40718 50263 41935 50315
rect 41987 50263 43524 50315
rect 40718 50222 43524 50263
rect 44605 50280 44812 50326
rect 44858 50280 44925 50326
rect 44971 50280 45038 50326
rect 45084 50280 45151 50326
rect 45197 50280 45264 50326
rect 45310 50280 45323 50326
rect 45584 50304 48546 50340
rect 51035 50329 51343 50370
rect 51035 50326 51073 50329
rect 51125 50326 51253 50329
rect 51305 50326 51343 50329
rect 51589 50354 51657 50365
rect 44341 50214 44509 50225
rect 44341 50168 44358 50214
rect 44498 50168 44509 50214
rect 44341 50124 44509 50168
rect 42229 50084 44509 50124
rect 42229 50032 43068 50084
rect 43120 50032 44509 50084
rect 42229 49991 44509 50032
rect 44605 49893 44721 50280
rect 48905 50254 49877 50294
rect 50454 50280 50467 50326
rect 50513 50280 50571 50326
rect 50617 50280 50674 50326
rect 50720 50280 50777 50326
rect 50823 50280 50880 50326
rect 50926 50280 50983 50326
rect 51029 50280 51073 50326
rect 51132 50280 51189 50326
rect 51235 50280 51253 50326
rect 51338 50280 51395 50326
rect 51441 50280 51454 50326
rect 48905 50239 48943 50254
rect 48995 50239 49154 50254
rect 49206 50239 49365 50254
rect 49417 50239 49576 50254
rect 49628 50239 49787 50254
rect 49839 50239 49877 50254
rect 48765 50193 48778 50239
rect 48824 50193 48881 50239
rect 48927 50202 48943 50239
rect 48927 50193 48984 50202
rect 49030 50193 49087 50239
rect 49133 50202 49154 50239
rect 49133 50193 49190 50202
rect 49236 50193 49293 50239
rect 49339 50202 49365 50239
rect 49339 50193 49396 50202
rect 49442 50193 49499 50239
rect 49545 50202 49576 50239
rect 49545 50193 49602 50202
rect 49852 50193 49877 50239
rect 51035 50277 51073 50280
rect 51125 50277 51253 50280
rect 51305 50277 51343 50280
rect 51035 50237 51343 50277
rect 48557 50147 48687 50188
rect 48905 50162 49877 50193
rect 44901 50102 45241 50131
rect 44799 50056 44812 50102
rect 44858 50056 44925 50102
rect 44971 50091 45038 50102
rect 44991 50056 45038 50091
rect 45084 50056 45151 50102
rect 45197 50091 45264 50102
rect 45203 50056 45264 50091
rect 45310 50056 45323 50102
rect 48557 50095 48596 50147
rect 48648 50095 48687 50147
rect 48557 50092 48687 50095
rect 44901 50039 44939 50056
rect 44991 50039 45151 50056
rect 45203 50039 45241 50056
rect 44901 49998 45241 50039
rect 45400 49983 48379 50016
rect 45400 49937 45464 49983
rect 45604 49975 48379 49983
rect 45400 49923 45597 49937
rect 45649 49923 48379 49975
rect 40046 49878 44918 49893
rect 45400 49882 48379 49923
rect 48557 49952 48622 50092
rect 48668 49952 48687 50092
rect 50262 50102 50812 50131
rect 50262 50091 50467 50102
rect 50513 50091 50571 50102
rect 49820 50015 50160 50056
rect 48765 49969 48778 50015
rect 48824 49969 48881 50015
rect 48927 49969 48984 50015
rect 49030 49969 49087 50015
rect 49133 49969 49190 50015
rect 49236 49969 49293 50015
rect 49339 49969 49396 50015
rect 49442 49969 49499 50015
rect 49545 49969 49602 50015
rect 49852 49969 50160 50015
rect 50262 50039 50300 50091
rect 50352 50056 50467 50091
rect 50563 50056 50571 50091
rect 50617 50056 50674 50102
rect 50720 50091 50777 50102
rect 50720 50056 50722 50091
rect 50352 50039 50511 50056
rect 50563 50039 50722 50056
rect 50774 50056 50777 50091
rect 50823 50056 50880 50102
rect 50926 50056 50983 50102
rect 51029 50056 51086 50102
rect 51132 50056 51189 50102
rect 51235 50056 51292 50102
rect 51338 50056 51395 50102
rect 51441 50056 51454 50102
rect 50774 50039 50812 50056
rect 50262 49998 50812 50039
rect 48557 49929 48687 49952
rect 49820 49937 50160 49969
rect 40046 49862 44812 49878
rect 39890 49860 44812 49862
rect 39809 49857 44812 49860
rect 39809 49811 43739 49857
rect 43785 49811 43906 49857
rect 43952 49811 44071 49857
rect 44117 49811 44236 49857
rect 44282 49832 44812 49857
rect 44858 49832 44925 49878
rect 44971 49832 45038 49878
rect 45084 49832 45151 49878
rect 45197 49832 45264 49878
rect 45310 49832 45323 49878
rect 48557 49877 48596 49929
rect 48648 49877 48687 49929
rect 48557 49837 48687 49877
rect 50044 49880 50160 49937
rect 51589 49932 51600 50354
rect 51646 49932 51657 50354
rect 51797 50326 52105 50363
rect 51789 50280 51802 50326
rect 53776 50280 53789 50326
rect 54085 50303 54540 50380
rect 51797 50270 51835 50280
rect 51887 50270 52015 50280
rect 52067 50270 52105 50280
rect 51797 50230 52105 50270
rect 54085 50262 54440 50303
rect 54085 50216 54223 50262
rect 54269 50257 54440 50262
rect 54486 50257 54540 50303
rect 54269 50216 54540 50257
rect 54085 50140 54540 50216
rect 54085 50124 54440 50140
rect 53585 50102 54440 50124
rect 51789 50056 51802 50102
rect 53776 50094 54440 50102
rect 54486 50094 54540 50140
rect 53776 50056 54540 50094
rect 53585 50005 54540 50056
rect 51589 49880 51657 49932
rect 54085 49977 54540 50005
rect 54085 49931 54440 49977
rect 54486 49931 54540 49977
rect 50044 49843 51657 49880
rect 51797 49878 52105 49900
rect 44282 49811 44918 49832
rect 38658 49791 39723 49805
rect 30683 49767 30855 49773
rect 30583 49727 30855 49767
rect 30901 49727 31040 49773
rect 33484 49760 34643 49789
rect 35260 49745 35273 49791
rect 35523 49745 35543 49791
rect 35626 49745 35683 49791
rect 35729 49745 35754 49791
rect 35832 49745 35889 49791
rect 35935 49745 35965 49791
rect 36038 49745 36095 49791
rect 36141 49745 36176 49791
rect 36244 49745 36301 49791
rect 36347 49745 36360 49791
rect 36438 49745 36854 49791
rect 36900 49745 36971 49791
rect 37017 49745 37088 49791
rect 37134 49745 37206 49791
rect 37252 49745 37324 49791
rect 37370 49745 37442 49791
rect 37488 49789 37909 49791
rect 37488 49745 37891 49789
rect 37955 49745 38026 49791
rect 38072 49789 38143 49791
rect 38123 49745 38143 49789
rect 38189 49745 38261 49791
rect 38307 49745 38379 49791
rect 38425 49745 38497 49791
rect 38543 49745 38556 49791
rect 38658 49745 39021 49791
rect 39067 49745 39144 49791
rect 39190 49745 39267 49791
rect 39313 49745 39641 49791
rect 39687 49745 39730 49791
rect 39809 49773 44918 49811
rect 48905 49791 49877 49831
rect 48765 49745 48778 49791
rect 48824 49745 48881 49791
rect 48927 49745 48943 49791
rect 49030 49745 49087 49791
rect 49133 49745 49154 49791
rect 49236 49745 49293 49791
rect 49339 49745 49365 49791
rect 49442 49745 49499 49791
rect 49545 49745 49576 49791
rect 49852 49745 49877 49791
rect 50044 49797 50516 49843
rect 50562 49797 50703 49843
rect 50749 49797 50890 49843
rect 50936 49797 51076 49843
rect 51122 49797 51263 49843
rect 51309 49797 51657 49843
rect 51789 49832 51802 49878
rect 53776 49832 53789 49878
rect 50044 49787 51657 49797
rect 50481 49760 51657 49787
rect 51797 49807 51835 49832
rect 51887 49807 52015 49832
rect 52067 49807 52105 49832
rect 51797 49767 52105 49807
rect 54085 49813 54540 49931
rect 54085 49773 54440 49813
rect 30583 49694 31040 49727
rect 35294 49739 35332 49745
rect 35384 49739 35543 49745
rect 35595 49739 35754 49745
rect 35806 49739 35965 49745
rect 36017 49739 36176 49745
rect 36228 49739 36266 49745
rect 34870 49694 35025 49701
rect 35294 49699 36266 49739
rect 36438 49705 36953 49745
rect 37439 49737 37891 49745
rect 37943 49737 38071 49745
rect 38123 49737 38161 49745
rect 37439 49705 38161 49737
rect 37853 49697 38161 49705
rect 27387 49601 27790 49653
rect 27842 49601 28001 49653
rect 28053 49601 28212 49653
rect 28264 49601 28423 49653
rect 28475 49601 28634 49653
rect 28686 49650 28845 49653
rect 28686 49604 28810 49650
rect 28686 49601 28845 49604
rect 28897 49601 29056 49653
rect 29108 49601 29196 49653
rect 27387 49487 29196 49601
rect 29283 49653 30365 49694
rect 29283 49650 29582 49653
rect 29283 49604 29317 49650
rect 29363 49604 29478 49650
rect 29524 49604 29582 49650
rect 29283 49601 29582 49604
rect 29634 49650 29793 49653
rect 29845 49650 30005 49653
rect 29634 49604 29638 49650
rect 29684 49604 29793 49650
rect 29845 49604 29959 49650
rect 29634 49601 29793 49604
rect 29845 49601 30005 49604
rect 30057 49650 30216 49653
rect 30057 49604 30121 49650
rect 30167 49604 30216 49650
rect 30057 49601 30216 49604
rect 30268 49650 30365 49653
rect 30268 49604 30284 49650
rect 30330 49604 30365 49650
rect 30268 49601 30365 49604
rect 29283 49561 30365 49601
rect 30583 49653 32842 49694
rect 30583 49650 30854 49653
rect 30583 49604 30637 49650
rect 30683 49604 30854 49650
rect 30583 49601 30854 49604
rect 30906 49601 31065 49653
rect 31117 49601 31276 49653
rect 31328 49601 31486 49653
rect 31538 49601 31697 49653
rect 31749 49601 31909 49653
rect 31961 49601 32120 49653
rect 32172 49601 32330 49653
rect 32382 49601 32541 49653
rect 32593 49601 32752 49653
rect 32804 49601 32842 49653
rect 29544 49560 30306 49561
rect 30583 49560 32842 49601
rect 34717 49653 35025 49694
rect 38658 49685 39723 49745
rect 48905 49739 48943 49745
rect 48995 49739 49154 49745
rect 49206 49739 49365 49745
rect 49417 49739 49576 49745
rect 49628 49739 49787 49745
rect 49839 49739 49877 49745
rect 48905 49699 49877 49739
rect 54085 49727 54223 49773
rect 54269 49767 54440 49773
rect 54486 49767 54540 49813
rect 54269 49727 54540 49767
rect 50099 49694 50255 49701
rect 54085 49694 54540 49727
rect 55927 50420 56267 50466
rect 56313 50420 57736 50466
rect 55927 50344 57736 50420
rect 55927 50298 55961 50344
rect 56007 50303 57736 50344
rect 56007 50298 56267 50303
rect 55927 50257 56267 50298
rect 56313 50257 57736 50303
rect 55927 50181 57736 50257
rect 55927 50135 55961 50181
rect 56007 50140 57736 50181
rect 56007 50135 56267 50140
rect 55927 50094 56267 50135
rect 56313 50094 57736 50140
rect 55927 50017 57736 50094
rect 55927 49971 55961 50017
rect 56007 49977 57736 50017
rect 56007 49971 56267 49977
rect 55927 49931 56267 49971
rect 56313 49931 57736 49977
rect 55927 49854 57736 49931
rect 55927 49808 55961 49854
rect 56007 49813 57736 49854
rect 56007 49808 56267 49813
rect 55927 49767 56267 49808
rect 56313 49767 57736 49813
rect 34717 49601 34755 49653
rect 34807 49650 34935 49653
rect 34807 49604 34916 49650
rect 34807 49601 34935 49604
rect 34987 49601 35025 49653
rect 34717 49560 35025 49601
rect 50099 49653 50408 49694
rect 50099 49601 50138 49653
rect 50190 49650 50318 49653
rect 50206 49604 50318 49650
rect 50190 49601 50318 49604
rect 50370 49601 50408 49653
rect 27387 49441 28810 49487
rect 28856 49444 29196 49487
rect 28856 49441 29116 49444
rect 27387 49398 29116 49441
rect 29162 49398 29196 49444
rect 27387 49323 29196 49398
rect 27387 49277 28810 49323
rect 28856 49281 29196 49323
rect 28856 49277 29116 49281
rect 27387 49235 29116 49277
rect 29162 49235 29196 49281
rect 27387 49160 29196 49235
rect 27387 49114 28810 49160
rect 28856 49117 29196 49160
rect 28856 49114 29116 49117
rect 27387 49071 29116 49114
rect 29162 49071 29196 49117
rect 27387 48997 29196 49071
rect 27387 48951 28810 48997
rect 28856 48954 29196 48997
rect 28856 48951 29116 48954
rect 27387 48908 29116 48951
rect 29162 48908 29196 48954
rect 27387 48834 29196 48908
rect 27387 48788 28810 48834
rect 28856 48788 29196 48834
rect 30583 49527 31040 49560
rect 34870 49553 35025 49560
rect 30583 49487 30855 49527
rect 30583 49441 30637 49487
rect 30683 49481 30855 49487
rect 30901 49481 31040 49527
rect 35294 49515 36266 49555
rect 37853 49549 38161 49557
rect 35294 49509 35332 49515
rect 35384 49509 35543 49515
rect 35595 49509 35754 49515
rect 35806 49509 35965 49515
rect 36017 49509 36176 49515
rect 36228 49509 36266 49515
rect 36438 49509 36953 49549
rect 37439 49517 38161 49549
rect 37439 49509 37891 49517
rect 37943 49509 38071 49517
rect 38123 49509 38161 49517
rect 38658 49509 39723 49569
rect 50099 49560 50408 49601
rect 52278 49653 54540 49694
rect 52278 49601 52316 49653
rect 52368 49601 52527 49653
rect 52579 49601 52738 49653
rect 52790 49601 52948 49653
rect 53000 49601 53159 49653
rect 53211 49601 53371 49653
rect 53423 49601 53582 49653
rect 53634 49601 53792 49653
rect 53844 49601 54003 49653
rect 54055 49601 54214 49653
rect 54266 49650 54540 49653
rect 54266 49604 54440 49650
rect 54486 49604 54540 49650
rect 54266 49601 54540 49604
rect 52278 49560 54540 49601
rect 54758 49653 55840 49694
rect 54758 49650 54855 49653
rect 54758 49604 54793 49650
rect 54839 49604 54855 49650
rect 54758 49601 54855 49604
rect 54907 49650 55066 49653
rect 54907 49604 54956 49650
rect 55002 49604 55066 49650
rect 54907 49601 55066 49604
rect 55118 49650 55278 49653
rect 55330 49650 55489 49653
rect 55164 49604 55278 49650
rect 55330 49604 55439 49650
rect 55485 49604 55489 49650
rect 55118 49601 55278 49604
rect 55330 49601 55489 49604
rect 55541 49650 55840 49653
rect 55541 49604 55599 49650
rect 55645 49604 55760 49650
rect 55806 49604 55840 49650
rect 55541 49601 55840 49604
rect 54758 49561 55840 49601
rect 55927 49653 57736 49767
rect 55927 49601 56015 49653
rect 56067 49601 56226 49653
rect 56278 49650 56437 49653
rect 56313 49604 56437 49650
rect 56278 49601 56437 49604
rect 56489 49601 56648 49653
rect 56700 49601 56859 49653
rect 56911 49601 57070 49653
rect 57122 49601 57281 49653
rect 57333 49601 57736 49653
rect 54817 49560 55579 49561
rect 48905 49515 49877 49555
rect 50099 49553 50255 49560
rect 48905 49509 48943 49515
rect 48995 49509 49154 49515
rect 49206 49509 49365 49515
rect 49417 49509 49576 49515
rect 49628 49509 49787 49515
rect 49839 49509 49877 49515
rect 30683 49441 31040 49481
rect 33484 49465 34643 49494
rect 30583 49364 31040 49441
rect 33019 49425 33327 49465
rect 33019 49422 33057 49425
rect 33109 49422 33237 49425
rect 33289 49422 33327 49425
rect 33484 49457 35082 49465
rect 35260 49463 35273 49509
rect 35523 49463 35543 49509
rect 35626 49463 35683 49509
rect 35729 49463 35754 49509
rect 35832 49463 35889 49509
rect 35935 49463 35965 49509
rect 36038 49463 36095 49509
rect 36141 49463 36176 49509
rect 36244 49463 36301 49509
rect 36347 49463 36360 49509
rect 36438 49463 36854 49509
rect 36900 49463 36971 49509
rect 37017 49463 37088 49509
rect 37134 49463 37206 49509
rect 37252 49463 37324 49509
rect 37370 49463 37442 49509
rect 37488 49465 37891 49509
rect 37488 49463 37909 49465
rect 37955 49463 38026 49509
rect 38123 49465 38143 49509
rect 38072 49463 38143 49465
rect 38189 49463 38261 49509
rect 38307 49463 38379 49509
rect 38425 49463 38497 49509
rect 38543 49463 38556 49509
rect 38658 49463 39021 49509
rect 39067 49463 39144 49509
rect 39190 49463 39267 49509
rect 39313 49463 39641 49509
rect 39687 49463 39730 49509
rect 31336 49376 31349 49422
rect 33323 49376 33336 49422
rect 33484 49411 33816 49457
rect 33862 49411 34002 49457
rect 34048 49411 34189 49457
rect 34235 49411 34376 49457
rect 34422 49411 34562 49457
rect 34608 49411 35082 49457
rect 35294 49423 36266 49463
rect 36438 49429 36953 49463
rect 37439 49429 38161 49463
rect 30583 49323 30855 49364
rect 30583 49277 30637 49323
rect 30683 49318 30855 49323
rect 30901 49318 31040 49364
rect 33019 49373 33057 49376
rect 33109 49373 33237 49376
rect 33289 49373 33327 49376
rect 33019 49332 33327 49373
rect 33484 49374 35082 49411
rect 30683 49277 31040 49318
rect 30583 49249 31040 49277
rect 33484 49292 33552 49374
rect 30583 49201 31493 49249
rect 30583 49160 30855 49201
rect 30583 49114 30637 49160
rect 30683 49155 30855 49160
rect 30901 49198 31493 49201
rect 30901 49155 31349 49198
rect 30683 49152 31349 49155
rect 33323 49152 33336 49198
rect 30683 49130 31493 49152
rect 30683 49114 31040 49130
rect 30583 49038 31040 49114
rect 30583 48997 30855 49038
rect 30583 48951 30637 48997
rect 30683 48992 30855 48997
rect 30901 48992 31040 49038
rect 30683 48951 31040 48992
rect 33019 48977 33327 49017
rect 33019 48974 33057 48977
rect 33109 48974 33237 48977
rect 33289 48974 33327 48977
rect 30583 48874 31040 48951
rect 31336 48928 31349 48974
rect 33323 48928 33336 48974
rect 33019 48925 33057 48928
rect 33109 48925 33237 48928
rect 33289 48925 33327 48928
rect 33019 48884 33327 48925
rect 30583 48834 30855 48874
rect 27387 48666 29196 48788
rect 27387 48620 28810 48666
rect 28856 48620 29196 48666
rect 29283 48753 30365 48794
rect 29283 48750 29582 48753
rect 29283 48704 29317 48750
rect 29363 48704 29478 48750
rect 29524 48704 29582 48750
rect 29283 48701 29582 48704
rect 29634 48750 29793 48753
rect 29845 48750 30005 48753
rect 29634 48704 29638 48750
rect 29684 48704 29793 48750
rect 29845 48704 29959 48750
rect 29634 48701 29793 48704
rect 29845 48701 30005 48704
rect 30057 48750 30216 48753
rect 30057 48704 30121 48750
rect 30167 48704 30216 48750
rect 30057 48701 30216 48704
rect 30268 48750 30365 48753
rect 30268 48704 30284 48750
rect 30330 48704 30365 48750
rect 30268 48701 30365 48704
rect 29283 48661 30365 48701
rect 30583 48788 30637 48834
rect 30683 48828 30855 48834
rect 30901 48828 31040 48874
rect 33484 48870 33495 49292
rect 33541 48870 33552 49292
rect 34964 49317 35082 49374
rect 36438 49329 36554 49429
rect 37853 49424 38161 49429
rect 38658 49449 39723 49463
rect 34964 49285 36360 49317
rect 34228 49215 34718 49256
rect 34228 49198 34267 49215
rect 34319 49198 34447 49215
rect 34499 49198 34627 49215
rect 33671 49152 33684 49198
rect 33730 49152 33787 49198
rect 33833 49152 33890 49198
rect 33936 49152 33993 49198
rect 34039 49152 34096 49198
rect 34142 49152 34199 49198
rect 34245 49163 34267 49198
rect 34245 49152 34302 49163
rect 34348 49152 34405 49198
rect 34499 49163 34508 49198
rect 34451 49152 34508 49163
rect 34554 49152 34612 49198
rect 34679 49163 34718 49215
rect 34964 49239 35273 49285
rect 35523 49239 35580 49285
rect 35626 49239 35683 49285
rect 35729 49239 35786 49285
rect 35832 49239 35889 49285
rect 35935 49239 35992 49285
rect 36038 49239 36095 49285
rect 36141 49239 36198 49285
rect 36244 49239 36301 49285
rect 36347 49239 36360 49285
rect 34964 49195 36360 49239
rect 34658 49152 34718 49163
rect 34228 49123 34718 49152
rect 36438 49189 36475 49329
rect 36521 49189 36554 49329
rect 35294 49061 36266 49095
rect 36438 49086 36554 49189
rect 36640 49329 36773 49349
rect 36640 49290 36697 49329
rect 36640 49238 36678 49290
rect 36640 49189 36697 49238
rect 36743 49189 36773 49329
rect 38658 49327 38726 49449
rect 39809 49443 44918 49481
rect 48765 49463 48778 49509
rect 48824 49463 48881 49509
rect 48927 49463 48943 49509
rect 49030 49463 49087 49509
rect 49133 49463 49154 49509
rect 49236 49463 49293 49509
rect 49339 49463 49365 49509
rect 49442 49463 49499 49509
rect 49545 49463 49576 49509
rect 49852 49463 49877 49509
rect 54085 49527 54540 49560
rect 50481 49467 51657 49494
rect 39809 49397 43739 49443
rect 43785 49397 43906 49443
rect 43952 49397 44071 49443
rect 44117 49397 44236 49443
rect 44282 49422 44918 49443
rect 48905 49423 49877 49463
rect 50044 49457 51657 49467
rect 44282 49397 44812 49422
rect 39809 49394 44812 49397
rect 39809 49348 39844 49394
rect 39890 49392 44812 49394
rect 39890 49348 39994 49392
rect 39809 49340 39994 49348
rect 40046 49376 44812 49392
rect 44858 49376 44925 49422
rect 44971 49376 45038 49422
rect 45084 49376 45151 49422
rect 45197 49376 45264 49422
rect 45310 49376 45323 49422
rect 48557 49377 48687 49417
rect 40046 49361 44918 49376
rect 40046 49340 40085 49361
rect 39809 49337 40085 49340
rect 36924 49317 37685 49324
rect 36923 49285 37931 49317
rect 36841 49239 36854 49285
rect 36900 49283 36971 49285
rect 36900 49239 36961 49283
rect 37017 49239 37088 49285
rect 37134 49283 37206 49285
rect 37134 49239 37172 49283
rect 37252 49239 37324 49285
rect 37370 49283 37442 49285
rect 37370 49239 37384 49283
rect 36923 49231 36961 49239
rect 37013 49231 37172 49239
rect 37224 49231 37384 49239
rect 37436 49239 37442 49283
rect 37488 49283 37909 49285
rect 37488 49239 37595 49283
rect 37436 49231 37595 49239
rect 37647 49239 37909 49283
rect 37955 49239 38026 49285
rect 38072 49239 38143 49285
rect 38189 49239 38261 49285
rect 38307 49239 38379 49285
rect 38425 49239 38497 49285
rect 38543 49239 38556 49285
rect 37647 49231 37931 49239
rect 36923 49198 37931 49231
rect 36923 49197 37685 49198
rect 36924 49191 37685 49197
rect 36640 49166 36773 49189
rect 38658 49187 38669 49327
rect 38715 49187 38726 49327
rect 39014 49285 39323 49317
rect 39492 49285 39608 49317
rect 39008 49239 39021 49285
rect 39067 49239 39144 49285
rect 39190 49239 39267 49285
rect 39313 49239 39326 49285
rect 39492 49239 39641 49285
rect 39687 49239 39730 49285
rect 38658 49176 38726 49187
rect 36438 49061 36953 49086
rect 37439 49083 37931 49086
rect 37439 49061 38161 49083
rect 35260 49015 35273 49061
rect 35523 49055 35580 49061
rect 35523 49015 35543 49055
rect 35626 49015 35683 49061
rect 35729 49055 35786 49061
rect 35729 49015 35754 49055
rect 35832 49015 35889 49061
rect 35935 49055 35992 49061
rect 35935 49015 35965 49055
rect 36038 49015 36095 49061
rect 36141 49055 36198 49061
rect 36141 49015 36176 49055
rect 36244 49015 36301 49061
rect 36347 49015 36360 49061
rect 36438 49015 36854 49061
rect 36900 49015 36971 49061
rect 37017 49015 37088 49061
rect 37134 49015 37206 49061
rect 37252 49015 37324 49061
rect 37370 49015 37442 49061
rect 37488 49043 37909 49061
rect 37488 49015 37891 49043
rect 37955 49015 38026 49061
rect 38072 49043 38143 49061
rect 38123 49015 38143 49043
rect 38189 49015 38261 49061
rect 38307 49015 38379 49061
rect 38425 49015 38497 49061
rect 38543 49015 38556 49061
rect 33781 48974 34089 49009
rect 35294 49003 35332 49015
rect 35384 49003 35543 49015
rect 35595 49003 35754 49015
rect 35806 49003 35965 49015
rect 36017 49003 36176 49015
rect 36228 49003 36266 49015
rect 33671 48928 33684 48974
rect 33730 48928 33787 48974
rect 33833 48969 33890 48974
rect 33871 48928 33890 48969
rect 33936 48928 33993 48974
rect 34039 48969 34096 48974
rect 34051 48928 34096 48969
rect 34142 48928 34199 48974
rect 34245 48928 34302 48974
rect 34348 48928 34405 48974
rect 34451 48928 34508 48974
rect 34554 48928 34612 48974
rect 34658 48928 34671 48974
rect 35294 48963 36266 49003
rect 36438 48966 36953 49015
rect 37439 48991 37891 49015
rect 37943 48991 38071 49015
rect 38123 48991 38161 49015
rect 37439 48966 38161 48991
rect 37853 48950 38161 48966
rect 33781 48917 33819 48928
rect 33871 48917 33999 48928
rect 34051 48917 34089 48928
rect 33781 48876 34089 48917
rect 33484 48859 33552 48870
rect 30683 48794 31040 48828
rect 30683 48788 32842 48794
rect 30583 48753 32842 48788
rect 34247 48787 35008 48794
rect 30583 48701 30854 48753
rect 30906 48701 31065 48753
rect 31117 48701 31276 48753
rect 31328 48750 31486 48753
rect 31538 48750 31697 48753
rect 31749 48750 31909 48753
rect 31961 48750 32120 48753
rect 32172 48750 32330 48753
rect 32382 48750 32541 48753
rect 32593 48750 32752 48753
rect 32804 48750 32842 48753
rect 34246 48753 35008 48787
rect 34246 48750 34284 48753
rect 34336 48750 34495 48753
rect 34547 48750 34707 48753
rect 31328 48704 31349 48750
rect 33323 48704 33336 48750
rect 33671 48704 33684 48750
rect 33730 48704 33787 48750
rect 33833 48704 33890 48750
rect 33936 48704 33993 48750
rect 34039 48704 34096 48750
rect 34142 48704 34199 48750
rect 34245 48704 34284 48750
rect 34348 48704 34405 48750
rect 34451 48704 34495 48750
rect 34554 48704 34612 48750
rect 34658 48704 34707 48750
rect 31328 48701 31486 48704
rect 31538 48701 31697 48704
rect 31749 48701 31909 48704
rect 31961 48701 32120 48704
rect 32172 48701 32330 48704
rect 32382 48701 32541 48704
rect 32593 48701 32752 48704
rect 32804 48701 32842 48704
rect 30583 48666 32842 48701
rect 34246 48701 34284 48704
rect 34336 48701 34495 48704
rect 34547 48701 34707 48704
rect 34759 48701 34918 48753
rect 34970 48701 35008 48753
rect 34246 48667 35008 48701
rect 29544 48660 30306 48661
rect 27387 48544 29196 48620
rect 27387 48503 29116 48544
rect 27387 48457 28810 48503
rect 28856 48498 29116 48503
rect 29162 48498 29196 48544
rect 28856 48457 29196 48498
rect 27387 48381 29196 48457
rect 27387 48340 29116 48381
rect 27387 48294 28810 48340
rect 28856 48335 29116 48340
rect 29162 48335 29196 48381
rect 28856 48294 29196 48335
rect 27387 48217 29196 48294
rect 27387 48177 29116 48217
rect 27387 48131 28810 48177
rect 28856 48171 29116 48177
rect 29162 48171 29196 48217
rect 28856 48131 29196 48171
rect 27387 48054 29196 48131
rect 27387 48013 29116 48054
rect 27387 47967 28810 48013
rect 28856 48008 29116 48013
rect 29162 48008 29196 48054
rect 28856 47967 29196 48008
rect 27387 47853 29196 47967
rect 30583 48620 30637 48666
rect 30683 48660 32842 48666
rect 34247 48660 35008 48667
rect 35182 48787 36364 48794
rect 35182 48753 36958 48787
rect 35182 48701 35220 48753
rect 35272 48701 35430 48753
rect 35482 48701 35641 48753
rect 35693 48701 35853 48753
rect 35905 48701 36064 48753
rect 36116 48701 36274 48753
rect 36326 48750 36958 48753
rect 36326 48704 36489 48750
rect 36723 48704 36958 48750
rect 36326 48701 36958 48704
rect 35182 48667 36958 48701
rect 37946 48753 38842 48794
rect 37946 48750 38330 48753
rect 38382 48750 38541 48753
rect 37946 48704 37957 48750
rect 38473 48704 38541 48750
rect 37946 48701 38330 48704
rect 38382 48701 38541 48704
rect 38593 48701 38752 48753
rect 38804 48701 38842 48753
rect 35182 48660 36364 48667
rect 37946 48660 38842 48701
rect 39014 48753 39323 49239
rect 39014 48701 39052 48753
rect 39104 48750 39232 48753
rect 39108 48704 39220 48750
rect 39104 48701 39232 48704
rect 39284 48701 39323 48753
rect 30683 48626 31040 48660
rect 30683 48620 30855 48626
rect 30583 48580 30855 48620
rect 30901 48580 31040 48626
rect 30583 48503 31040 48580
rect 33484 48584 33552 48595
rect 33019 48529 33327 48570
rect 33019 48526 33057 48529
rect 33109 48526 33237 48529
rect 33289 48526 33327 48529
rect 30583 48457 30637 48503
rect 30683 48462 31040 48503
rect 31336 48480 31349 48526
rect 33323 48480 33336 48526
rect 30683 48457 30855 48462
rect 30583 48416 30855 48457
rect 30901 48416 31040 48462
rect 33019 48477 33057 48480
rect 33109 48477 33237 48480
rect 33289 48477 33327 48480
rect 33019 48437 33327 48477
rect 30583 48340 31040 48416
rect 30583 48294 30637 48340
rect 30683 48324 31040 48340
rect 30683 48302 31493 48324
rect 30683 48299 31349 48302
rect 30683 48294 30855 48299
rect 30583 48253 30855 48294
rect 30901 48256 31349 48299
rect 33323 48256 33336 48302
rect 30901 48253 31493 48256
rect 30583 48205 31493 48253
rect 30583 48177 31040 48205
rect 30583 48131 30637 48177
rect 30683 48136 31040 48177
rect 30683 48131 30855 48136
rect 30583 48090 30855 48131
rect 30901 48090 31040 48136
rect 33484 48162 33495 48584
rect 33541 48162 33552 48584
rect 33781 48537 34089 48578
rect 33781 48526 33819 48537
rect 33871 48526 33999 48537
rect 34051 48526 34089 48537
rect 33671 48480 33684 48526
rect 33730 48480 33787 48526
rect 33871 48485 33890 48526
rect 33833 48480 33890 48485
rect 33936 48480 33993 48526
rect 34051 48485 34096 48526
rect 34039 48480 34096 48485
rect 34142 48480 34199 48526
rect 34245 48480 34302 48526
rect 34348 48480 34405 48526
rect 34451 48480 34508 48526
rect 34554 48480 34612 48526
rect 34658 48480 34671 48526
rect 33781 48445 34089 48480
rect 35294 48451 36266 48491
rect 37853 48488 38161 48504
rect 35294 48439 35332 48451
rect 35384 48439 35543 48451
rect 35595 48439 35754 48451
rect 35806 48439 35965 48451
rect 36017 48439 36176 48451
rect 36228 48439 36266 48451
rect 36438 48439 36953 48488
rect 37439 48463 38161 48488
rect 37439 48439 37891 48463
rect 37943 48439 38071 48463
rect 38123 48439 38161 48463
rect 35260 48393 35273 48439
rect 35523 48399 35543 48439
rect 35523 48393 35580 48399
rect 35626 48393 35683 48439
rect 35729 48399 35754 48439
rect 35729 48393 35786 48399
rect 35832 48393 35889 48439
rect 35935 48399 35965 48439
rect 35935 48393 35992 48399
rect 36038 48393 36095 48439
rect 36141 48399 36176 48439
rect 36141 48393 36198 48399
rect 36244 48393 36301 48439
rect 36347 48393 36360 48439
rect 36438 48393 36854 48439
rect 36900 48393 36971 48439
rect 37017 48393 37088 48439
rect 37134 48393 37206 48439
rect 37252 48393 37324 48439
rect 37370 48393 37442 48439
rect 37488 48411 37891 48439
rect 37488 48393 37909 48411
rect 37955 48393 38026 48439
rect 38123 48411 38143 48439
rect 38072 48393 38143 48411
rect 38189 48393 38261 48439
rect 38307 48393 38379 48439
rect 38425 48393 38497 48439
rect 38543 48393 38556 48439
rect 35294 48359 36266 48393
rect 36438 48368 36953 48393
rect 37439 48371 38161 48393
rect 37439 48368 37931 48371
rect 34228 48302 34718 48331
rect 33671 48256 33684 48302
rect 33730 48256 33787 48302
rect 33833 48256 33890 48302
rect 33936 48256 33993 48302
rect 34039 48256 34096 48302
rect 34142 48256 34199 48302
rect 34245 48291 34302 48302
rect 34245 48256 34267 48291
rect 34348 48256 34405 48302
rect 34451 48291 34508 48302
rect 34499 48256 34508 48291
rect 34554 48256 34612 48302
rect 34658 48291 34718 48302
rect 34228 48239 34267 48256
rect 34319 48239 34447 48256
rect 34499 48239 34627 48256
rect 34679 48239 34718 48291
rect 36438 48265 36554 48368
rect 34228 48198 34718 48239
rect 34964 48215 36360 48259
rect 30583 48013 31040 48090
rect 33019 48081 33327 48122
rect 33019 48078 33057 48081
rect 33109 48078 33237 48081
rect 33289 48078 33327 48081
rect 33484 48080 33552 48162
rect 34964 48169 35273 48215
rect 35523 48169 35580 48215
rect 35626 48169 35683 48215
rect 35729 48169 35786 48215
rect 35832 48169 35889 48215
rect 35935 48169 35992 48215
rect 36038 48169 36095 48215
rect 36141 48169 36198 48215
rect 36244 48169 36301 48215
rect 36347 48169 36360 48215
rect 34964 48137 36360 48169
rect 34964 48080 35082 48137
rect 31336 48032 31349 48078
rect 33323 48032 33336 48078
rect 33484 48043 35082 48080
rect 30583 47967 30637 48013
rect 30683 47973 31040 48013
rect 33019 48029 33057 48032
rect 33109 48029 33237 48032
rect 33289 48029 33327 48032
rect 33019 47989 33327 48029
rect 33484 47997 33816 48043
rect 33862 47997 34002 48043
rect 34048 47997 34189 48043
rect 34235 47997 34376 48043
rect 34422 47997 34562 48043
rect 34608 47997 35082 48043
rect 36438 48125 36475 48265
rect 36521 48125 36554 48265
rect 33484 47989 35082 47997
rect 35294 47991 36266 48031
rect 36438 48025 36554 48125
rect 36640 48265 36773 48288
rect 36640 48216 36697 48265
rect 36640 48164 36678 48216
rect 36640 48125 36697 48164
rect 36743 48125 36773 48265
rect 38658 48267 38726 48278
rect 36924 48257 37685 48263
rect 36923 48256 37685 48257
rect 36923 48223 37931 48256
rect 36923 48215 36961 48223
rect 37013 48215 37172 48223
rect 37224 48215 37384 48223
rect 36841 48169 36854 48215
rect 36900 48171 36961 48215
rect 36900 48169 36971 48171
rect 37017 48169 37088 48215
rect 37134 48171 37172 48215
rect 37134 48169 37206 48171
rect 37252 48169 37324 48215
rect 37370 48171 37384 48215
rect 37436 48215 37595 48223
rect 37436 48171 37442 48215
rect 37370 48169 37442 48171
rect 37488 48171 37595 48215
rect 37647 48215 37931 48223
rect 37647 48171 37909 48215
rect 37488 48169 37909 48171
rect 37955 48169 38026 48215
rect 38072 48169 38143 48215
rect 38189 48169 38261 48215
rect 38307 48169 38379 48215
rect 38425 48169 38497 48215
rect 38543 48169 38556 48215
rect 36923 48137 37931 48169
rect 36924 48130 37685 48137
rect 36640 48105 36773 48125
rect 38658 48127 38669 48267
rect 38715 48127 38726 48267
rect 39014 48215 39323 48701
rect 39492 48787 39608 49239
rect 39923 49206 40085 49337
rect 39923 49154 39994 49206
rect 40046 49154 40085 49206
rect 39923 49114 40085 49154
rect 39737 49018 39865 49031
rect 39737 48991 39866 49018
rect 39737 48974 39775 48991
rect 39827 48974 39866 48991
rect 39727 48928 39740 48974
rect 39827 48939 39862 48974
rect 39786 48928 39862 48939
rect 39908 48928 39985 48974
rect 40031 48928 40108 48974
rect 40154 48928 40167 48974
rect 40246 48963 40362 49361
rect 42229 49222 44509 49263
rect 42229 49170 43068 49222
rect 43120 49170 44509 49222
rect 42229 49130 44509 49170
rect 44341 49086 44509 49130
rect 44341 49040 44358 49086
rect 44498 49040 44509 49086
rect 39737 48899 39866 48928
rect 40246 48917 40281 48963
rect 40327 48917 40362 48963
rect 40246 48880 40362 48917
rect 40718 48991 43524 49032
rect 44341 49029 44509 49040
rect 40718 48939 41935 48991
rect 41987 48939 43524 48991
rect 40718 48898 43524 48939
rect 44605 48974 44721 49361
rect 45400 49331 48379 49372
rect 45400 49317 45975 49331
rect 45400 49271 45464 49317
rect 45604 49279 45975 49317
rect 46027 49279 48379 49331
rect 45604 49271 48379 49279
rect 44901 49215 45241 49256
rect 45400 49238 48379 49271
rect 48557 49325 48596 49377
rect 48648 49325 48687 49377
rect 48557 49302 48687 49325
rect 50044 49411 50516 49457
rect 50562 49411 50703 49457
rect 50749 49411 50890 49457
rect 50936 49411 51076 49457
rect 51122 49411 51263 49457
rect 51309 49411 51657 49457
rect 51797 49447 52105 49487
rect 51797 49422 51835 49447
rect 51887 49422 52015 49447
rect 52067 49422 52105 49447
rect 54085 49481 54223 49527
rect 54269 49487 54540 49527
rect 54269 49481 54440 49487
rect 54085 49441 54440 49481
rect 54486 49441 54540 49487
rect 50044 49374 51657 49411
rect 51789 49376 51802 49422
rect 53776 49376 53789 49422
rect 50044 49317 50160 49374
rect 44901 49198 44939 49215
rect 44991 49198 45151 49215
rect 45203 49198 45241 49215
rect 44799 49152 44812 49198
rect 44858 49152 44925 49198
rect 44991 49163 45038 49198
rect 44971 49152 45038 49163
rect 45084 49152 45151 49198
rect 45203 49163 45264 49198
rect 45197 49152 45264 49163
rect 45310 49152 45323 49198
rect 48557 49162 48622 49302
rect 48668 49162 48687 49302
rect 49820 49285 50160 49317
rect 48765 49239 48778 49285
rect 48824 49239 48881 49285
rect 48927 49239 48984 49285
rect 49030 49239 49087 49285
rect 49133 49239 49190 49285
rect 49236 49239 49293 49285
rect 49339 49239 49396 49285
rect 49442 49239 49499 49285
rect 49545 49239 49602 49285
rect 49852 49239 50160 49285
rect 51589 49322 51657 49374
rect 51797 49354 52105 49376
rect 49820 49198 50160 49239
rect 50262 49215 50812 49256
rect 48557 49159 48687 49162
rect 44901 49123 45241 49152
rect 48557 49107 48596 49159
rect 48648 49107 48687 49159
rect 50262 49163 50300 49215
rect 50352 49198 50511 49215
rect 50563 49198 50722 49215
rect 50352 49163 50467 49198
rect 50563 49163 50571 49198
rect 50262 49152 50467 49163
rect 50513 49152 50571 49163
rect 50617 49152 50674 49198
rect 50720 49163 50722 49198
rect 50774 49198 50812 49215
rect 50774 49163 50777 49198
rect 50720 49152 50777 49163
rect 50823 49152 50880 49198
rect 50926 49152 50983 49198
rect 51029 49152 51086 49198
rect 51132 49152 51189 49198
rect 51235 49152 51292 49198
rect 51338 49152 51395 49198
rect 51441 49152 51454 49198
rect 50262 49123 50812 49152
rect 48557 49066 48687 49107
rect 48905 49061 49877 49092
rect 48765 49015 48778 49061
rect 48824 49015 48881 49061
rect 48927 49052 48984 49061
rect 48927 49015 48943 49052
rect 49030 49015 49087 49061
rect 49133 49052 49190 49061
rect 49133 49015 49154 49052
rect 49236 49015 49293 49061
rect 49339 49052 49396 49061
rect 49339 49015 49365 49052
rect 49442 49015 49499 49061
rect 49545 49052 49602 49061
rect 49545 49015 49576 49052
rect 49852 49015 49877 49061
rect 48905 49000 48943 49015
rect 48995 49000 49154 49015
rect 49206 49000 49365 49015
rect 49417 49000 49576 49015
rect 49628 49000 49787 49015
rect 49839 49000 49877 49015
rect 44605 48928 44812 48974
rect 44858 48928 44925 48974
rect 44971 48928 45038 48974
rect 45084 48928 45151 48974
rect 45197 48928 45264 48974
rect 45310 48928 45323 48974
rect 48905 48960 49877 49000
rect 51035 48977 51343 49017
rect 51035 48974 51073 48977
rect 51125 48974 51253 48977
rect 51305 48974 51343 48977
rect 43362 48891 43524 48898
rect 43362 48845 43373 48891
rect 43513 48845 43524 48891
rect 43362 48834 43524 48845
rect 45584 48914 48546 48950
rect 50454 48928 50467 48974
rect 50513 48928 50571 48974
rect 50617 48928 50674 48974
rect 50720 48928 50777 48974
rect 50823 48928 50880 48974
rect 50926 48928 50983 48974
rect 51029 48928 51073 48974
rect 51132 48928 51189 48974
rect 51235 48928 51253 48974
rect 51338 48928 51395 48974
rect 51441 48928 51454 48974
rect 45584 48868 45619 48914
rect 45665 48868 45777 48914
rect 45823 48868 45935 48914
rect 45981 48868 46093 48914
rect 46139 48868 46251 48914
rect 46297 48868 46409 48914
rect 46455 48868 46568 48914
rect 46614 48868 46726 48914
rect 46772 48868 46884 48914
rect 46930 48868 47042 48914
rect 47088 48868 47200 48914
rect 47246 48868 47358 48914
rect 47404 48868 47516 48914
rect 47562 48868 47675 48914
rect 47721 48868 47833 48914
rect 47879 48868 47991 48914
rect 48037 48868 48149 48914
rect 48195 48868 48307 48914
rect 48353 48868 48465 48914
rect 48511 48868 48546 48914
rect 51035 48925 51073 48928
rect 51125 48925 51253 48928
rect 51305 48925 51343 48928
rect 51035 48884 51343 48925
rect 51589 48900 51600 49322
rect 51646 48900 51657 49322
rect 54085 49323 54540 49441
rect 54085 49277 54440 49323
rect 54486 49277 54540 49323
rect 54085 49249 54540 49277
rect 53585 49198 54540 49249
rect 51789 49152 51802 49198
rect 53776 49160 54540 49198
rect 53776 49152 54440 49160
rect 53585 49130 54440 49152
rect 54085 49114 54440 49130
rect 54486 49114 54540 49160
rect 54085 49038 54540 49114
rect 51797 48984 52105 49024
rect 51797 48974 51835 48984
rect 51887 48974 52015 48984
rect 52067 48974 52105 48984
rect 54085 48992 54223 49038
rect 54269 48997 54540 49038
rect 54269 48992 54440 48997
rect 51789 48928 51802 48974
rect 53776 48928 53789 48974
rect 54085 48951 54440 48992
rect 54486 48951 54540 48997
rect 51589 48889 51657 48900
rect 51797 48891 52105 48928
rect 40215 48787 40523 48794
rect 40788 48787 42986 48801
rect 43753 48787 44514 48794
rect 39492 48764 42986 48787
rect 43704 48764 44514 48787
rect 39492 48753 44514 48764
rect 39492 48750 40253 48753
rect 39492 48704 39740 48750
rect 39786 48704 39862 48750
rect 39908 48704 39985 48750
rect 40031 48704 40108 48750
rect 40154 48704 40253 48750
rect 39492 48701 40253 48704
rect 40305 48701 40433 48753
rect 40485 48750 43790 48753
rect 40485 48704 40836 48750
rect 40882 48704 40994 48750
rect 41040 48704 41152 48750
rect 41198 48704 41310 48750
rect 41356 48704 41469 48750
rect 41515 48704 41627 48750
rect 41673 48704 41785 48750
rect 41831 48704 41943 48750
rect 41989 48704 42101 48750
rect 42147 48704 42259 48750
rect 42305 48704 42418 48750
rect 42464 48704 42576 48750
rect 42622 48704 42734 48750
rect 42780 48704 42892 48750
rect 42938 48704 43739 48750
rect 43785 48704 43790 48750
rect 40485 48701 43790 48704
rect 43842 48750 44001 48753
rect 43842 48704 43906 48750
rect 43952 48704 44001 48750
rect 43842 48701 44001 48704
rect 44053 48750 44213 48753
rect 44265 48750 44424 48753
rect 44053 48704 44071 48750
rect 44117 48704 44213 48750
rect 44282 48704 44424 48750
rect 44053 48701 44213 48704
rect 44265 48701 44424 48704
rect 44476 48701 44514 48753
rect 39492 48690 44514 48701
rect 39492 48667 42986 48690
rect 43704 48667 44514 48690
rect 39492 48215 39608 48667
rect 40215 48660 40523 48667
rect 40788 48653 42986 48667
rect 43753 48660 44514 48667
rect 44796 48787 45346 48794
rect 45584 48787 48546 48868
rect 54085 48874 54540 48951
rect 54085 48828 54223 48874
rect 54269 48834 54540 48874
rect 54269 48828 54440 48834
rect 54085 48794 54440 48828
rect 48800 48787 49982 48794
rect 50308 48787 50859 48794
rect 44796 48753 49982 48787
rect 44796 48750 44834 48753
rect 44886 48750 45045 48753
rect 45097 48750 45256 48753
rect 45308 48750 48838 48753
rect 44796 48704 44812 48750
rect 44886 48704 44925 48750
rect 44971 48704 45038 48750
rect 45097 48704 45151 48750
rect 45197 48704 45256 48750
rect 45310 48704 45619 48750
rect 45665 48704 45777 48750
rect 45823 48704 45935 48750
rect 45981 48704 46093 48750
rect 46139 48704 46251 48750
rect 46297 48704 46409 48750
rect 46455 48704 46568 48750
rect 46614 48704 46726 48750
rect 46772 48704 46884 48750
rect 46930 48704 47042 48750
rect 47088 48704 47200 48750
rect 47246 48704 47358 48750
rect 47404 48704 47516 48750
rect 47562 48704 47675 48750
rect 47721 48704 47833 48750
rect 47879 48704 47991 48750
rect 48037 48704 48149 48750
rect 48195 48704 48307 48750
rect 48353 48704 48465 48750
rect 48511 48704 48838 48750
rect 44796 48701 44834 48704
rect 44886 48701 45045 48704
rect 45097 48701 45256 48704
rect 45308 48701 48838 48704
rect 48890 48701 49048 48753
rect 49100 48701 49259 48753
rect 49311 48701 49471 48753
rect 49523 48701 49682 48753
rect 49734 48701 49892 48753
rect 49944 48701 49982 48753
rect 44796 48667 49982 48701
rect 50307 48753 50859 48787
rect 50307 48701 50346 48753
rect 50398 48750 50557 48753
rect 50609 48750 50768 48753
rect 50820 48750 50859 48753
rect 52278 48788 54440 48794
rect 54486 48788 54540 48834
rect 55927 49487 57736 49601
rect 55927 49444 56267 49487
rect 55927 49398 55961 49444
rect 56007 49441 56267 49444
rect 56313 49441 57736 49487
rect 56007 49398 57736 49441
rect 55927 49323 57736 49398
rect 55927 49281 56267 49323
rect 55927 49235 55961 49281
rect 56007 49277 56267 49281
rect 56313 49277 57736 49323
rect 56007 49235 57736 49277
rect 55927 49160 57736 49235
rect 55927 49117 56267 49160
rect 55927 49071 55961 49117
rect 56007 49114 56267 49117
rect 56313 49114 57736 49160
rect 56007 49071 57736 49114
rect 55927 48997 57736 49071
rect 55927 48954 56267 48997
rect 55927 48908 55961 48954
rect 56007 48951 56267 48954
rect 56313 48951 57736 48997
rect 56007 48908 57736 48951
rect 55927 48834 57736 48908
rect 52278 48753 54540 48788
rect 52278 48750 52316 48753
rect 52368 48750 52527 48753
rect 52579 48750 52738 48753
rect 52790 48750 52948 48753
rect 53000 48750 53159 48753
rect 53211 48750 53371 48753
rect 53423 48750 53582 48753
rect 53634 48750 53792 48753
rect 50398 48704 50467 48750
rect 50513 48704 50557 48750
rect 50617 48704 50674 48750
rect 50720 48704 50768 48750
rect 50823 48704 50880 48750
rect 50926 48704 50983 48750
rect 51029 48704 51086 48750
rect 51132 48704 51189 48750
rect 51235 48704 51292 48750
rect 51338 48704 51395 48750
rect 51441 48704 51454 48750
rect 51789 48704 51802 48750
rect 53776 48704 53792 48750
rect 50398 48701 50557 48704
rect 50609 48701 50768 48704
rect 50820 48701 50859 48704
rect 50307 48667 50859 48701
rect 44796 48660 45346 48667
rect 43362 48609 43524 48620
rect 39737 48526 39866 48555
rect 40246 48537 40362 48574
rect 43362 48563 43373 48609
rect 43513 48563 43524 48609
rect 43362 48556 43524 48563
rect 39727 48480 39740 48526
rect 39786 48515 39862 48526
rect 39827 48480 39862 48515
rect 39908 48480 39985 48526
rect 40031 48480 40108 48526
rect 40154 48480 40167 48526
rect 40246 48491 40281 48537
rect 40327 48491 40362 48537
rect 39737 48463 39775 48480
rect 39827 48463 39866 48480
rect 39737 48436 39866 48463
rect 39737 48423 39865 48436
rect 39923 48300 40085 48340
rect 39923 48248 39994 48300
rect 40046 48248 40085 48300
rect 39008 48169 39021 48215
rect 39067 48169 39144 48215
rect 39190 48169 39267 48215
rect 39313 48169 39326 48215
rect 39492 48169 39641 48215
rect 39687 48169 39730 48215
rect 39014 48137 39323 48169
rect 39492 48137 39608 48169
rect 37853 48025 38161 48030
rect 36438 47991 36953 48025
rect 37439 47991 38161 48025
rect 38658 48005 38726 48127
rect 39923 48117 40085 48248
rect 39809 48114 40085 48117
rect 39809 48106 39994 48114
rect 39809 48060 39844 48106
rect 39890 48062 39994 48106
rect 40046 48093 40085 48114
rect 40246 48093 40362 48491
rect 40718 48515 43524 48556
rect 45584 48586 48546 48667
rect 48800 48660 49982 48667
rect 50308 48660 50859 48667
rect 52278 48701 52316 48704
rect 52368 48701 52527 48704
rect 52579 48701 52738 48704
rect 52790 48701 52948 48704
rect 53000 48701 53159 48704
rect 53211 48701 53371 48704
rect 53423 48701 53582 48704
rect 53634 48701 53792 48704
rect 53844 48701 54003 48753
rect 54055 48701 54214 48753
rect 54266 48701 54540 48753
rect 52278 48666 54540 48701
rect 52278 48660 54440 48666
rect 45584 48540 45619 48586
rect 45665 48540 45777 48586
rect 45823 48540 45935 48586
rect 45981 48540 46093 48586
rect 46139 48540 46251 48586
rect 46297 48540 46409 48586
rect 46455 48540 46568 48586
rect 46614 48540 46726 48586
rect 46772 48540 46884 48586
rect 46930 48540 47042 48586
rect 47088 48540 47200 48586
rect 47246 48540 47358 48586
rect 47404 48540 47516 48586
rect 47562 48540 47675 48586
rect 47721 48540 47833 48586
rect 47879 48540 47991 48586
rect 48037 48540 48149 48586
rect 48195 48540 48307 48586
rect 48353 48540 48465 48586
rect 48511 48540 48546 48586
rect 54085 48626 54440 48660
rect 54085 48580 54223 48626
rect 54269 48620 54440 48626
rect 54486 48620 54540 48666
rect 54758 48753 55840 48794
rect 54758 48750 54855 48753
rect 54758 48704 54793 48750
rect 54839 48704 54855 48750
rect 54758 48701 54855 48704
rect 54907 48750 55066 48753
rect 54907 48704 54956 48750
rect 55002 48704 55066 48750
rect 54907 48701 55066 48704
rect 55118 48750 55278 48753
rect 55330 48750 55489 48753
rect 55164 48704 55278 48750
rect 55330 48704 55439 48750
rect 55485 48704 55489 48750
rect 55118 48701 55278 48704
rect 55330 48701 55489 48704
rect 55541 48750 55840 48753
rect 55541 48704 55599 48750
rect 55645 48704 55760 48750
rect 55806 48704 55840 48750
rect 55541 48701 55840 48704
rect 54758 48661 55840 48701
rect 55927 48788 56267 48834
rect 56313 48788 57736 48834
rect 55927 48666 57736 48788
rect 54817 48660 55579 48661
rect 54269 48580 54540 48620
rect 40718 48463 41935 48515
rect 41987 48463 43524 48515
rect 40718 48422 43524 48463
rect 44605 48480 44812 48526
rect 44858 48480 44925 48526
rect 44971 48480 45038 48526
rect 45084 48480 45151 48526
rect 45197 48480 45264 48526
rect 45310 48480 45323 48526
rect 45584 48504 48546 48540
rect 51035 48529 51343 48570
rect 51035 48526 51073 48529
rect 51125 48526 51253 48529
rect 51305 48526 51343 48529
rect 51589 48554 51657 48565
rect 44341 48414 44509 48425
rect 44341 48368 44358 48414
rect 44498 48368 44509 48414
rect 44341 48324 44509 48368
rect 42229 48284 44509 48324
rect 42229 48232 43068 48284
rect 43120 48232 44509 48284
rect 42229 48191 44509 48232
rect 44605 48093 44721 48480
rect 48905 48454 49877 48494
rect 50454 48480 50467 48526
rect 50513 48480 50571 48526
rect 50617 48480 50674 48526
rect 50720 48480 50777 48526
rect 50823 48480 50880 48526
rect 50926 48480 50983 48526
rect 51029 48480 51073 48526
rect 51132 48480 51189 48526
rect 51235 48480 51253 48526
rect 51338 48480 51395 48526
rect 51441 48480 51454 48526
rect 48905 48439 48943 48454
rect 48995 48439 49154 48454
rect 49206 48439 49365 48454
rect 49417 48439 49576 48454
rect 49628 48439 49787 48454
rect 49839 48439 49877 48454
rect 48765 48393 48778 48439
rect 48824 48393 48881 48439
rect 48927 48402 48943 48439
rect 48927 48393 48984 48402
rect 49030 48393 49087 48439
rect 49133 48402 49154 48439
rect 49133 48393 49190 48402
rect 49236 48393 49293 48439
rect 49339 48402 49365 48439
rect 49339 48393 49396 48402
rect 49442 48393 49499 48439
rect 49545 48402 49576 48439
rect 49545 48393 49602 48402
rect 49852 48393 49877 48439
rect 51035 48477 51073 48480
rect 51125 48477 51253 48480
rect 51305 48477 51343 48480
rect 51035 48437 51343 48477
rect 48557 48347 48687 48388
rect 48905 48362 49877 48393
rect 44901 48302 45241 48331
rect 44799 48256 44812 48302
rect 44858 48256 44925 48302
rect 44971 48291 45038 48302
rect 44991 48256 45038 48291
rect 45084 48256 45151 48302
rect 45197 48291 45264 48302
rect 45203 48256 45264 48291
rect 45310 48256 45323 48302
rect 48557 48295 48596 48347
rect 48648 48295 48687 48347
rect 48557 48292 48687 48295
rect 44901 48239 44939 48256
rect 44991 48239 45151 48256
rect 45203 48239 45241 48256
rect 44901 48198 45241 48239
rect 45400 48183 48379 48216
rect 45400 48137 45464 48183
rect 45604 48175 48379 48183
rect 45604 48137 46353 48175
rect 45400 48123 46353 48137
rect 46405 48123 48379 48175
rect 40046 48078 44918 48093
rect 45400 48082 48379 48123
rect 48557 48152 48622 48292
rect 48668 48152 48687 48292
rect 50262 48302 50812 48331
rect 50262 48291 50467 48302
rect 50513 48291 50571 48302
rect 49820 48215 50160 48256
rect 48765 48169 48778 48215
rect 48824 48169 48881 48215
rect 48927 48169 48984 48215
rect 49030 48169 49087 48215
rect 49133 48169 49190 48215
rect 49236 48169 49293 48215
rect 49339 48169 49396 48215
rect 49442 48169 49499 48215
rect 49545 48169 49602 48215
rect 49852 48169 50160 48215
rect 50262 48239 50300 48291
rect 50352 48256 50467 48291
rect 50563 48256 50571 48291
rect 50617 48256 50674 48302
rect 50720 48291 50777 48302
rect 50720 48256 50722 48291
rect 50352 48239 50511 48256
rect 50563 48239 50722 48256
rect 50774 48256 50777 48291
rect 50823 48256 50880 48302
rect 50926 48256 50983 48302
rect 51029 48256 51086 48302
rect 51132 48256 51189 48302
rect 51235 48256 51292 48302
rect 51338 48256 51395 48302
rect 51441 48256 51454 48302
rect 50774 48239 50812 48256
rect 50262 48198 50812 48239
rect 48557 48129 48687 48152
rect 49820 48137 50160 48169
rect 40046 48062 44812 48078
rect 39890 48060 44812 48062
rect 39809 48057 44812 48060
rect 39809 48011 43739 48057
rect 43785 48011 43906 48057
rect 43952 48011 44071 48057
rect 44117 48011 44236 48057
rect 44282 48032 44812 48057
rect 44858 48032 44925 48078
rect 44971 48032 45038 48078
rect 45084 48032 45151 48078
rect 45197 48032 45264 48078
rect 45310 48032 45323 48078
rect 48557 48077 48596 48129
rect 48648 48077 48687 48129
rect 48557 48037 48687 48077
rect 50044 48080 50160 48137
rect 51589 48132 51600 48554
rect 51646 48132 51657 48554
rect 51797 48526 52105 48563
rect 51789 48480 51802 48526
rect 53776 48480 53789 48526
rect 54085 48503 54540 48580
rect 51797 48470 51835 48480
rect 51887 48470 52015 48480
rect 52067 48470 52105 48480
rect 51797 48430 52105 48470
rect 54085 48462 54440 48503
rect 54085 48416 54223 48462
rect 54269 48457 54440 48462
rect 54486 48457 54540 48503
rect 54269 48416 54540 48457
rect 54085 48340 54540 48416
rect 54085 48324 54440 48340
rect 53585 48302 54440 48324
rect 51789 48256 51802 48302
rect 53776 48294 54440 48302
rect 54486 48294 54540 48340
rect 53776 48256 54540 48294
rect 53585 48205 54540 48256
rect 51589 48080 51657 48132
rect 54085 48177 54540 48205
rect 54085 48131 54440 48177
rect 54486 48131 54540 48177
rect 50044 48043 51657 48080
rect 51797 48078 52105 48100
rect 44282 48011 44918 48032
rect 38658 47991 39723 48005
rect 30683 47967 30855 47973
rect 30583 47927 30855 47967
rect 30901 47927 31040 47973
rect 33484 47960 34643 47989
rect 35260 47945 35273 47991
rect 35523 47945 35543 47991
rect 35626 47945 35683 47991
rect 35729 47945 35754 47991
rect 35832 47945 35889 47991
rect 35935 47945 35965 47991
rect 36038 47945 36095 47991
rect 36141 47945 36176 47991
rect 36244 47945 36301 47991
rect 36347 47945 36360 47991
rect 36438 47945 36854 47991
rect 36900 47945 36971 47991
rect 37017 47945 37088 47991
rect 37134 47945 37206 47991
rect 37252 47945 37324 47991
rect 37370 47945 37442 47991
rect 37488 47989 37909 47991
rect 37488 47945 37891 47989
rect 37955 47945 38026 47991
rect 38072 47989 38143 47991
rect 38123 47945 38143 47989
rect 38189 47945 38261 47991
rect 38307 47945 38379 47991
rect 38425 47945 38497 47991
rect 38543 47945 38556 47991
rect 38658 47945 39021 47991
rect 39067 47945 39144 47991
rect 39190 47945 39267 47991
rect 39313 47945 39641 47991
rect 39687 47945 39730 47991
rect 39809 47973 44918 48011
rect 48905 47991 49877 48031
rect 48765 47945 48778 47991
rect 48824 47945 48881 47991
rect 48927 47945 48943 47991
rect 49030 47945 49087 47991
rect 49133 47945 49154 47991
rect 49236 47945 49293 47991
rect 49339 47945 49365 47991
rect 49442 47945 49499 47991
rect 49545 47945 49576 47991
rect 49852 47945 49877 47991
rect 50044 47997 50516 48043
rect 50562 47997 50703 48043
rect 50749 47997 50890 48043
rect 50936 47997 51076 48043
rect 51122 47997 51263 48043
rect 51309 47997 51657 48043
rect 51789 48032 51802 48078
rect 53776 48032 53789 48078
rect 50044 47987 51657 47997
rect 50481 47960 51657 47987
rect 51797 48007 51835 48032
rect 51887 48007 52015 48032
rect 52067 48007 52105 48032
rect 51797 47967 52105 48007
rect 54085 48013 54540 48131
rect 54085 47973 54440 48013
rect 30583 47894 31040 47927
rect 35294 47939 35332 47945
rect 35384 47939 35543 47945
rect 35595 47939 35754 47945
rect 35806 47939 35965 47945
rect 36017 47939 36176 47945
rect 36228 47939 36266 47945
rect 34870 47894 35025 47901
rect 35294 47899 36266 47939
rect 36438 47905 36953 47945
rect 37439 47937 37891 47945
rect 37943 47937 38071 47945
rect 38123 47937 38161 47945
rect 37439 47905 38161 47937
rect 37853 47897 38161 47905
rect 27387 47801 27790 47853
rect 27842 47801 28001 47853
rect 28053 47801 28212 47853
rect 28264 47801 28423 47853
rect 28475 47801 28634 47853
rect 28686 47850 28845 47853
rect 28686 47804 28810 47850
rect 28686 47801 28845 47804
rect 28897 47801 29056 47853
rect 29108 47801 29196 47853
rect 27387 47687 29196 47801
rect 29283 47853 30365 47894
rect 29283 47850 29582 47853
rect 29283 47804 29317 47850
rect 29363 47804 29478 47850
rect 29524 47804 29582 47850
rect 29283 47801 29582 47804
rect 29634 47850 29793 47853
rect 29845 47850 30005 47853
rect 29634 47804 29638 47850
rect 29684 47804 29793 47850
rect 29845 47804 29959 47850
rect 29634 47801 29793 47804
rect 29845 47801 30005 47804
rect 30057 47850 30216 47853
rect 30057 47804 30121 47850
rect 30167 47804 30216 47850
rect 30057 47801 30216 47804
rect 30268 47850 30365 47853
rect 30268 47804 30284 47850
rect 30330 47804 30365 47850
rect 30268 47801 30365 47804
rect 29283 47761 30365 47801
rect 30583 47853 32842 47894
rect 30583 47850 30854 47853
rect 30583 47804 30637 47850
rect 30683 47804 30854 47850
rect 30583 47801 30854 47804
rect 30906 47801 31065 47853
rect 31117 47801 31276 47853
rect 31328 47801 31486 47853
rect 31538 47801 31697 47853
rect 31749 47801 31909 47853
rect 31961 47801 32120 47853
rect 32172 47801 32330 47853
rect 32382 47801 32541 47853
rect 32593 47801 32752 47853
rect 32804 47801 32842 47853
rect 29544 47760 30306 47761
rect 30583 47760 32842 47801
rect 34717 47853 35025 47894
rect 38658 47885 39723 47945
rect 48905 47939 48943 47945
rect 48995 47939 49154 47945
rect 49206 47939 49365 47945
rect 49417 47939 49576 47945
rect 49628 47939 49787 47945
rect 49839 47939 49877 47945
rect 48905 47899 49877 47939
rect 54085 47927 54223 47973
rect 54269 47967 54440 47973
rect 54486 47967 54540 48013
rect 54269 47927 54540 47967
rect 50099 47894 50255 47901
rect 54085 47894 54540 47927
rect 55927 48620 56267 48666
rect 56313 48620 57736 48666
rect 55927 48544 57736 48620
rect 55927 48498 55961 48544
rect 56007 48503 57736 48544
rect 56007 48498 56267 48503
rect 55927 48457 56267 48498
rect 56313 48457 57736 48503
rect 55927 48381 57736 48457
rect 55927 48335 55961 48381
rect 56007 48340 57736 48381
rect 56007 48335 56267 48340
rect 55927 48294 56267 48335
rect 56313 48294 57736 48340
rect 55927 48217 57736 48294
rect 55927 48171 55961 48217
rect 56007 48177 57736 48217
rect 56007 48171 56267 48177
rect 55927 48131 56267 48171
rect 56313 48131 57736 48177
rect 55927 48054 57736 48131
rect 55927 48008 55961 48054
rect 56007 48013 57736 48054
rect 56007 48008 56267 48013
rect 55927 47967 56267 48008
rect 56313 47967 57736 48013
rect 34717 47801 34755 47853
rect 34807 47850 34935 47853
rect 34807 47804 34916 47850
rect 34807 47801 34935 47804
rect 34987 47801 35025 47853
rect 34717 47760 35025 47801
rect 50099 47853 50408 47894
rect 50099 47801 50138 47853
rect 50190 47850 50318 47853
rect 50206 47804 50318 47850
rect 50190 47801 50318 47804
rect 50370 47801 50408 47853
rect 27387 47641 28810 47687
rect 28856 47644 29196 47687
rect 28856 47641 29116 47644
rect 27387 47598 29116 47641
rect 29162 47598 29196 47644
rect 27387 47523 29196 47598
rect 27387 47477 28810 47523
rect 28856 47481 29196 47523
rect 28856 47477 29116 47481
rect 27387 47435 29116 47477
rect 29162 47435 29196 47481
rect 27387 47360 29196 47435
rect 27387 47314 28810 47360
rect 28856 47317 29196 47360
rect 28856 47314 29116 47317
rect 27387 47271 29116 47314
rect 29162 47271 29196 47317
rect 27387 47197 29196 47271
rect 27387 47151 28810 47197
rect 28856 47154 29196 47197
rect 28856 47151 29116 47154
rect 27387 47108 29116 47151
rect 29162 47108 29196 47154
rect 27387 47034 29196 47108
rect 27387 46988 28810 47034
rect 28856 46988 29196 47034
rect 30583 47727 31040 47760
rect 34870 47753 35025 47760
rect 30583 47687 30855 47727
rect 30583 47641 30637 47687
rect 30683 47681 30855 47687
rect 30901 47681 31040 47727
rect 35294 47715 36266 47755
rect 37853 47749 38161 47757
rect 35294 47709 35332 47715
rect 35384 47709 35543 47715
rect 35595 47709 35754 47715
rect 35806 47709 35965 47715
rect 36017 47709 36176 47715
rect 36228 47709 36266 47715
rect 36438 47709 36953 47749
rect 37439 47717 38161 47749
rect 37439 47709 37891 47717
rect 37943 47709 38071 47717
rect 38123 47709 38161 47717
rect 38658 47709 39723 47769
rect 50099 47760 50408 47801
rect 52278 47853 54540 47894
rect 52278 47801 52316 47853
rect 52368 47801 52527 47853
rect 52579 47801 52738 47853
rect 52790 47801 52948 47853
rect 53000 47801 53159 47853
rect 53211 47801 53371 47853
rect 53423 47801 53582 47853
rect 53634 47801 53792 47853
rect 53844 47801 54003 47853
rect 54055 47801 54214 47853
rect 54266 47850 54540 47853
rect 54266 47804 54440 47850
rect 54486 47804 54540 47850
rect 54266 47801 54540 47804
rect 52278 47760 54540 47801
rect 54758 47853 55840 47894
rect 54758 47850 54855 47853
rect 54758 47804 54793 47850
rect 54839 47804 54855 47850
rect 54758 47801 54855 47804
rect 54907 47850 55066 47853
rect 54907 47804 54956 47850
rect 55002 47804 55066 47850
rect 54907 47801 55066 47804
rect 55118 47850 55278 47853
rect 55330 47850 55489 47853
rect 55164 47804 55278 47850
rect 55330 47804 55439 47850
rect 55485 47804 55489 47850
rect 55118 47801 55278 47804
rect 55330 47801 55489 47804
rect 55541 47850 55840 47853
rect 55541 47804 55599 47850
rect 55645 47804 55760 47850
rect 55806 47804 55840 47850
rect 55541 47801 55840 47804
rect 54758 47761 55840 47801
rect 55927 47853 57736 47967
rect 55927 47801 56015 47853
rect 56067 47801 56226 47853
rect 56278 47850 56437 47853
rect 56313 47804 56437 47850
rect 56278 47801 56437 47804
rect 56489 47801 56648 47853
rect 56700 47801 56859 47853
rect 56911 47801 57070 47853
rect 57122 47801 57281 47853
rect 57333 47801 57736 47853
rect 54817 47760 55579 47761
rect 48905 47715 49877 47755
rect 50099 47753 50255 47760
rect 48905 47709 48943 47715
rect 48995 47709 49154 47715
rect 49206 47709 49365 47715
rect 49417 47709 49576 47715
rect 49628 47709 49787 47715
rect 49839 47709 49877 47715
rect 30683 47641 31040 47681
rect 33484 47665 34643 47694
rect 30583 47564 31040 47641
rect 33019 47625 33327 47665
rect 33019 47622 33057 47625
rect 33109 47622 33237 47625
rect 33289 47622 33327 47625
rect 33484 47657 35082 47665
rect 35260 47663 35273 47709
rect 35523 47663 35543 47709
rect 35626 47663 35683 47709
rect 35729 47663 35754 47709
rect 35832 47663 35889 47709
rect 35935 47663 35965 47709
rect 36038 47663 36095 47709
rect 36141 47663 36176 47709
rect 36244 47663 36301 47709
rect 36347 47663 36360 47709
rect 36438 47663 36854 47709
rect 36900 47663 36971 47709
rect 37017 47663 37088 47709
rect 37134 47663 37206 47709
rect 37252 47663 37324 47709
rect 37370 47663 37442 47709
rect 37488 47665 37891 47709
rect 37488 47663 37909 47665
rect 37955 47663 38026 47709
rect 38123 47665 38143 47709
rect 38072 47663 38143 47665
rect 38189 47663 38261 47709
rect 38307 47663 38379 47709
rect 38425 47663 38497 47709
rect 38543 47663 38556 47709
rect 38658 47663 39021 47709
rect 39067 47663 39144 47709
rect 39190 47663 39267 47709
rect 39313 47663 39641 47709
rect 39687 47663 39730 47709
rect 31336 47576 31349 47622
rect 33323 47576 33336 47622
rect 33484 47611 33816 47657
rect 33862 47611 34002 47657
rect 34048 47611 34189 47657
rect 34235 47611 34376 47657
rect 34422 47611 34562 47657
rect 34608 47611 35082 47657
rect 35294 47623 36266 47663
rect 36438 47629 36953 47663
rect 37439 47629 38161 47663
rect 30583 47523 30855 47564
rect 30583 47477 30637 47523
rect 30683 47518 30855 47523
rect 30901 47518 31040 47564
rect 33019 47573 33057 47576
rect 33109 47573 33237 47576
rect 33289 47573 33327 47576
rect 33019 47532 33327 47573
rect 33484 47574 35082 47611
rect 30683 47477 31040 47518
rect 30583 47449 31040 47477
rect 33484 47492 33552 47574
rect 30583 47401 31493 47449
rect 30583 47360 30855 47401
rect 30583 47314 30637 47360
rect 30683 47355 30855 47360
rect 30901 47398 31493 47401
rect 30901 47355 31349 47398
rect 30683 47352 31349 47355
rect 33323 47352 33336 47398
rect 30683 47330 31493 47352
rect 30683 47314 31040 47330
rect 30583 47238 31040 47314
rect 30583 47197 30855 47238
rect 30583 47151 30637 47197
rect 30683 47192 30855 47197
rect 30901 47192 31040 47238
rect 30683 47151 31040 47192
rect 33019 47177 33327 47217
rect 33019 47174 33057 47177
rect 33109 47174 33237 47177
rect 33289 47174 33327 47177
rect 30583 47074 31040 47151
rect 31336 47128 31349 47174
rect 33323 47128 33336 47174
rect 33019 47125 33057 47128
rect 33109 47125 33237 47128
rect 33289 47125 33327 47128
rect 33019 47084 33327 47125
rect 30583 47034 30855 47074
rect 27387 46866 29196 46988
rect 27387 46820 28810 46866
rect 28856 46820 29196 46866
rect 29283 46953 30365 46994
rect 29283 46950 29582 46953
rect 29283 46904 29317 46950
rect 29363 46904 29478 46950
rect 29524 46904 29582 46950
rect 29283 46901 29582 46904
rect 29634 46950 29793 46953
rect 29845 46950 30005 46953
rect 29634 46904 29638 46950
rect 29684 46904 29793 46950
rect 29845 46904 29959 46950
rect 29634 46901 29793 46904
rect 29845 46901 30005 46904
rect 30057 46950 30216 46953
rect 30057 46904 30121 46950
rect 30167 46904 30216 46950
rect 30057 46901 30216 46904
rect 30268 46950 30365 46953
rect 30268 46904 30284 46950
rect 30330 46904 30365 46950
rect 30268 46901 30365 46904
rect 29283 46861 30365 46901
rect 30583 46988 30637 47034
rect 30683 47028 30855 47034
rect 30901 47028 31040 47074
rect 33484 47070 33495 47492
rect 33541 47070 33552 47492
rect 34964 47517 35082 47574
rect 36438 47529 36554 47629
rect 37853 47624 38161 47629
rect 38658 47649 39723 47663
rect 34964 47485 36360 47517
rect 34228 47415 34718 47456
rect 34228 47398 34267 47415
rect 34319 47398 34447 47415
rect 34499 47398 34627 47415
rect 33671 47352 33684 47398
rect 33730 47352 33787 47398
rect 33833 47352 33890 47398
rect 33936 47352 33993 47398
rect 34039 47352 34096 47398
rect 34142 47352 34199 47398
rect 34245 47363 34267 47398
rect 34245 47352 34302 47363
rect 34348 47352 34405 47398
rect 34499 47363 34508 47398
rect 34451 47352 34508 47363
rect 34554 47352 34612 47398
rect 34679 47363 34718 47415
rect 34964 47439 35273 47485
rect 35523 47439 35580 47485
rect 35626 47439 35683 47485
rect 35729 47439 35786 47485
rect 35832 47439 35889 47485
rect 35935 47439 35992 47485
rect 36038 47439 36095 47485
rect 36141 47439 36198 47485
rect 36244 47439 36301 47485
rect 36347 47439 36360 47485
rect 34964 47395 36360 47439
rect 34658 47352 34718 47363
rect 34228 47323 34718 47352
rect 36438 47389 36475 47529
rect 36521 47389 36554 47529
rect 35294 47261 36266 47295
rect 36438 47286 36554 47389
rect 36640 47529 36773 47549
rect 36640 47490 36697 47529
rect 36640 47438 36678 47490
rect 36640 47389 36697 47438
rect 36743 47389 36773 47529
rect 38658 47527 38726 47649
rect 39809 47643 44918 47681
rect 48765 47663 48778 47709
rect 48824 47663 48881 47709
rect 48927 47663 48943 47709
rect 49030 47663 49087 47709
rect 49133 47663 49154 47709
rect 49236 47663 49293 47709
rect 49339 47663 49365 47709
rect 49442 47663 49499 47709
rect 49545 47663 49576 47709
rect 49852 47663 49877 47709
rect 54085 47727 54540 47760
rect 50481 47667 51657 47694
rect 39809 47597 43739 47643
rect 43785 47597 43906 47643
rect 43952 47597 44071 47643
rect 44117 47597 44236 47643
rect 44282 47622 44918 47643
rect 48905 47623 49877 47663
rect 50044 47657 51657 47667
rect 44282 47597 44812 47622
rect 39809 47594 44812 47597
rect 39809 47548 39844 47594
rect 39890 47592 44812 47594
rect 39890 47548 39994 47592
rect 39809 47540 39994 47548
rect 40046 47576 44812 47592
rect 44858 47576 44925 47622
rect 44971 47576 45038 47622
rect 45084 47576 45151 47622
rect 45197 47576 45264 47622
rect 45310 47576 45323 47622
rect 48557 47577 48687 47617
rect 40046 47561 44918 47576
rect 40046 47540 40085 47561
rect 39809 47537 40085 47540
rect 36924 47517 37685 47524
rect 36923 47485 37931 47517
rect 36841 47439 36854 47485
rect 36900 47483 36971 47485
rect 36900 47439 36961 47483
rect 37017 47439 37088 47485
rect 37134 47483 37206 47485
rect 37134 47439 37172 47483
rect 37252 47439 37324 47485
rect 37370 47483 37442 47485
rect 37370 47439 37384 47483
rect 36923 47431 36961 47439
rect 37013 47431 37172 47439
rect 37224 47431 37384 47439
rect 37436 47439 37442 47483
rect 37488 47483 37909 47485
rect 37488 47439 37595 47483
rect 37436 47431 37595 47439
rect 37647 47439 37909 47483
rect 37955 47439 38026 47485
rect 38072 47439 38143 47485
rect 38189 47439 38261 47485
rect 38307 47439 38379 47485
rect 38425 47439 38497 47485
rect 38543 47439 38556 47485
rect 37647 47431 37931 47439
rect 36923 47398 37931 47431
rect 36923 47397 37685 47398
rect 36924 47391 37685 47397
rect 36640 47366 36773 47389
rect 38658 47387 38669 47527
rect 38715 47387 38726 47527
rect 39014 47485 39323 47517
rect 39492 47485 39608 47517
rect 39008 47439 39021 47485
rect 39067 47439 39144 47485
rect 39190 47439 39267 47485
rect 39313 47439 39326 47485
rect 39492 47439 39641 47485
rect 39687 47439 39730 47485
rect 38658 47376 38726 47387
rect 36438 47261 36953 47286
rect 37439 47283 37931 47286
rect 37439 47261 38161 47283
rect 35260 47215 35273 47261
rect 35523 47255 35580 47261
rect 35523 47215 35543 47255
rect 35626 47215 35683 47261
rect 35729 47255 35786 47261
rect 35729 47215 35754 47255
rect 35832 47215 35889 47261
rect 35935 47255 35992 47261
rect 35935 47215 35965 47255
rect 36038 47215 36095 47261
rect 36141 47255 36198 47261
rect 36141 47215 36176 47255
rect 36244 47215 36301 47261
rect 36347 47215 36360 47261
rect 36438 47215 36854 47261
rect 36900 47215 36971 47261
rect 37017 47215 37088 47261
rect 37134 47215 37206 47261
rect 37252 47215 37324 47261
rect 37370 47215 37442 47261
rect 37488 47243 37909 47261
rect 37488 47215 37891 47243
rect 37955 47215 38026 47261
rect 38072 47243 38143 47261
rect 38123 47215 38143 47243
rect 38189 47215 38261 47261
rect 38307 47215 38379 47261
rect 38425 47215 38497 47261
rect 38543 47215 38556 47261
rect 33781 47174 34089 47209
rect 35294 47203 35332 47215
rect 35384 47203 35543 47215
rect 35595 47203 35754 47215
rect 35806 47203 35965 47215
rect 36017 47203 36176 47215
rect 36228 47203 36266 47215
rect 33671 47128 33684 47174
rect 33730 47128 33787 47174
rect 33833 47169 33890 47174
rect 33871 47128 33890 47169
rect 33936 47128 33993 47174
rect 34039 47169 34096 47174
rect 34051 47128 34096 47169
rect 34142 47128 34199 47174
rect 34245 47128 34302 47174
rect 34348 47128 34405 47174
rect 34451 47128 34508 47174
rect 34554 47128 34612 47174
rect 34658 47128 34671 47174
rect 35294 47163 36266 47203
rect 36438 47166 36953 47215
rect 37439 47191 37891 47215
rect 37943 47191 38071 47215
rect 38123 47191 38161 47215
rect 37439 47166 38161 47191
rect 37853 47150 38161 47166
rect 33781 47117 33819 47128
rect 33871 47117 33999 47128
rect 34051 47117 34089 47128
rect 33781 47076 34089 47117
rect 33484 47059 33552 47070
rect 30683 46994 31040 47028
rect 30683 46988 32842 46994
rect 30583 46953 32842 46988
rect 34247 46987 35008 46994
rect 30583 46901 30854 46953
rect 30906 46901 31065 46953
rect 31117 46901 31276 46953
rect 31328 46950 31486 46953
rect 31538 46950 31697 46953
rect 31749 46950 31909 46953
rect 31961 46950 32120 46953
rect 32172 46950 32330 46953
rect 32382 46950 32541 46953
rect 32593 46950 32752 46953
rect 32804 46950 32842 46953
rect 34246 46953 35008 46987
rect 34246 46950 34284 46953
rect 34336 46950 34495 46953
rect 34547 46950 34707 46953
rect 31328 46904 31349 46950
rect 33323 46904 33336 46950
rect 33671 46904 33684 46950
rect 33730 46904 33787 46950
rect 33833 46904 33890 46950
rect 33936 46904 33993 46950
rect 34039 46904 34096 46950
rect 34142 46904 34199 46950
rect 34245 46904 34284 46950
rect 34348 46904 34405 46950
rect 34451 46904 34495 46950
rect 34554 46904 34612 46950
rect 34658 46904 34707 46950
rect 31328 46901 31486 46904
rect 31538 46901 31697 46904
rect 31749 46901 31909 46904
rect 31961 46901 32120 46904
rect 32172 46901 32330 46904
rect 32382 46901 32541 46904
rect 32593 46901 32752 46904
rect 32804 46901 32842 46904
rect 30583 46866 32842 46901
rect 34246 46901 34284 46904
rect 34336 46901 34495 46904
rect 34547 46901 34707 46904
rect 34759 46901 34918 46953
rect 34970 46901 35008 46953
rect 34246 46867 35008 46901
rect 29544 46860 30306 46861
rect 27387 46744 29196 46820
rect 27387 46703 29116 46744
rect 27387 46657 28810 46703
rect 28856 46698 29116 46703
rect 29162 46698 29196 46744
rect 28856 46657 29196 46698
rect 27387 46581 29196 46657
rect 27387 46540 29116 46581
rect 27387 46494 28810 46540
rect 28856 46535 29116 46540
rect 29162 46535 29196 46581
rect 28856 46494 29196 46535
rect 27387 46417 29196 46494
rect 27387 46377 29116 46417
rect 27387 46331 28810 46377
rect 28856 46371 29116 46377
rect 29162 46371 29196 46417
rect 28856 46331 29196 46371
rect 27387 46254 29196 46331
rect 27387 46213 29116 46254
rect 27387 46167 28810 46213
rect 28856 46208 29116 46213
rect 29162 46208 29196 46254
rect 28856 46167 29196 46208
rect 27387 46053 29196 46167
rect 30583 46820 30637 46866
rect 30683 46860 32842 46866
rect 34247 46860 35008 46867
rect 35182 46987 36364 46994
rect 35182 46953 36958 46987
rect 35182 46901 35220 46953
rect 35272 46901 35430 46953
rect 35482 46901 35641 46953
rect 35693 46901 35853 46953
rect 35905 46901 36064 46953
rect 36116 46901 36274 46953
rect 36326 46950 36958 46953
rect 36326 46904 36489 46950
rect 36723 46904 36958 46950
rect 36326 46901 36958 46904
rect 35182 46867 36958 46901
rect 37946 46953 38842 46994
rect 37946 46950 38330 46953
rect 38382 46950 38541 46953
rect 37946 46904 37957 46950
rect 38473 46904 38541 46950
rect 37946 46901 38330 46904
rect 38382 46901 38541 46904
rect 38593 46901 38752 46953
rect 38804 46901 38842 46953
rect 35182 46860 36364 46867
rect 37946 46860 38842 46901
rect 39014 46953 39323 47439
rect 39014 46901 39052 46953
rect 39104 46950 39232 46953
rect 39108 46904 39220 46950
rect 39104 46901 39232 46904
rect 39284 46901 39323 46953
rect 30683 46826 31040 46860
rect 30683 46820 30855 46826
rect 30583 46780 30855 46820
rect 30901 46780 31040 46826
rect 30583 46703 31040 46780
rect 33484 46784 33552 46795
rect 33019 46729 33327 46770
rect 33019 46726 33057 46729
rect 33109 46726 33237 46729
rect 33289 46726 33327 46729
rect 30583 46657 30637 46703
rect 30683 46662 31040 46703
rect 31336 46680 31349 46726
rect 33323 46680 33336 46726
rect 30683 46657 30855 46662
rect 30583 46616 30855 46657
rect 30901 46616 31040 46662
rect 33019 46677 33057 46680
rect 33109 46677 33237 46680
rect 33289 46677 33327 46680
rect 33019 46637 33327 46677
rect 30583 46540 31040 46616
rect 30583 46494 30637 46540
rect 30683 46524 31040 46540
rect 30683 46502 31493 46524
rect 30683 46499 31349 46502
rect 30683 46494 30855 46499
rect 30583 46453 30855 46494
rect 30901 46456 31349 46499
rect 33323 46456 33336 46502
rect 30901 46453 31493 46456
rect 30583 46405 31493 46453
rect 30583 46377 31040 46405
rect 30583 46331 30637 46377
rect 30683 46336 31040 46377
rect 30683 46331 30855 46336
rect 30583 46290 30855 46331
rect 30901 46290 31040 46336
rect 33484 46362 33495 46784
rect 33541 46362 33552 46784
rect 33781 46737 34089 46778
rect 33781 46726 33819 46737
rect 33871 46726 33999 46737
rect 34051 46726 34089 46737
rect 33671 46680 33684 46726
rect 33730 46680 33787 46726
rect 33871 46685 33890 46726
rect 33833 46680 33890 46685
rect 33936 46680 33993 46726
rect 34051 46685 34096 46726
rect 34039 46680 34096 46685
rect 34142 46680 34199 46726
rect 34245 46680 34302 46726
rect 34348 46680 34405 46726
rect 34451 46680 34508 46726
rect 34554 46680 34612 46726
rect 34658 46680 34671 46726
rect 33781 46645 34089 46680
rect 35294 46651 36266 46691
rect 37853 46688 38161 46704
rect 35294 46639 35332 46651
rect 35384 46639 35543 46651
rect 35595 46639 35754 46651
rect 35806 46639 35965 46651
rect 36017 46639 36176 46651
rect 36228 46639 36266 46651
rect 36438 46639 36953 46688
rect 37439 46663 38161 46688
rect 37439 46639 37891 46663
rect 37943 46639 38071 46663
rect 38123 46639 38161 46663
rect 35260 46593 35273 46639
rect 35523 46599 35543 46639
rect 35523 46593 35580 46599
rect 35626 46593 35683 46639
rect 35729 46599 35754 46639
rect 35729 46593 35786 46599
rect 35832 46593 35889 46639
rect 35935 46599 35965 46639
rect 35935 46593 35992 46599
rect 36038 46593 36095 46639
rect 36141 46599 36176 46639
rect 36141 46593 36198 46599
rect 36244 46593 36301 46639
rect 36347 46593 36360 46639
rect 36438 46593 36854 46639
rect 36900 46593 36971 46639
rect 37017 46593 37088 46639
rect 37134 46593 37206 46639
rect 37252 46593 37324 46639
rect 37370 46593 37442 46639
rect 37488 46611 37891 46639
rect 37488 46593 37909 46611
rect 37955 46593 38026 46639
rect 38123 46611 38143 46639
rect 38072 46593 38143 46611
rect 38189 46593 38261 46639
rect 38307 46593 38379 46639
rect 38425 46593 38497 46639
rect 38543 46593 38556 46639
rect 35294 46559 36266 46593
rect 36438 46568 36953 46593
rect 37439 46571 38161 46593
rect 37439 46568 37931 46571
rect 34228 46502 34718 46531
rect 33671 46456 33684 46502
rect 33730 46456 33787 46502
rect 33833 46456 33890 46502
rect 33936 46456 33993 46502
rect 34039 46456 34096 46502
rect 34142 46456 34199 46502
rect 34245 46491 34302 46502
rect 34245 46456 34267 46491
rect 34348 46456 34405 46502
rect 34451 46491 34508 46502
rect 34499 46456 34508 46491
rect 34554 46456 34612 46502
rect 34658 46491 34718 46502
rect 34228 46439 34267 46456
rect 34319 46439 34447 46456
rect 34499 46439 34627 46456
rect 34679 46439 34718 46491
rect 36438 46465 36554 46568
rect 34228 46398 34718 46439
rect 34964 46415 36360 46459
rect 30583 46213 31040 46290
rect 33019 46281 33327 46322
rect 33019 46278 33057 46281
rect 33109 46278 33237 46281
rect 33289 46278 33327 46281
rect 33484 46280 33552 46362
rect 34964 46369 35273 46415
rect 35523 46369 35580 46415
rect 35626 46369 35683 46415
rect 35729 46369 35786 46415
rect 35832 46369 35889 46415
rect 35935 46369 35992 46415
rect 36038 46369 36095 46415
rect 36141 46369 36198 46415
rect 36244 46369 36301 46415
rect 36347 46369 36360 46415
rect 34964 46337 36360 46369
rect 34964 46280 35082 46337
rect 31336 46232 31349 46278
rect 33323 46232 33336 46278
rect 33484 46243 35082 46280
rect 30583 46167 30637 46213
rect 30683 46173 31040 46213
rect 33019 46229 33057 46232
rect 33109 46229 33237 46232
rect 33289 46229 33327 46232
rect 33019 46189 33327 46229
rect 33484 46197 33816 46243
rect 33862 46197 34002 46243
rect 34048 46197 34189 46243
rect 34235 46197 34376 46243
rect 34422 46197 34562 46243
rect 34608 46197 35082 46243
rect 36438 46325 36475 46465
rect 36521 46325 36554 46465
rect 33484 46189 35082 46197
rect 35294 46191 36266 46231
rect 36438 46225 36554 46325
rect 36640 46465 36773 46488
rect 36640 46416 36697 46465
rect 36640 46364 36678 46416
rect 36640 46325 36697 46364
rect 36743 46325 36773 46465
rect 38658 46467 38726 46478
rect 36924 46457 37685 46463
rect 36923 46456 37685 46457
rect 36923 46423 37931 46456
rect 36923 46415 36961 46423
rect 37013 46415 37172 46423
rect 37224 46415 37384 46423
rect 36841 46369 36854 46415
rect 36900 46371 36961 46415
rect 36900 46369 36971 46371
rect 37017 46369 37088 46415
rect 37134 46371 37172 46415
rect 37134 46369 37206 46371
rect 37252 46369 37324 46415
rect 37370 46371 37384 46415
rect 37436 46415 37595 46423
rect 37436 46371 37442 46415
rect 37370 46369 37442 46371
rect 37488 46371 37595 46415
rect 37647 46415 37931 46423
rect 37647 46371 37909 46415
rect 37488 46369 37909 46371
rect 37955 46369 38026 46415
rect 38072 46369 38143 46415
rect 38189 46369 38261 46415
rect 38307 46369 38379 46415
rect 38425 46369 38497 46415
rect 38543 46369 38556 46415
rect 36923 46337 37931 46369
rect 36924 46330 37685 46337
rect 36640 46305 36773 46325
rect 38658 46327 38669 46467
rect 38715 46327 38726 46467
rect 39014 46415 39323 46901
rect 39492 46987 39608 47439
rect 39923 47406 40085 47537
rect 39923 47354 39994 47406
rect 40046 47354 40085 47406
rect 39923 47314 40085 47354
rect 39737 47218 39865 47231
rect 39737 47191 39866 47218
rect 39737 47174 39775 47191
rect 39827 47174 39866 47191
rect 39727 47128 39740 47174
rect 39827 47139 39862 47174
rect 39786 47128 39862 47139
rect 39908 47128 39985 47174
rect 40031 47128 40108 47174
rect 40154 47128 40167 47174
rect 40246 47163 40362 47561
rect 42229 47422 44509 47463
rect 42229 47370 43068 47422
rect 43120 47370 44509 47422
rect 42229 47330 44509 47370
rect 44341 47286 44509 47330
rect 44341 47240 44358 47286
rect 44498 47240 44509 47286
rect 39737 47099 39866 47128
rect 40246 47117 40281 47163
rect 40327 47117 40362 47163
rect 40246 47080 40362 47117
rect 40718 47191 43524 47232
rect 44341 47229 44509 47240
rect 40718 47139 41935 47191
rect 41987 47139 43524 47191
rect 40718 47098 43524 47139
rect 44605 47174 44721 47561
rect 45400 47531 48379 47572
rect 45400 47517 46731 47531
rect 45400 47471 45464 47517
rect 45604 47479 46731 47517
rect 46783 47479 48379 47531
rect 45604 47471 48379 47479
rect 44901 47415 45241 47456
rect 45400 47438 48379 47471
rect 48557 47525 48596 47577
rect 48648 47525 48687 47577
rect 48557 47502 48687 47525
rect 50044 47611 50516 47657
rect 50562 47611 50703 47657
rect 50749 47611 50890 47657
rect 50936 47611 51076 47657
rect 51122 47611 51263 47657
rect 51309 47611 51657 47657
rect 51797 47647 52105 47687
rect 51797 47622 51835 47647
rect 51887 47622 52015 47647
rect 52067 47622 52105 47647
rect 54085 47681 54223 47727
rect 54269 47687 54540 47727
rect 54269 47681 54440 47687
rect 54085 47641 54440 47681
rect 54486 47641 54540 47687
rect 50044 47574 51657 47611
rect 51789 47576 51802 47622
rect 53776 47576 53789 47622
rect 50044 47517 50160 47574
rect 44901 47398 44939 47415
rect 44991 47398 45151 47415
rect 45203 47398 45241 47415
rect 44799 47352 44812 47398
rect 44858 47352 44925 47398
rect 44991 47363 45038 47398
rect 44971 47352 45038 47363
rect 45084 47352 45151 47398
rect 45203 47363 45264 47398
rect 45197 47352 45264 47363
rect 45310 47352 45323 47398
rect 48557 47362 48622 47502
rect 48668 47362 48687 47502
rect 49820 47485 50160 47517
rect 48765 47439 48778 47485
rect 48824 47439 48881 47485
rect 48927 47439 48984 47485
rect 49030 47439 49087 47485
rect 49133 47439 49190 47485
rect 49236 47439 49293 47485
rect 49339 47439 49396 47485
rect 49442 47439 49499 47485
rect 49545 47439 49602 47485
rect 49852 47439 50160 47485
rect 51589 47522 51657 47574
rect 51797 47554 52105 47576
rect 49820 47398 50160 47439
rect 50262 47415 50812 47456
rect 48557 47359 48687 47362
rect 44901 47323 45241 47352
rect 48557 47307 48596 47359
rect 48648 47307 48687 47359
rect 50262 47363 50300 47415
rect 50352 47398 50511 47415
rect 50563 47398 50722 47415
rect 50352 47363 50467 47398
rect 50563 47363 50571 47398
rect 50262 47352 50467 47363
rect 50513 47352 50571 47363
rect 50617 47352 50674 47398
rect 50720 47363 50722 47398
rect 50774 47398 50812 47415
rect 50774 47363 50777 47398
rect 50720 47352 50777 47363
rect 50823 47352 50880 47398
rect 50926 47352 50983 47398
rect 51029 47352 51086 47398
rect 51132 47352 51189 47398
rect 51235 47352 51292 47398
rect 51338 47352 51395 47398
rect 51441 47352 51454 47398
rect 50262 47323 50812 47352
rect 48557 47266 48687 47307
rect 48905 47261 49877 47292
rect 48765 47215 48778 47261
rect 48824 47215 48881 47261
rect 48927 47252 48984 47261
rect 48927 47215 48943 47252
rect 49030 47215 49087 47261
rect 49133 47252 49190 47261
rect 49133 47215 49154 47252
rect 49236 47215 49293 47261
rect 49339 47252 49396 47261
rect 49339 47215 49365 47252
rect 49442 47215 49499 47261
rect 49545 47252 49602 47261
rect 49545 47215 49576 47252
rect 49852 47215 49877 47261
rect 48905 47200 48943 47215
rect 48995 47200 49154 47215
rect 49206 47200 49365 47215
rect 49417 47200 49576 47215
rect 49628 47200 49787 47215
rect 49839 47200 49877 47215
rect 44605 47128 44812 47174
rect 44858 47128 44925 47174
rect 44971 47128 45038 47174
rect 45084 47128 45151 47174
rect 45197 47128 45264 47174
rect 45310 47128 45323 47174
rect 48905 47160 49877 47200
rect 51035 47177 51343 47217
rect 51035 47174 51073 47177
rect 51125 47174 51253 47177
rect 51305 47174 51343 47177
rect 43362 47091 43524 47098
rect 43362 47045 43373 47091
rect 43513 47045 43524 47091
rect 43362 47034 43524 47045
rect 45584 47114 48546 47150
rect 50454 47128 50467 47174
rect 50513 47128 50571 47174
rect 50617 47128 50674 47174
rect 50720 47128 50777 47174
rect 50823 47128 50880 47174
rect 50926 47128 50983 47174
rect 51029 47128 51073 47174
rect 51132 47128 51189 47174
rect 51235 47128 51253 47174
rect 51338 47128 51395 47174
rect 51441 47128 51454 47174
rect 45584 47068 45619 47114
rect 45665 47068 45777 47114
rect 45823 47068 45935 47114
rect 45981 47068 46093 47114
rect 46139 47068 46251 47114
rect 46297 47068 46409 47114
rect 46455 47068 46568 47114
rect 46614 47068 46726 47114
rect 46772 47068 46884 47114
rect 46930 47068 47042 47114
rect 47088 47068 47200 47114
rect 47246 47068 47358 47114
rect 47404 47068 47516 47114
rect 47562 47068 47675 47114
rect 47721 47068 47833 47114
rect 47879 47068 47991 47114
rect 48037 47068 48149 47114
rect 48195 47068 48307 47114
rect 48353 47068 48465 47114
rect 48511 47068 48546 47114
rect 51035 47125 51073 47128
rect 51125 47125 51253 47128
rect 51305 47125 51343 47128
rect 51035 47084 51343 47125
rect 51589 47100 51600 47522
rect 51646 47100 51657 47522
rect 54085 47523 54540 47641
rect 54085 47477 54440 47523
rect 54486 47477 54540 47523
rect 54085 47449 54540 47477
rect 53585 47398 54540 47449
rect 51789 47352 51802 47398
rect 53776 47360 54540 47398
rect 53776 47352 54440 47360
rect 53585 47330 54440 47352
rect 54085 47314 54440 47330
rect 54486 47314 54540 47360
rect 54085 47238 54540 47314
rect 51797 47184 52105 47224
rect 51797 47174 51835 47184
rect 51887 47174 52015 47184
rect 52067 47174 52105 47184
rect 54085 47192 54223 47238
rect 54269 47197 54540 47238
rect 54269 47192 54440 47197
rect 51789 47128 51802 47174
rect 53776 47128 53789 47174
rect 54085 47151 54440 47192
rect 54486 47151 54540 47197
rect 51589 47089 51657 47100
rect 51797 47091 52105 47128
rect 40215 46987 40523 46994
rect 40788 46987 42986 47001
rect 43753 46987 44514 46994
rect 39492 46964 42986 46987
rect 43704 46964 44514 46987
rect 39492 46953 44514 46964
rect 39492 46950 40253 46953
rect 39492 46904 39740 46950
rect 39786 46904 39862 46950
rect 39908 46904 39985 46950
rect 40031 46904 40108 46950
rect 40154 46904 40253 46950
rect 39492 46901 40253 46904
rect 40305 46901 40433 46953
rect 40485 46950 43790 46953
rect 40485 46904 40836 46950
rect 40882 46904 40994 46950
rect 41040 46904 41152 46950
rect 41198 46904 41310 46950
rect 41356 46904 41469 46950
rect 41515 46904 41627 46950
rect 41673 46904 41785 46950
rect 41831 46904 41943 46950
rect 41989 46904 42101 46950
rect 42147 46904 42259 46950
rect 42305 46904 42418 46950
rect 42464 46904 42576 46950
rect 42622 46904 42734 46950
rect 42780 46904 42892 46950
rect 42938 46904 43739 46950
rect 43785 46904 43790 46950
rect 40485 46901 43790 46904
rect 43842 46950 44001 46953
rect 43842 46904 43906 46950
rect 43952 46904 44001 46950
rect 43842 46901 44001 46904
rect 44053 46950 44213 46953
rect 44265 46950 44424 46953
rect 44053 46904 44071 46950
rect 44117 46904 44213 46950
rect 44282 46904 44424 46950
rect 44053 46901 44213 46904
rect 44265 46901 44424 46904
rect 44476 46901 44514 46953
rect 39492 46890 44514 46901
rect 39492 46867 42986 46890
rect 43704 46867 44514 46890
rect 39492 46415 39608 46867
rect 40215 46860 40523 46867
rect 40788 46853 42986 46867
rect 43753 46860 44514 46867
rect 44796 46987 45346 46994
rect 45584 46987 48546 47068
rect 54085 47074 54540 47151
rect 54085 47028 54223 47074
rect 54269 47034 54540 47074
rect 54269 47028 54440 47034
rect 54085 46994 54440 47028
rect 48800 46987 49982 46994
rect 50308 46987 50859 46994
rect 44796 46953 49982 46987
rect 44796 46950 44834 46953
rect 44886 46950 45045 46953
rect 45097 46950 45256 46953
rect 45308 46950 48838 46953
rect 44796 46904 44812 46950
rect 44886 46904 44925 46950
rect 44971 46904 45038 46950
rect 45097 46904 45151 46950
rect 45197 46904 45256 46950
rect 45310 46904 45619 46950
rect 45665 46904 45777 46950
rect 45823 46904 45935 46950
rect 45981 46904 46093 46950
rect 46139 46904 46251 46950
rect 46297 46904 46409 46950
rect 46455 46904 46568 46950
rect 46614 46904 46726 46950
rect 46772 46904 46884 46950
rect 46930 46904 47042 46950
rect 47088 46904 47200 46950
rect 47246 46904 47358 46950
rect 47404 46904 47516 46950
rect 47562 46904 47675 46950
rect 47721 46904 47833 46950
rect 47879 46904 47991 46950
rect 48037 46904 48149 46950
rect 48195 46904 48307 46950
rect 48353 46904 48465 46950
rect 48511 46904 48838 46950
rect 44796 46901 44834 46904
rect 44886 46901 45045 46904
rect 45097 46901 45256 46904
rect 45308 46901 48838 46904
rect 48890 46901 49048 46953
rect 49100 46901 49259 46953
rect 49311 46901 49471 46953
rect 49523 46901 49682 46953
rect 49734 46901 49892 46953
rect 49944 46901 49982 46953
rect 44796 46867 49982 46901
rect 50307 46953 50859 46987
rect 50307 46901 50346 46953
rect 50398 46950 50557 46953
rect 50609 46950 50768 46953
rect 50820 46950 50859 46953
rect 52278 46988 54440 46994
rect 54486 46988 54540 47034
rect 55927 47687 57736 47801
rect 55927 47644 56267 47687
rect 55927 47598 55961 47644
rect 56007 47641 56267 47644
rect 56313 47641 57736 47687
rect 56007 47598 57736 47641
rect 55927 47523 57736 47598
rect 55927 47481 56267 47523
rect 55927 47435 55961 47481
rect 56007 47477 56267 47481
rect 56313 47477 57736 47523
rect 56007 47435 57736 47477
rect 55927 47360 57736 47435
rect 55927 47317 56267 47360
rect 55927 47271 55961 47317
rect 56007 47314 56267 47317
rect 56313 47314 57736 47360
rect 56007 47271 57736 47314
rect 55927 47197 57736 47271
rect 55927 47154 56267 47197
rect 55927 47108 55961 47154
rect 56007 47151 56267 47154
rect 56313 47151 57736 47197
rect 56007 47108 57736 47151
rect 55927 47034 57736 47108
rect 52278 46953 54540 46988
rect 52278 46950 52316 46953
rect 52368 46950 52527 46953
rect 52579 46950 52738 46953
rect 52790 46950 52948 46953
rect 53000 46950 53159 46953
rect 53211 46950 53371 46953
rect 53423 46950 53582 46953
rect 53634 46950 53792 46953
rect 50398 46904 50467 46950
rect 50513 46904 50557 46950
rect 50617 46904 50674 46950
rect 50720 46904 50768 46950
rect 50823 46904 50880 46950
rect 50926 46904 50983 46950
rect 51029 46904 51086 46950
rect 51132 46904 51189 46950
rect 51235 46904 51292 46950
rect 51338 46904 51395 46950
rect 51441 46904 51454 46950
rect 51789 46904 51802 46950
rect 53776 46904 53792 46950
rect 50398 46901 50557 46904
rect 50609 46901 50768 46904
rect 50820 46901 50859 46904
rect 50307 46867 50859 46901
rect 44796 46860 45346 46867
rect 43362 46809 43524 46820
rect 39737 46726 39866 46755
rect 40246 46737 40362 46774
rect 43362 46763 43373 46809
rect 43513 46763 43524 46809
rect 43362 46756 43524 46763
rect 39727 46680 39740 46726
rect 39786 46715 39862 46726
rect 39827 46680 39862 46715
rect 39908 46680 39985 46726
rect 40031 46680 40108 46726
rect 40154 46680 40167 46726
rect 40246 46691 40281 46737
rect 40327 46691 40362 46737
rect 39737 46663 39775 46680
rect 39827 46663 39866 46680
rect 39737 46636 39866 46663
rect 39737 46623 39865 46636
rect 39923 46500 40085 46540
rect 39923 46448 39994 46500
rect 40046 46448 40085 46500
rect 39008 46369 39021 46415
rect 39067 46369 39144 46415
rect 39190 46369 39267 46415
rect 39313 46369 39326 46415
rect 39492 46369 39641 46415
rect 39687 46369 39730 46415
rect 39014 46337 39323 46369
rect 39492 46337 39608 46369
rect 37853 46225 38161 46230
rect 36438 46191 36953 46225
rect 37439 46191 38161 46225
rect 38658 46205 38726 46327
rect 39923 46317 40085 46448
rect 39809 46314 40085 46317
rect 39809 46306 39994 46314
rect 39809 46260 39844 46306
rect 39890 46262 39994 46306
rect 40046 46293 40085 46314
rect 40246 46293 40362 46691
rect 40718 46715 43524 46756
rect 45584 46786 48546 46867
rect 48800 46860 49982 46867
rect 50308 46860 50859 46867
rect 52278 46901 52316 46904
rect 52368 46901 52527 46904
rect 52579 46901 52738 46904
rect 52790 46901 52948 46904
rect 53000 46901 53159 46904
rect 53211 46901 53371 46904
rect 53423 46901 53582 46904
rect 53634 46901 53792 46904
rect 53844 46901 54003 46953
rect 54055 46901 54214 46953
rect 54266 46901 54540 46953
rect 52278 46866 54540 46901
rect 52278 46860 54440 46866
rect 45584 46740 45619 46786
rect 45665 46740 45777 46786
rect 45823 46740 45935 46786
rect 45981 46740 46093 46786
rect 46139 46740 46251 46786
rect 46297 46740 46409 46786
rect 46455 46740 46568 46786
rect 46614 46740 46726 46786
rect 46772 46740 46884 46786
rect 46930 46740 47042 46786
rect 47088 46740 47200 46786
rect 47246 46740 47358 46786
rect 47404 46740 47516 46786
rect 47562 46740 47675 46786
rect 47721 46740 47833 46786
rect 47879 46740 47991 46786
rect 48037 46740 48149 46786
rect 48195 46740 48307 46786
rect 48353 46740 48465 46786
rect 48511 46740 48546 46786
rect 54085 46826 54440 46860
rect 54085 46780 54223 46826
rect 54269 46820 54440 46826
rect 54486 46820 54540 46866
rect 54758 46953 55840 46994
rect 54758 46950 54855 46953
rect 54758 46904 54793 46950
rect 54839 46904 54855 46950
rect 54758 46901 54855 46904
rect 54907 46950 55066 46953
rect 54907 46904 54956 46950
rect 55002 46904 55066 46950
rect 54907 46901 55066 46904
rect 55118 46950 55278 46953
rect 55330 46950 55489 46953
rect 55164 46904 55278 46950
rect 55330 46904 55439 46950
rect 55485 46904 55489 46950
rect 55118 46901 55278 46904
rect 55330 46901 55489 46904
rect 55541 46950 55840 46953
rect 55541 46904 55599 46950
rect 55645 46904 55760 46950
rect 55806 46904 55840 46950
rect 55541 46901 55840 46904
rect 54758 46861 55840 46901
rect 55927 46988 56267 47034
rect 56313 46988 57736 47034
rect 55927 46866 57736 46988
rect 54817 46860 55579 46861
rect 54269 46780 54540 46820
rect 40718 46663 41935 46715
rect 41987 46663 43524 46715
rect 40718 46622 43524 46663
rect 44605 46680 44812 46726
rect 44858 46680 44925 46726
rect 44971 46680 45038 46726
rect 45084 46680 45151 46726
rect 45197 46680 45264 46726
rect 45310 46680 45323 46726
rect 45584 46704 48546 46740
rect 51035 46729 51343 46770
rect 51035 46726 51073 46729
rect 51125 46726 51253 46729
rect 51305 46726 51343 46729
rect 51589 46754 51657 46765
rect 44341 46614 44509 46625
rect 44341 46568 44358 46614
rect 44498 46568 44509 46614
rect 44341 46524 44509 46568
rect 42229 46484 44509 46524
rect 42229 46432 43068 46484
rect 43120 46432 44509 46484
rect 42229 46391 44509 46432
rect 44605 46293 44721 46680
rect 48905 46654 49877 46694
rect 50454 46680 50467 46726
rect 50513 46680 50571 46726
rect 50617 46680 50674 46726
rect 50720 46680 50777 46726
rect 50823 46680 50880 46726
rect 50926 46680 50983 46726
rect 51029 46680 51073 46726
rect 51132 46680 51189 46726
rect 51235 46680 51253 46726
rect 51338 46680 51395 46726
rect 51441 46680 51454 46726
rect 48905 46639 48943 46654
rect 48995 46639 49154 46654
rect 49206 46639 49365 46654
rect 49417 46639 49576 46654
rect 49628 46639 49787 46654
rect 49839 46639 49877 46654
rect 48765 46593 48778 46639
rect 48824 46593 48881 46639
rect 48927 46602 48943 46639
rect 48927 46593 48984 46602
rect 49030 46593 49087 46639
rect 49133 46602 49154 46639
rect 49133 46593 49190 46602
rect 49236 46593 49293 46639
rect 49339 46602 49365 46639
rect 49339 46593 49396 46602
rect 49442 46593 49499 46639
rect 49545 46602 49576 46639
rect 49545 46593 49602 46602
rect 49852 46593 49877 46639
rect 51035 46677 51073 46680
rect 51125 46677 51253 46680
rect 51305 46677 51343 46680
rect 51035 46637 51343 46677
rect 48557 46547 48687 46588
rect 48905 46562 49877 46593
rect 44901 46502 45241 46531
rect 44799 46456 44812 46502
rect 44858 46456 44925 46502
rect 44971 46491 45038 46502
rect 44991 46456 45038 46491
rect 45084 46456 45151 46502
rect 45197 46491 45264 46502
rect 45203 46456 45264 46491
rect 45310 46456 45323 46502
rect 48557 46495 48596 46547
rect 48648 46495 48687 46547
rect 48557 46492 48687 46495
rect 44901 46439 44939 46456
rect 44991 46439 45151 46456
rect 45203 46439 45241 46456
rect 44901 46398 45241 46439
rect 45400 46383 48379 46416
rect 45400 46337 45464 46383
rect 45604 46375 48379 46383
rect 45604 46337 47108 46375
rect 45400 46323 47108 46337
rect 47160 46323 48379 46375
rect 40046 46278 44918 46293
rect 45400 46282 48379 46323
rect 48557 46352 48622 46492
rect 48668 46352 48687 46492
rect 50262 46502 50812 46531
rect 50262 46491 50467 46502
rect 50513 46491 50571 46502
rect 49820 46415 50160 46456
rect 48765 46369 48778 46415
rect 48824 46369 48881 46415
rect 48927 46369 48984 46415
rect 49030 46369 49087 46415
rect 49133 46369 49190 46415
rect 49236 46369 49293 46415
rect 49339 46369 49396 46415
rect 49442 46369 49499 46415
rect 49545 46369 49602 46415
rect 49852 46369 50160 46415
rect 50262 46439 50300 46491
rect 50352 46456 50467 46491
rect 50563 46456 50571 46491
rect 50617 46456 50674 46502
rect 50720 46491 50777 46502
rect 50720 46456 50722 46491
rect 50352 46439 50511 46456
rect 50563 46439 50722 46456
rect 50774 46456 50777 46491
rect 50823 46456 50880 46502
rect 50926 46456 50983 46502
rect 51029 46456 51086 46502
rect 51132 46456 51189 46502
rect 51235 46456 51292 46502
rect 51338 46456 51395 46502
rect 51441 46456 51454 46502
rect 50774 46439 50812 46456
rect 50262 46398 50812 46439
rect 48557 46329 48687 46352
rect 49820 46337 50160 46369
rect 40046 46262 44812 46278
rect 39890 46260 44812 46262
rect 39809 46257 44812 46260
rect 39809 46211 43739 46257
rect 43785 46211 43906 46257
rect 43952 46211 44071 46257
rect 44117 46211 44236 46257
rect 44282 46232 44812 46257
rect 44858 46232 44925 46278
rect 44971 46232 45038 46278
rect 45084 46232 45151 46278
rect 45197 46232 45264 46278
rect 45310 46232 45323 46278
rect 48557 46277 48596 46329
rect 48648 46277 48687 46329
rect 48557 46237 48687 46277
rect 50044 46280 50160 46337
rect 51589 46332 51600 46754
rect 51646 46332 51657 46754
rect 51797 46726 52105 46763
rect 51789 46680 51802 46726
rect 53776 46680 53789 46726
rect 54085 46703 54540 46780
rect 51797 46670 51835 46680
rect 51887 46670 52015 46680
rect 52067 46670 52105 46680
rect 51797 46630 52105 46670
rect 54085 46662 54440 46703
rect 54085 46616 54223 46662
rect 54269 46657 54440 46662
rect 54486 46657 54540 46703
rect 54269 46616 54540 46657
rect 54085 46540 54540 46616
rect 54085 46524 54440 46540
rect 53585 46502 54440 46524
rect 51789 46456 51802 46502
rect 53776 46494 54440 46502
rect 54486 46494 54540 46540
rect 53776 46456 54540 46494
rect 53585 46405 54540 46456
rect 51589 46280 51657 46332
rect 54085 46377 54540 46405
rect 54085 46331 54440 46377
rect 54486 46331 54540 46377
rect 50044 46243 51657 46280
rect 51797 46278 52105 46300
rect 44282 46211 44918 46232
rect 38658 46191 39723 46205
rect 30683 46167 30855 46173
rect 30583 46127 30855 46167
rect 30901 46127 31040 46173
rect 33484 46160 34643 46189
rect 35260 46145 35273 46191
rect 35523 46145 35543 46191
rect 35626 46145 35683 46191
rect 35729 46145 35754 46191
rect 35832 46145 35889 46191
rect 35935 46145 35965 46191
rect 36038 46145 36095 46191
rect 36141 46145 36176 46191
rect 36244 46145 36301 46191
rect 36347 46145 36360 46191
rect 36438 46145 36854 46191
rect 36900 46145 36971 46191
rect 37017 46145 37088 46191
rect 37134 46145 37206 46191
rect 37252 46145 37324 46191
rect 37370 46145 37442 46191
rect 37488 46189 37909 46191
rect 37488 46145 37891 46189
rect 37955 46145 38026 46191
rect 38072 46189 38143 46191
rect 38123 46145 38143 46189
rect 38189 46145 38261 46191
rect 38307 46145 38379 46191
rect 38425 46145 38497 46191
rect 38543 46145 38556 46191
rect 38658 46145 39021 46191
rect 39067 46145 39144 46191
rect 39190 46145 39267 46191
rect 39313 46145 39641 46191
rect 39687 46145 39730 46191
rect 39809 46173 44918 46211
rect 48905 46191 49877 46231
rect 48765 46145 48778 46191
rect 48824 46145 48881 46191
rect 48927 46145 48943 46191
rect 49030 46145 49087 46191
rect 49133 46145 49154 46191
rect 49236 46145 49293 46191
rect 49339 46145 49365 46191
rect 49442 46145 49499 46191
rect 49545 46145 49576 46191
rect 49852 46145 49877 46191
rect 50044 46197 50516 46243
rect 50562 46197 50703 46243
rect 50749 46197 50890 46243
rect 50936 46197 51076 46243
rect 51122 46197 51263 46243
rect 51309 46197 51657 46243
rect 51789 46232 51802 46278
rect 53776 46232 53789 46278
rect 50044 46187 51657 46197
rect 50481 46160 51657 46187
rect 51797 46207 51835 46232
rect 51887 46207 52015 46232
rect 52067 46207 52105 46232
rect 51797 46167 52105 46207
rect 54085 46213 54540 46331
rect 54085 46173 54440 46213
rect 30583 46094 31040 46127
rect 35294 46139 35332 46145
rect 35384 46139 35543 46145
rect 35595 46139 35754 46145
rect 35806 46139 35965 46145
rect 36017 46139 36176 46145
rect 36228 46139 36266 46145
rect 34870 46094 35025 46101
rect 35294 46099 36266 46139
rect 36438 46105 36953 46145
rect 37439 46137 37891 46145
rect 37943 46137 38071 46145
rect 38123 46137 38161 46145
rect 37439 46105 38161 46137
rect 37853 46097 38161 46105
rect 27387 46001 27790 46053
rect 27842 46001 28001 46053
rect 28053 46001 28212 46053
rect 28264 46001 28423 46053
rect 28475 46001 28634 46053
rect 28686 46050 28845 46053
rect 28686 46004 28810 46050
rect 28686 46001 28845 46004
rect 28897 46001 29056 46053
rect 29108 46001 29196 46053
rect 27387 45887 29196 46001
rect 29283 46053 30365 46094
rect 29283 46050 29582 46053
rect 29283 46004 29317 46050
rect 29363 46004 29478 46050
rect 29524 46004 29582 46050
rect 29283 46001 29582 46004
rect 29634 46050 29793 46053
rect 29845 46050 30005 46053
rect 29634 46004 29638 46050
rect 29684 46004 29793 46050
rect 29845 46004 29959 46050
rect 29634 46001 29793 46004
rect 29845 46001 30005 46004
rect 30057 46050 30216 46053
rect 30057 46004 30121 46050
rect 30167 46004 30216 46050
rect 30057 46001 30216 46004
rect 30268 46050 30365 46053
rect 30268 46004 30284 46050
rect 30330 46004 30365 46050
rect 30268 46001 30365 46004
rect 29283 45961 30365 46001
rect 30583 46053 32842 46094
rect 30583 46050 30854 46053
rect 30583 46004 30637 46050
rect 30683 46004 30854 46050
rect 30583 46001 30854 46004
rect 30906 46001 31065 46053
rect 31117 46001 31276 46053
rect 31328 46001 31486 46053
rect 31538 46001 31697 46053
rect 31749 46001 31909 46053
rect 31961 46001 32120 46053
rect 32172 46001 32330 46053
rect 32382 46001 32541 46053
rect 32593 46001 32752 46053
rect 32804 46001 32842 46053
rect 29544 45960 30306 45961
rect 30583 45960 32842 46001
rect 34717 46053 35025 46094
rect 38658 46085 39723 46145
rect 48905 46139 48943 46145
rect 48995 46139 49154 46145
rect 49206 46139 49365 46145
rect 49417 46139 49576 46145
rect 49628 46139 49787 46145
rect 49839 46139 49877 46145
rect 48905 46099 49877 46139
rect 54085 46127 54223 46173
rect 54269 46167 54440 46173
rect 54486 46167 54540 46213
rect 54269 46127 54540 46167
rect 50099 46094 50255 46101
rect 54085 46094 54540 46127
rect 55927 46820 56267 46866
rect 56313 46820 57736 46866
rect 55927 46744 57736 46820
rect 55927 46698 55961 46744
rect 56007 46703 57736 46744
rect 56007 46698 56267 46703
rect 55927 46657 56267 46698
rect 56313 46657 57736 46703
rect 55927 46581 57736 46657
rect 55927 46535 55961 46581
rect 56007 46540 57736 46581
rect 56007 46535 56267 46540
rect 55927 46494 56267 46535
rect 56313 46494 57736 46540
rect 55927 46417 57736 46494
rect 55927 46371 55961 46417
rect 56007 46377 57736 46417
rect 56007 46371 56267 46377
rect 55927 46331 56267 46371
rect 56313 46331 57736 46377
rect 55927 46254 57736 46331
rect 55927 46208 55961 46254
rect 56007 46213 57736 46254
rect 56007 46208 56267 46213
rect 55927 46167 56267 46208
rect 56313 46167 57736 46213
rect 34717 46001 34755 46053
rect 34807 46050 34935 46053
rect 34807 46004 34916 46050
rect 34807 46001 34935 46004
rect 34987 46001 35025 46053
rect 34717 45960 35025 46001
rect 50099 46053 50408 46094
rect 50099 46001 50138 46053
rect 50190 46050 50318 46053
rect 50206 46004 50318 46050
rect 50190 46001 50318 46004
rect 50370 46001 50408 46053
rect 27387 45841 28810 45887
rect 28856 45844 29196 45887
rect 28856 45841 29116 45844
rect 27387 45798 29116 45841
rect 29162 45798 29196 45844
rect 27387 45723 29196 45798
rect 27387 45677 28810 45723
rect 28856 45681 29196 45723
rect 28856 45677 29116 45681
rect 27387 45635 29116 45677
rect 29162 45635 29196 45681
rect 27387 45560 29196 45635
rect 27387 45514 28810 45560
rect 28856 45517 29196 45560
rect 28856 45514 29116 45517
rect 27387 45471 29116 45514
rect 29162 45471 29196 45517
rect 27387 45397 29196 45471
rect 27387 45351 28810 45397
rect 28856 45354 29196 45397
rect 28856 45351 29116 45354
rect 27387 45308 29116 45351
rect 29162 45308 29196 45354
rect 27387 45234 29196 45308
rect 27387 45188 28810 45234
rect 28856 45188 29196 45234
rect 30583 45927 31040 45960
rect 34870 45953 35025 45960
rect 30583 45887 30855 45927
rect 30583 45841 30637 45887
rect 30683 45881 30855 45887
rect 30901 45881 31040 45927
rect 35294 45915 36266 45955
rect 37853 45949 38161 45957
rect 35294 45909 35332 45915
rect 35384 45909 35543 45915
rect 35595 45909 35754 45915
rect 35806 45909 35965 45915
rect 36017 45909 36176 45915
rect 36228 45909 36266 45915
rect 36438 45909 36953 45949
rect 37439 45917 38161 45949
rect 37439 45909 37891 45917
rect 37943 45909 38071 45917
rect 38123 45909 38161 45917
rect 38658 45909 39723 45969
rect 50099 45960 50408 46001
rect 52278 46053 54540 46094
rect 52278 46001 52316 46053
rect 52368 46001 52527 46053
rect 52579 46001 52738 46053
rect 52790 46001 52948 46053
rect 53000 46001 53159 46053
rect 53211 46001 53371 46053
rect 53423 46001 53582 46053
rect 53634 46001 53792 46053
rect 53844 46001 54003 46053
rect 54055 46001 54214 46053
rect 54266 46050 54540 46053
rect 54266 46004 54440 46050
rect 54486 46004 54540 46050
rect 54266 46001 54540 46004
rect 52278 45960 54540 46001
rect 54758 46053 55840 46094
rect 54758 46050 54855 46053
rect 54758 46004 54793 46050
rect 54839 46004 54855 46050
rect 54758 46001 54855 46004
rect 54907 46050 55066 46053
rect 54907 46004 54956 46050
rect 55002 46004 55066 46050
rect 54907 46001 55066 46004
rect 55118 46050 55278 46053
rect 55330 46050 55489 46053
rect 55164 46004 55278 46050
rect 55330 46004 55439 46050
rect 55485 46004 55489 46050
rect 55118 46001 55278 46004
rect 55330 46001 55489 46004
rect 55541 46050 55840 46053
rect 55541 46004 55599 46050
rect 55645 46004 55760 46050
rect 55806 46004 55840 46050
rect 55541 46001 55840 46004
rect 54758 45961 55840 46001
rect 55927 46053 57736 46167
rect 55927 46001 56015 46053
rect 56067 46001 56226 46053
rect 56278 46050 56437 46053
rect 56313 46004 56437 46050
rect 56278 46001 56437 46004
rect 56489 46001 56648 46053
rect 56700 46001 56859 46053
rect 56911 46001 57070 46053
rect 57122 46001 57281 46053
rect 57333 46001 57736 46053
rect 54817 45960 55579 45961
rect 48905 45915 49877 45955
rect 50099 45953 50255 45960
rect 48905 45909 48943 45915
rect 48995 45909 49154 45915
rect 49206 45909 49365 45915
rect 49417 45909 49576 45915
rect 49628 45909 49787 45915
rect 49839 45909 49877 45915
rect 30683 45841 31040 45881
rect 33484 45865 34643 45894
rect 30583 45764 31040 45841
rect 33019 45825 33327 45865
rect 33019 45822 33057 45825
rect 33109 45822 33237 45825
rect 33289 45822 33327 45825
rect 33484 45857 35082 45865
rect 35260 45863 35273 45909
rect 35523 45863 35543 45909
rect 35626 45863 35683 45909
rect 35729 45863 35754 45909
rect 35832 45863 35889 45909
rect 35935 45863 35965 45909
rect 36038 45863 36095 45909
rect 36141 45863 36176 45909
rect 36244 45863 36301 45909
rect 36347 45863 36360 45909
rect 36438 45863 36854 45909
rect 36900 45863 36971 45909
rect 37017 45863 37088 45909
rect 37134 45863 37206 45909
rect 37252 45863 37324 45909
rect 37370 45863 37442 45909
rect 37488 45865 37891 45909
rect 37488 45863 37909 45865
rect 37955 45863 38026 45909
rect 38123 45865 38143 45909
rect 38072 45863 38143 45865
rect 38189 45863 38261 45909
rect 38307 45863 38379 45909
rect 38425 45863 38497 45909
rect 38543 45863 38556 45909
rect 38658 45863 39021 45909
rect 39067 45863 39144 45909
rect 39190 45863 39267 45909
rect 39313 45863 39641 45909
rect 39687 45863 39730 45909
rect 31336 45776 31349 45822
rect 33323 45776 33336 45822
rect 33484 45811 33816 45857
rect 33862 45811 34002 45857
rect 34048 45811 34189 45857
rect 34235 45811 34376 45857
rect 34422 45811 34562 45857
rect 34608 45811 35082 45857
rect 35294 45823 36266 45863
rect 36438 45829 36953 45863
rect 37439 45829 38161 45863
rect 30583 45723 30855 45764
rect 30583 45677 30637 45723
rect 30683 45718 30855 45723
rect 30901 45718 31040 45764
rect 33019 45773 33057 45776
rect 33109 45773 33237 45776
rect 33289 45773 33327 45776
rect 33019 45732 33327 45773
rect 33484 45774 35082 45811
rect 30683 45677 31040 45718
rect 30583 45649 31040 45677
rect 33484 45692 33552 45774
rect 30583 45601 31493 45649
rect 30583 45560 30855 45601
rect 30583 45514 30637 45560
rect 30683 45555 30855 45560
rect 30901 45598 31493 45601
rect 30901 45555 31349 45598
rect 30683 45552 31349 45555
rect 33323 45552 33336 45598
rect 30683 45530 31493 45552
rect 30683 45514 31040 45530
rect 30583 45438 31040 45514
rect 30583 45397 30855 45438
rect 30583 45351 30637 45397
rect 30683 45392 30855 45397
rect 30901 45392 31040 45438
rect 30683 45351 31040 45392
rect 33019 45377 33327 45417
rect 33019 45374 33057 45377
rect 33109 45374 33237 45377
rect 33289 45374 33327 45377
rect 30583 45274 31040 45351
rect 31336 45328 31349 45374
rect 33323 45328 33336 45374
rect 33019 45325 33057 45328
rect 33109 45325 33237 45328
rect 33289 45325 33327 45328
rect 33019 45284 33327 45325
rect 30583 45234 30855 45274
rect 27387 45066 29196 45188
rect 27387 45020 28810 45066
rect 28856 45020 29196 45066
rect 29283 45153 30365 45194
rect 29283 45150 29582 45153
rect 29283 45104 29317 45150
rect 29363 45104 29478 45150
rect 29524 45104 29582 45150
rect 29283 45101 29582 45104
rect 29634 45150 29793 45153
rect 29845 45150 30005 45153
rect 29634 45104 29638 45150
rect 29684 45104 29793 45150
rect 29845 45104 29959 45150
rect 29634 45101 29793 45104
rect 29845 45101 30005 45104
rect 30057 45150 30216 45153
rect 30057 45104 30121 45150
rect 30167 45104 30216 45150
rect 30057 45101 30216 45104
rect 30268 45150 30365 45153
rect 30268 45104 30284 45150
rect 30330 45104 30365 45150
rect 30268 45101 30365 45104
rect 29283 45061 30365 45101
rect 30583 45188 30637 45234
rect 30683 45228 30855 45234
rect 30901 45228 31040 45274
rect 33484 45270 33495 45692
rect 33541 45270 33552 45692
rect 34964 45717 35082 45774
rect 36438 45729 36554 45829
rect 37853 45824 38161 45829
rect 38658 45849 39723 45863
rect 34964 45685 36360 45717
rect 34228 45615 34718 45656
rect 34228 45598 34267 45615
rect 34319 45598 34447 45615
rect 34499 45598 34627 45615
rect 33671 45552 33684 45598
rect 33730 45552 33787 45598
rect 33833 45552 33890 45598
rect 33936 45552 33993 45598
rect 34039 45552 34096 45598
rect 34142 45552 34199 45598
rect 34245 45563 34267 45598
rect 34245 45552 34302 45563
rect 34348 45552 34405 45598
rect 34499 45563 34508 45598
rect 34451 45552 34508 45563
rect 34554 45552 34612 45598
rect 34679 45563 34718 45615
rect 34964 45639 35273 45685
rect 35523 45639 35580 45685
rect 35626 45639 35683 45685
rect 35729 45639 35786 45685
rect 35832 45639 35889 45685
rect 35935 45639 35992 45685
rect 36038 45639 36095 45685
rect 36141 45639 36198 45685
rect 36244 45639 36301 45685
rect 36347 45639 36360 45685
rect 34964 45595 36360 45639
rect 34658 45552 34718 45563
rect 34228 45523 34718 45552
rect 36438 45589 36475 45729
rect 36521 45589 36554 45729
rect 35294 45461 36266 45495
rect 36438 45486 36554 45589
rect 36640 45729 36773 45749
rect 36640 45690 36697 45729
rect 36640 45638 36678 45690
rect 36640 45589 36697 45638
rect 36743 45589 36773 45729
rect 38658 45727 38726 45849
rect 39809 45843 44918 45881
rect 48765 45863 48778 45909
rect 48824 45863 48881 45909
rect 48927 45863 48943 45909
rect 49030 45863 49087 45909
rect 49133 45863 49154 45909
rect 49236 45863 49293 45909
rect 49339 45863 49365 45909
rect 49442 45863 49499 45909
rect 49545 45863 49576 45909
rect 49852 45863 49877 45909
rect 54085 45927 54540 45960
rect 50481 45867 51657 45894
rect 39809 45797 43739 45843
rect 43785 45797 43906 45843
rect 43952 45797 44071 45843
rect 44117 45797 44236 45843
rect 44282 45822 44918 45843
rect 48905 45823 49877 45863
rect 50044 45857 51657 45867
rect 44282 45797 44812 45822
rect 39809 45794 44812 45797
rect 39809 45748 39844 45794
rect 39890 45792 44812 45794
rect 39890 45748 39994 45792
rect 39809 45740 39994 45748
rect 40046 45776 44812 45792
rect 44858 45776 44925 45822
rect 44971 45776 45038 45822
rect 45084 45776 45151 45822
rect 45197 45776 45264 45822
rect 45310 45776 45323 45822
rect 48557 45777 48687 45817
rect 40046 45761 44918 45776
rect 40046 45740 40085 45761
rect 39809 45737 40085 45740
rect 36924 45717 37685 45724
rect 36923 45685 37931 45717
rect 36841 45639 36854 45685
rect 36900 45683 36971 45685
rect 36900 45639 36961 45683
rect 37017 45639 37088 45685
rect 37134 45683 37206 45685
rect 37134 45639 37172 45683
rect 37252 45639 37324 45685
rect 37370 45683 37442 45685
rect 37370 45639 37384 45683
rect 36923 45631 36961 45639
rect 37013 45631 37172 45639
rect 37224 45631 37384 45639
rect 37436 45639 37442 45683
rect 37488 45683 37909 45685
rect 37488 45639 37595 45683
rect 37436 45631 37595 45639
rect 37647 45639 37909 45683
rect 37955 45639 38026 45685
rect 38072 45639 38143 45685
rect 38189 45639 38261 45685
rect 38307 45639 38379 45685
rect 38425 45639 38497 45685
rect 38543 45639 38556 45685
rect 37647 45631 37931 45639
rect 36923 45598 37931 45631
rect 36923 45597 37685 45598
rect 36924 45591 37685 45597
rect 36640 45566 36773 45589
rect 38658 45587 38669 45727
rect 38715 45587 38726 45727
rect 39014 45685 39323 45717
rect 39492 45685 39608 45717
rect 39008 45639 39021 45685
rect 39067 45639 39144 45685
rect 39190 45639 39267 45685
rect 39313 45639 39326 45685
rect 39492 45639 39641 45685
rect 39687 45639 39730 45685
rect 38658 45576 38726 45587
rect 36438 45461 36953 45486
rect 37439 45483 37931 45486
rect 37439 45461 38161 45483
rect 35260 45415 35273 45461
rect 35523 45455 35580 45461
rect 35523 45415 35543 45455
rect 35626 45415 35683 45461
rect 35729 45455 35786 45461
rect 35729 45415 35754 45455
rect 35832 45415 35889 45461
rect 35935 45455 35992 45461
rect 35935 45415 35965 45455
rect 36038 45415 36095 45461
rect 36141 45455 36198 45461
rect 36141 45415 36176 45455
rect 36244 45415 36301 45461
rect 36347 45415 36360 45461
rect 36438 45415 36854 45461
rect 36900 45415 36971 45461
rect 37017 45415 37088 45461
rect 37134 45415 37206 45461
rect 37252 45415 37324 45461
rect 37370 45415 37442 45461
rect 37488 45443 37909 45461
rect 37488 45415 37891 45443
rect 37955 45415 38026 45461
rect 38072 45443 38143 45461
rect 38123 45415 38143 45443
rect 38189 45415 38261 45461
rect 38307 45415 38379 45461
rect 38425 45415 38497 45461
rect 38543 45415 38556 45461
rect 33781 45374 34089 45409
rect 35294 45403 35332 45415
rect 35384 45403 35543 45415
rect 35595 45403 35754 45415
rect 35806 45403 35965 45415
rect 36017 45403 36176 45415
rect 36228 45403 36266 45415
rect 33671 45328 33684 45374
rect 33730 45328 33787 45374
rect 33833 45369 33890 45374
rect 33871 45328 33890 45369
rect 33936 45328 33993 45374
rect 34039 45369 34096 45374
rect 34051 45328 34096 45369
rect 34142 45328 34199 45374
rect 34245 45328 34302 45374
rect 34348 45328 34405 45374
rect 34451 45328 34508 45374
rect 34554 45328 34612 45374
rect 34658 45328 34671 45374
rect 35294 45363 36266 45403
rect 36438 45366 36953 45415
rect 37439 45391 37891 45415
rect 37943 45391 38071 45415
rect 38123 45391 38161 45415
rect 37439 45366 38161 45391
rect 37853 45350 38161 45366
rect 33781 45317 33819 45328
rect 33871 45317 33999 45328
rect 34051 45317 34089 45328
rect 33781 45276 34089 45317
rect 33484 45259 33552 45270
rect 30683 45194 31040 45228
rect 30683 45188 32842 45194
rect 30583 45153 32842 45188
rect 34247 45187 35008 45194
rect 30583 45101 30854 45153
rect 30906 45101 31065 45153
rect 31117 45101 31276 45153
rect 31328 45150 31486 45153
rect 31538 45150 31697 45153
rect 31749 45150 31909 45153
rect 31961 45150 32120 45153
rect 32172 45150 32330 45153
rect 32382 45150 32541 45153
rect 32593 45150 32752 45153
rect 32804 45150 32842 45153
rect 34246 45153 35008 45187
rect 34246 45150 34284 45153
rect 34336 45150 34495 45153
rect 34547 45150 34707 45153
rect 31328 45104 31349 45150
rect 33323 45104 33336 45150
rect 33671 45104 33684 45150
rect 33730 45104 33787 45150
rect 33833 45104 33890 45150
rect 33936 45104 33993 45150
rect 34039 45104 34096 45150
rect 34142 45104 34199 45150
rect 34245 45104 34284 45150
rect 34348 45104 34405 45150
rect 34451 45104 34495 45150
rect 34554 45104 34612 45150
rect 34658 45104 34707 45150
rect 31328 45101 31486 45104
rect 31538 45101 31697 45104
rect 31749 45101 31909 45104
rect 31961 45101 32120 45104
rect 32172 45101 32330 45104
rect 32382 45101 32541 45104
rect 32593 45101 32752 45104
rect 32804 45101 32842 45104
rect 30583 45066 32842 45101
rect 34246 45101 34284 45104
rect 34336 45101 34495 45104
rect 34547 45101 34707 45104
rect 34759 45101 34918 45153
rect 34970 45101 35008 45153
rect 34246 45067 35008 45101
rect 29544 45060 30306 45061
rect 27387 44944 29196 45020
rect 27387 44903 29116 44944
rect 27387 44857 28810 44903
rect 28856 44898 29116 44903
rect 29162 44898 29196 44944
rect 28856 44857 29196 44898
rect 27387 44781 29196 44857
rect 27387 44740 29116 44781
rect 27387 44694 28810 44740
rect 28856 44735 29116 44740
rect 29162 44735 29196 44781
rect 28856 44694 29196 44735
rect 27387 44617 29196 44694
rect 27387 44577 29116 44617
rect 27387 44531 28810 44577
rect 28856 44571 29116 44577
rect 29162 44571 29196 44617
rect 28856 44531 29196 44571
rect 27387 44454 29196 44531
rect 27387 44413 29116 44454
rect 27387 44367 28810 44413
rect 28856 44408 29116 44413
rect 29162 44408 29196 44454
rect 28856 44367 29196 44408
rect 27387 44253 29196 44367
rect 30583 45020 30637 45066
rect 30683 45060 32842 45066
rect 34247 45060 35008 45067
rect 35182 45187 36364 45194
rect 35182 45153 36958 45187
rect 35182 45101 35220 45153
rect 35272 45101 35430 45153
rect 35482 45101 35641 45153
rect 35693 45101 35853 45153
rect 35905 45101 36064 45153
rect 36116 45101 36274 45153
rect 36326 45150 36958 45153
rect 36326 45104 36489 45150
rect 36723 45104 36958 45150
rect 36326 45101 36958 45104
rect 35182 45067 36958 45101
rect 37946 45153 38842 45194
rect 37946 45150 38330 45153
rect 38382 45150 38541 45153
rect 37946 45104 37957 45150
rect 38473 45104 38541 45150
rect 37946 45101 38330 45104
rect 38382 45101 38541 45104
rect 38593 45101 38752 45153
rect 38804 45101 38842 45153
rect 35182 45060 36364 45067
rect 37946 45060 38842 45101
rect 39014 45153 39323 45639
rect 39014 45101 39052 45153
rect 39104 45150 39232 45153
rect 39108 45104 39220 45150
rect 39104 45101 39232 45104
rect 39284 45101 39323 45153
rect 30683 45026 31040 45060
rect 30683 45020 30855 45026
rect 30583 44980 30855 45020
rect 30901 44980 31040 45026
rect 30583 44903 31040 44980
rect 33484 44984 33552 44995
rect 33019 44929 33327 44970
rect 33019 44926 33057 44929
rect 33109 44926 33237 44929
rect 33289 44926 33327 44929
rect 30583 44857 30637 44903
rect 30683 44862 31040 44903
rect 31336 44880 31349 44926
rect 33323 44880 33336 44926
rect 30683 44857 30855 44862
rect 30583 44816 30855 44857
rect 30901 44816 31040 44862
rect 33019 44877 33057 44880
rect 33109 44877 33237 44880
rect 33289 44877 33327 44880
rect 33019 44837 33327 44877
rect 30583 44740 31040 44816
rect 30583 44694 30637 44740
rect 30683 44724 31040 44740
rect 30683 44702 31493 44724
rect 30683 44699 31349 44702
rect 30683 44694 30855 44699
rect 30583 44653 30855 44694
rect 30901 44656 31349 44699
rect 33323 44656 33336 44702
rect 30901 44653 31493 44656
rect 30583 44605 31493 44653
rect 30583 44577 31040 44605
rect 30583 44531 30637 44577
rect 30683 44536 31040 44577
rect 30683 44531 30855 44536
rect 30583 44490 30855 44531
rect 30901 44490 31040 44536
rect 33484 44562 33495 44984
rect 33541 44562 33552 44984
rect 33781 44937 34089 44978
rect 33781 44926 33819 44937
rect 33871 44926 33999 44937
rect 34051 44926 34089 44937
rect 33671 44880 33684 44926
rect 33730 44880 33787 44926
rect 33871 44885 33890 44926
rect 33833 44880 33890 44885
rect 33936 44880 33993 44926
rect 34051 44885 34096 44926
rect 34039 44880 34096 44885
rect 34142 44880 34199 44926
rect 34245 44880 34302 44926
rect 34348 44880 34405 44926
rect 34451 44880 34508 44926
rect 34554 44880 34612 44926
rect 34658 44880 34671 44926
rect 33781 44845 34089 44880
rect 35294 44851 36266 44891
rect 37853 44888 38161 44904
rect 35294 44839 35332 44851
rect 35384 44839 35543 44851
rect 35595 44839 35754 44851
rect 35806 44839 35965 44851
rect 36017 44839 36176 44851
rect 36228 44839 36266 44851
rect 36438 44839 36953 44888
rect 37439 44863 38161 44888
rect 37439 44839 37891 44863
rect 37943 44839 38071 44863
rect 38123 44839 38161 44863
rect 35260 44793 35273 44839
rect 35523 44799 35543 44839
rect 35523 44793 35580 44799
rect 35626 44793 35683 44839
rect 35729 44799 35754 44839
rect 35729 44793 35786 44799
rect 35832 44793 35889 44839
rect 35935 44799 35965 44839
rect 35935 44793 35992 44799
rect 36038 44793 36095 44839
rect 36141 44799 36176 44839
rect 36141 44793 36198 44799
rect 36244 44793 36301 44839
rect 36347 44793 36360 44839
rect 36438 44793 36854 44839
rect 36900 44793 36971 44839
rect 37017 44793 37088 44839
rect 37134 44793 37206 44839
rect 37252 44793 37324 44839
rect 37370 44793 37442 44839
rect 37488 44811 37891 44839
rect 37488 44793 37909 44811
rect 37955 44793 38026 44839
rect 38123 44811 38143 44839
rect 38072 44793 38143 44811
rect 38189 44793 38261 44839
rect 38307 44793 38379 44839
rect 38425 44793 38497 44839
rect 38543 44793 38556 44839
rect 35294 44759 36266 44793
rect 36438 44768 36953 44793
rect 37439 44771 38161 44793
rect 37439 44768 37931 44771
rect 34228 44702 34718 44731
rect 33671 44656 33684 44702
rect 33730 44656 33787 44702
rect 33833 44656 33890 44702
rect 33936 44656 33993 44702
rect 34039 44656 34096 44702
rect 34142 44656 34199 44702
rect 34245 44691 34302 44702
rect 34245 44656 34267 44691
rect 34348 44656 34405 44702
rect 34451 44691 34508 44702
rect 34499 44656 34508 44691
rect 34554 44656 34612 44702
rect 34658 44691 34718 44702
rect 34228 44639 34267 44656
rect 34319 44639 34447 44656
rect 34499 44639 34627 44656
rect 34679 44639 34718 44691
rect 36438 44665 36554 44768
rect 34228 44598 34718 44639
rect 34964 44615 36360 44659
rect 30583 44413 31040 44490
rect 33019 44481 33327 44522
rect 33019 44478 33057 44481
rect 33109 44478 33237 44481
rect 33289 44478 33327 44481
rect 33484 44480 33552 44562
rect 34964 44569 35273 44615
rect 35523 44569 35580 44615
rect 35626 44569 35683 44615
rect 35729 44569 35786 44615
rect 35832 44569 35889 44615
rect 35935 44569 35992 44615
rect 36038 44569 36095 44615
rect 36141 44569 36198 44615
rect 36244 44569 36301 44615
rect 36347 44569 36360 44615
rect 34964 44537 36360 44569
rect 34964 44480 35082 44537
rect 31336 44432 31349 44478
rect 33323 44432 33336 44478
rect 33484 44443 35082 44480
rect 30583 44367 30637 44413
rect 30683 44373 31040 44413
rect 33019 44429 33057 44432
rect 33109 44429 33237 44432
rect 33289 44429 33327 44432
rect 33019 44389 33327 44429
rect 33484 44397 33816 44443
rect 33862 44397 34002 44443
rect 34048 44397 34189 44443
rect 34235 44397 34376 44443
rect 34422 44397 34562 44443
rect 34608 44397 35082 44443
rect 36438 44525 36475 44665
rect 36521 44525 36554 44665
rect 33484 44389 35082 44397
rect 35294 44391 36266 44431
rect 36438 44425 36554 44525
rect 36640 44665 36773 44688
rect 36640 44616 36697 44665
rect 36640 44564 36678 44616
rect 36640 44525 36697 44564
rect 36743 44525 36773 44665
rect 38658 44667 38726 44678
rect 36924 44657 37685 44663
rect 36923 44656 37685 44657
rect 36923 44623 37931 44656
rect 36923 44615 36961 44623
rect 37013 44615 37172 44623
rect 37224 44615 37384 44623
rect 36841 44569 36854 44615
rect 36900 44571 36961 44615
rect 36900 44569 36971 44571
rect 37017 44569 37088 44615
rect 37134 44571 37172 44615
rect 37134 44569 37206 44571
rect 37252 44569 37324 44615
rect 37370 44571 37384 44615
rect 37436 44615 37595 44623
rect 37436 44571 37442 44615
rect 37370 44569 37442 44571
rect 37488 44571 37595 44615
rect 37647 44615 37931 44623
rect 37647 44571 37909 44615
rect 37488 44569 37909 44571
rect 37955 44569 38026 44615
rect 38072 44569 38143 44615
rect 38189 44569 38261 44615
rect 38307 44569 38379 44615
rect 38425 44569 38497 44615
rect 38543 44569 38556 44615
rect 36923 44537 37931 44569
rect 36924 44530 37685 44537
rect 36640 44505 36773 44525
rect 38658 44527 38669 44667
rect 38715 44527 38726 44667
rect 39014 44615 39323 45101
rect 39492 45187 39608 45639
rect 39923 45606 40085 45737
rect 39923 45554 39994 45606
rect 40046 45554 40085 45606
rect 39923 45514 40085 45554
rect 39737 45418 39865 45431
rect 39737 45391 39866 45418
rect 39737 45374 39775 45391
rect 39827 45374 39866 45391
rect 39727 45328 39740 45374
rect 39827 45339 39862 45374
rect 39786 45328 39862 45339
rect 39908 45328 39985 45374
rect 40031 45328 40108 45374
rect 40154 45328 40167 45374
rect 40246 45363 40362 45761
rect 42229 45622 44509 45663
rect 42229 45570 43068 45622
rect 43120 45570 44509 45622
rect 42229 45530 44509 45570
rect 44341 45486 44509 45530
rect 44341 45440 44358 45486
rect 44498 45440 44509 45486
rect 39737 45299 39866 45328
rect 40246 45317 40281 45363
rect 40327 45317 40362 45363
rect 40246 45280 40362 45317
rect 40718 45391 43524 45432
rect 44341 45429 44509 45440
rect 40718 45339 41935 45391
rect 41987 45339 43524 45391
rect 40718 45298 43524 45339
rect 44605 45374 44721 45761
rect 45400 45731 48379 45772
rect 45400 45717 47486 45731
rect 45400 45671 45464 45717
rect 45604 45679 47486 45717
rect 47538 45679 48379 45731
rect 45604 45671 48379 45679
rect 44901 45615 45241 45656
rect 45400 45638 48379 45671
rect 48557 45725 48596 45777
rect 48648 45725 48687 45777
rect 48557 45702 48687 45725
rect 50044 45811 50516 45857
rect 50562 45811 50703 45857
rect 50749 45811 50890 45857
rect 50936 45811 51076 45857
rect 51122 45811 51263 45857
rect 51309 45811 51657 45857
rect 51797 45847 52105 45887
rect 51797 45822 51835 45847
rect 51887 45822 52015 45847
rect 52067 45822 52105 45847
rect 54085 45881 54223 45927
rect 54269 45887 54540 45927
rect 54269 45881 54440 45887
rect 54085 45841 54440 45881
rect 54486 45841 54540 45887
rect 50044 45774 51657 45811
rect 51789 45776 51802 45822
rect 53776 45776 53789 45822
rect 50044 45717 50160 45774
rect 44901 45598 44939 45615
rect 44991 45598 45151 45615
rect 45203 45598 45241 45615
rect 44799 45552 44812 45598
rect 44858 45552 44925 45598
rect 44991 45563 45038 45598
rect 44971 45552 45038 45563
rect 45084 45552 45151 45598
rect 45203 45563 45264 45598
rect 45197 45552 45264 45563
rect 45310 45552 45323 45598
rect 48557 45562 48622 45702
rect 48668 45562 48687 45702
rect 49820 45685 50160 45717
rect 48765 45639 48778 45685
rect 48824 45639 48881 45685
rect 48927 45639 48984 45685
rect 49030 45639 49087 45685
rect 49133 45639 49190 45685
rect 49236 45639 49293 45685
rect 49339 45639 49396 45685
rect 49442 45639 49499 45685
rect 49545 45639 49602 45685
rect 49852 45639 50160 45685
rect 51589 45722 51657 45774
rect 51797 45754 52105 45776
rect 49820 45598 50160 45639
rect 50262 45615 50812 45656
rect 48557 45559 48687 45562
rect 44901 45523 45241 45552
rect 48557 45507 48596 45559
rect 48648 45507 48687 45559
rect 50262 45563 50300 45615
rect 50352 45598 50511 45615
rect 50563 45598 50722 45615
rect 50352 45563 50467 45598
rect 50563 45563 50571 45598
rect 50262 45552 50467 45563
rect 50513 45552 50571 45563
rect 50617 45552 50674 45598
rect 50720 45563 50722 45598
rect 50774 45598 50812 45615
rect 50774 45563 50777 45598
rect 50720 45552 50777 45563
rect 50823 45552 50880 45598
rect 50926 45552 50983 45598
rect 51029 45552 51086 45598
rect 51132 45552 51189 45598
rect 51235 45552 51292 45598
rect 51338 45552 51395 45598
rect 51441 45552 51454 45598
rect 50262 45523 50812 45552
rect 48557 45466 48687 45507
rect 48905 45461 49877 45492
rect 48765 45415 48778 45461
rect 48824 45415 48881 45461
rect 48927 45452 48984 45461
rect 48927 45415 48943 45452
rect 49030 45415 49087 45461
rect 49133 45452 49190 45461
rect 49133 45415 49154 45452
rect 49236 45415 49293 45461
rect 49339 45452 49396 45461
rect 49339 45415 49365 45452
rect 49442 45415 49499 45461
rect 49545 45452 49602 45461
rect 49545 45415 49576 45452
rect 49852 45415 49877 45461
rect 48905 45400 48943 45415
rect 48995 45400 49154 45415
rect 49206 45400 49365 45415
rect 49417 45400 49576 45415
rect 49628 45400 49787 45415
rect 49839 45400 49877 45415
rect 44605 45328 44812 45374
rect 44858 45328 44925 45374
rect 44971 45328 45038 45374
rect 45084 45328 45151 45374
rect 45197 45328 45264 45374
rect 45310 45328 45323 45374
rect 48905 45360 49877 45400
rect 51035 45377 51343 45417
rect 51035 45374 51073 45377
rect 51125 45374 51253 45377
rect 51305 45374 51343 45377
rect 43362 45291 43524 45298
rect 43362 45245 43373 45291
rect 43513 45245 43524 45291
rect 43362 45234 43524 45245
rect 45584 45314 48546 45350
rect 50454 45328 50467 45374
rect 50513 45328 50571 45374
rect 50617 45328 50674 45374
rect 50720 45328 50777 45374
rect 50823 45328 50880 45374
rect 50926 45328 50983 45374
rect 51029 45328 51073 45374
rect 51132 45328 51189 45374
rect 51235 45328 51253 45374
rect 51338 45328 51395 45374
rect 51441 45328 51454 45374
rect 45584 45268 45619 45314
rect 45665 45268 45777 45314
rect 45823 45268 45935 45314
rect 45981 45268 46093 45314
rect 46139 45268 46251 45314
rect 46297 45268 46409 45314
rect 46455 45268 46568 45314
rect 46614 45268 46726 45314
rect 46772 45268 46884 45314
rect 46930 45268 47042 45314
rect 47088 45268 47200 45314
rect 47246 45268 47358 45314
rect 47404 45268 47516 45314
rect 47562 45268 47675 45314
rect 47721 45268 47833 45314
rect 47879 45268 47991 45314
rect 48037 45268 48149 45314
rect 48195 45268 48307 45314
rect 48353 45268 48465 45314
rect 48511 45268 48546 45314
rect 51035 45325 51073 45328
rect 51125 45325 51253 45328
rect 51305 45325 51343 45328
rect 51035 45284 51343 45325
rect 51589 45300 51600 45722
rect 51646 45300 51657 45722
rect 54085 45723 54540 45841
rect 54085 45677 54440 45723
rect 54486 45677 54540 45723
rect 54085 45649 54540 45677
rect 53585 45598 54540 45649
rect 51789 45552 51802 45598
rect 53776 45560 54540 45598
rect 53776 45552 54440 45560
rect 53585 45530 54440 45552
rect 54085 45514 54440 45530
rect 54486 45514 54540 45560
rect 54085 45438 54540 45514
rect 51797 45384 52105 45424
rect 51797 45374 51835 45384
rect 51887 45374 52015 45384
rect 52067 45374 52105 45384
rect 54085 45392 54223 45438
rect 54269 45397 54540 45438
rect 54269 45392 54440 45397
rect 51789 45328 51802 45374
rect 53776 45328 53789 45374
rect 54085 45351 54440 45392
rect 54486 45351 54540 45397
rect 51589 45289 51657 45300
rect 51797 45291 52105 45328
rect 40215 45187 40523 45194
rect 40788 45187 42986 45201
rect 43753 45187 44514 45194
rect 39492 45164 42986 45187
rect 43704 45164 44514 45187
rect 39492 45153 44514 45164
rect 39492 45150 40253 45153
rect 39492 45104 39740 45150
rect 39786 45104 39862 45150
rect 39908 45104 39985 45150
rect 40031 45104 40108 45150
rect 40154 45104 40253 45150
rect 39492 45101 40253 45104
rect 40305 45101 40433 45153
rect 40485 45150 43790 45153
rect 40485 45104 40836 45150
rect 40882 45104 40994 45150
rect 41040 45104 41152 45150
rect 41198 45104 41310 45150
rect 41356 45104 41469 45150
rect 41515 45104 41627 45150
rect 41673 45104 41785 45150
rect 41831 45104 41943 45150
rect 41989 45104 42101 45150
rect 42147 45104 42259 45150
rect 42305 45104 42418 45150
rect 42464 45104 42576 45150
rect 42622 45104 42734 45150
rect 42780 45104 42892 45150
rect 42938 45104 43739 45150
rect 43785 45104 43790 45150
rect 40485 45101 43790 45104
rect 43842 45150 44001 45153
rect 43842 45104 43906 45150
rect 43952 45104 44001 45150
rect 43842 45101 44001 45104
rect 44053 45150 44213 45153
rect 44265 45150 44424 45153
rect 44053 45104 44071 45150
rect 44117 45104 44213 45150
rect 44282 45104 44424 45150
rect 44053 45101 44213 45104
rect 44265 45101 44424 45104
rect 44476 45101 44514 45153
rect 39492 45090 44514 45101
rect 39492 45067 42986 45090
rect 43704 45067 44514 45090
rect 39492 44615 39608 45067
rect 40215 45060 40523 45067
rect 40788 45053 42986 45067
rect 43753 45060 44514 45067
rect 44796 45187 45346 45194
rect 45584 45187 48546 45268
rect 54085 45274 54540 45351
rect 54085 45228 54223 45274
rect 54269 45234 54540 45274
rect 54269 45228 54440 45234
rect 54085 45194 54440 45228
rect 48800 45187 49982 45194
rect 50308 45187 50859 45194
rect 44796 45153 49982 45187
rect 44796 45150 44834 45153
rect 44886 45150 45045 45153
rect 45097 45150 45256 45153
rect 45308 45150 48838 45153
rect 44796 45104 44812 45150
rect 44886 45104 44925 45150
rect 44971 45104 45038 45150
rect 45097 45104 45151 45150
rect 45197 45104 45256 45150
rect 45310 45104 45619 45150
rect 45665 45104 45777 45150
rect 45823 45104 45935 45150
rect 45981 45104 46093 45150
rect 46139 45104 46251 45150
rect 46297 45104 46409 45150
rect 46455 45104 46568 45150
rect 46614 45104 46726 45150
rect 46772 45104 46884 45150
rect 46930 45104 47042 45150
rect 47088 45104 47200 45150
rect 47246 45104 47358 45150
rect 47404 45104 47516 45150
rect 47562 45104 47675 45150
rect 47721 45104 47833 45150
rect 47879 45104 47991 45150
rect 48037 45104 48149 45150
rect 48195 45104 48307 45150
rect 48353 45104 48465 45150
rect 48511 45104 48838 45150
rect 44796 45101 44834 45104
rect 44886 45101 45045 45104
rect 45097 45101 45256 45104
rect 45308 45101 48838 45104
rect 48890 45101 49048 45153
rect 49100 45101 49259 45153
rect 49311 45101 49471 45153
rect 49523 45101 49682 45153
rect 49734 45101 49892 45153
rect 49944 45101 49982 45153
rect 44796 45067 49982 45101
rect 50307 45153 50859 45187
rect 50307 45101 50346 45153
rect 50398 45150 50557 45153
rect 50609 45150 50768 45153
rect 50820 45150 50859 45153
rect 52278 45188 54440 45194
rect 54486 45188 54540 45234
rect 55927 45887 57736 46001
rect 55927 45844 56267 45887
rect 55927 45798 55961 45844
rect 56007 45841 56267 45844
rect 56313 45841 57736 45887
rect 56007 45798 57736 45841
rect 55927 45723 57736 45798
rect 55927 45681 56267 45723
rect 55927 45635 55961 45681
rect 56007 45677 56267 45681
rect 56313 45677 57736 45723
rect 56007 45635 57736 45677
rect 55927 45560 57736 45635
rect 55927 45517 56267 45560
rect 55927 45471 55961 45517
rect 56007 45514 56267 45517
rect 56313 45514 57736 45560
rect 56007 45471 57736 45514
rect 55927 45397 57736 45471
rect 55927 45354 56267 45397
rect 55927 45308 55961 45354
rect 56007 45351 56267 45354
rect 56313 45351 57736 45397
rect 56007 45308 57736 45351
rect 55927 45234 57736 45308
rect 52278 45153 54540 45188
rect 52278 45150 52316 45153
rect 52368 45150 52527 45153
rect 52579 45150 52738 45153
rect 52790 45150 52948 45153
rect 53000 45150 53159 45153
rect 53211 45150 53371 45153
rect 53423 45150 53582 45153
rect 53634 45150 53792 45153
rect 50398 45104 50467 45150
rect 50513 45104 50557 45150
rect 50617 45104 50674 45150
rect 50720 45104 50768 45150
rect 50823 45104 50880 45150
rect 50926 45104 50983 45150
rect 51029 45104 51086 45150
rect 51132 45104 51189 45150
rect 51235 45104 51292 45150
rect 51338 45104 51395 45150
rect 51441 45104 51454 45150
rect 51789 45104 51802 45150
rect 53776 45104 53792 45150
rect 50398 45101 50557 45104
rect 50609 45101 50768 45104
rect 50820 45101 50859 45104
rect 50307 45067 50859 45101
rect 44796 45060 45346 45067
rect 43362 45009 43524 45020
rect 39737 44926 39866 44955
rect 40246 44937 40362 44974
rect 43362 44963 43373 45009
rect 43513 44963 43524 45009
rect 43362 44956 43524 44963
rect 39727 44880 39740 44926
rect 39786 44915 39862 44926
rect 39827 44880 39862 44915
rect 39908 44880 39985 44926
rect 40031 44880 40108 44926
rect 40154 44880 40167 44926
rect 40246 44891 40281 44937
rect 40327 44891 40362 44937
rect 39737 44863 39775 44880
rect 39827 44863 39866 44880
rect 39737 44836 39866 44863
rect 39737 44823 39865 44836
rect 39923 44700 40085 44740
rect 39923 44648 39994 44700
rect 40046 44648 40085 44700
rect 39008 44569 39021 44615
rect 39067 44569 39144 44615
rect 39190 44569 39267 44615
rect 39313 44569 39326 44615
rect 39492 44569 39641 44615
rect 39687 44569 39730 44615
rect 39014 44537 39323 44569
rect 39492 44537 39608 44569
rect 37853 44425 38161 44430
rect 36438 44391 36953 44425
rect 37439 44391 38161 44425
rect 38658 44405 38726 44527
rect 39923 44517 40085 44648
rect 39809 44514 40085 44517
rect 39809 44506 39994 44514
rect 39809 44460 39844 44506
rect 39890 44462 39994 44506
rect 40046 44493 40085 44514
rect 40246 44493 40362 44891
rect 40718 44915 43524 44956
rect 45584 44986 48546 45067
rect 48800 45060 49982 45067
rect 50308 45060 50859 45067
rect 52278 45101 52316 45104
rect 52368 45101 52527 45104
rect 52579 45101 52738 45104
rect 52790 45101 52948 45104
rect 53000 45101 53159 45104
rect 53211 45101 53371 45104
rect 53423 45101 53582 45104
rect 53634 45101 53792 45104
rect 53844 45101 54003 45153
rect 54055 45101 54214 45153
rect 54266 45101 54540 45153
rect 52278 45066 54540 45101
rect 52278 45060 54440 45066
rect 45584 44940 45619 44986
rect 45665 44940 45777 44986
rect 45823 44940 45935 44986
rect 45981 44940 46093 44986
rect 46139 44940 46251 44986
rect 46297 44940 46409 44986
rect 46455 44940 46568 44986
rect 46614 44940 46726 44986
rect 46772 44940 46884 44986
rect 46930 44940 47042 44986
rect 47088 44940 47200 44986
rect 47246 44940 47358 44986
rect 47404 44940 47516 44986
rect 47562 44940 47675 44986
rect 47721 44940 47833 44986
rect 47879 44940 47991 44986
rect 48037 44940 48149 44986
rect 48195 44940 48307 44986
rect 48353 44940 48465 44986
rect 48511 44940 48546 44986
rect 54085 45026 54440 45060
rect 54085 44980 54223 45026
rect 54269 45020 54440 45026
rect 54486 45020 54540 45066
rect 54758 45153 55840 45194
rect 54758 45150 54855 45153
rect 54758 45104 54793 45150
rect 54839 45104 54855 45150
rect 54758 45101 54855 45104
rect 54907 45150 55066 45153
rect 54907 45104 54956 45150
rect 55002 45104 55066 45150
rect 54907 45101 55066 45104
rect 55118 45150 55278 45153
rect 55330 45150 55489 45153
rect 55164 45104 55278 45150
rect 55330 45104 55439 45150
rect 55485 45104 55489 45150
rect 55118 45101 55278 45104
rect 55330 45101 55489 45104
rect 55541 45150 55840 45153
rect 55541 45104 55599 45150
rect 55645 45104 55760 45150
rect 55806 45104 55840 45150
rect 55541 45101 55840 45104
rect 54758 45061 55840 45101
rect 55927 45188 56267 45234
rect 56313 45188 57736 45234
rect 55927 45066 57736 45188
rect 54817 45060 55579 45061
rect 54269 44980 54540 45020
rect 40718 44863 41935 44915
rect 41987 44863 43524 44915
rect 40718 44822 43524 44863
rect 44605 44880 44812 44926
rect 44858 44880 44925 44926
rect 44971 44880 45038 44926
rect 45084 44880 45151 44926
rect 45197 44880 45264 44926
rect 45310 44880 45323 44926
rect 45584 44904 48546 44940
rect 51035 44929 51343 44970
rect 51035 44926 51073 44929
rect 51125 44926 51253 44929
rect 51305 44926 51343 44929
rect 51589 44954 51657 44965
rect 44341 44814 44509 44825
rect 44341 44768 44358 44814
rect 44498 44768 44509 44814
rect 44341 44724 44509 44768
rect 42229 44684 44509 44724
rect 42229 44632 43068 44684
rect 43120 44632 44509 44684
rect 42229 44591 44509 44632
rect 44605 44493 44721 44880
rect 48905 44854 49877 44894
rect 50454 44880 50467 44926
rect 50513 44880 50571 44926
rect 50617 44880 50674 44926
rect 50720 44880 50777 44926
rect 50823 44880 50880 44926
rect 50926 44880 50983 44926
rect 51029 44880 51073 44926
rect 51132 44880 51189 44926
rect 51235 44880 51253 44926
rect 51338 44880 51395 44926
rect 51441 44880 51454 44926
rect 48905 44839 48943 44854
rect 48995 44839 49154 44854
rect 49206 44839 49365 44854
rect 49417 44839 49576 44854
rect 49628 44839 49787 44854
rect 49839 44839 49877 44854
rect 48765 44793 48778 44839
rect 48824 44793 48881 44839
rect 48927 44802 48943 44839
rect 48927 44793 48984 44802
rect 49030 44793 49087 44839
rect 49133 44802 49154 44839
rect 49133 44793 49190 44802
rect 49236 44793 49293 44839
rect 49339 44802 49365 44839
rect 49339 44793 49396 44802
rect 49442 44793 49499 44839
rect 49545 44802 49576 44839
rect 49545 44793 49602 44802
rect 49852 44793 49877 44839
rect 51035 44877 51073 44880
rect 51125 44877 51253 44880
rect 51305 44877 51343 44880
rect 51035 44837 51343 44877
rect 48557 44747 48687 44788
rect 48905 44762 49877 44793
rect 44901 44702 45241 44731
rect 44799 44656 44812 44702
rect 44858 44656 44925 44702
rect 44971 44691 45038 44702
rect 44991 44656 45038 44691
rect 45084 44656 45151 44702
rect 45197 44691 45264 44702
rect 45203 44656 45264 44691
rect 45310 44656 45323 44702
rect 48557 44695 48596 44747
rect 48648 44695 48687 44747
rect 48557 44692 48687 44695
rect 44901 44639 44939 44656
rect 44991 44639 45151 44656
rect 45203 44639 45241 44656
rect 44901 44598 45241 44639
rect 45400 44583 48379 44616
rect 45400 44537 45464 44583
rect 45604 44575 48379 44583
rect 45604 44537 47864 44575
rect 45400 44523 47864 44537
rect 47916 44523 48379 44575
rect 40046 44478 44918 44493
rect 45400 44482 48379 44523
rect 48557 44552 48622 44692
rect 48668 44552 48687 44692
rect 50262 44702 50812 44731
rect 50262 44691 50467 44702
rect 50513 44691 50571 44702
rect 49820 44615 50160 44656
rect 48765 44569 48778 44615
rect 48824 44569 48881 44615
rect 48927 44569 48984 44615
rect 49030 44569 49087 44615
rect 49133 44569 49190 44615
rect 49236 44569 49293 44615
rect 49339 44569 49396 44615
rect 49442 44569 49499 44615
rect 49545 44569 49602 44615
rect 49852 44569 50160 44615
rect 50262 44639 50300 44691
rect 50352 44656 50467 44691
rect 50563 44656 50571 44691
rect 50617 44656 50674 44702
rect 50720 44691 50777 44702
rect 50720 44656 50722 44691
rect 50352 44639 50511 44656
rect 50563 44639 50722 44656
rect 50774 44656 50777 44691
rect 50823 44656 50880 44702
rect 50926 44656 50983 44702
rect 51029 44656 51086 44702
rect 51132 44656 51189 44702
rect 51235 44656 51292 44702
rect 51338 44656 51395 44702
rect 51441 44656 51454 44702
rect 50774 44639 50812 44656
rect 50262 44598 50812 44639
rect 48557 44529 48687 44552
rect 49820 44537 50160 44569
rect 40046 44462 44812 44478
rect 39890 44460 44812 44462
rect 39809 44457 44812 44460
rect 39809 44411 43739 44457
rect 43785 44411 43906 44457
rect 43952 44411 44071 44457
rect 44117 44411 44236 44457
rect 44282 44432 44812 44457
rect 44858 44432 44925 44478
rect 44971 44432 45038 44478
rect 45084 44432 45151 44478
rect 45197 44432 45264 44478
rect 45310 44432 45323 44478
rect 48557 44477 48596 44529
rect 48648 44477 48687 44529
rect 48557 44437 48687 44477
rect 50044 44480 50160 44537
rect 51589 44532 51600 44954
rect 51646 44532 51657 44954
rect 51797 44926 52105 44963
rect 51789 44880 51802 44926
rect 53776 44880 53789 44926
rect 54085 44903 54540 44980
rect 51797 44870 51835 44880
rect 51887 44870 52015 44880
rect 52067 44870 52105 44880
rect 51797 44830 52105 44870
rect 54085 44862 54440 44903
rect 54085 44816 54223 44862
rect 54269 44857 54440 44862
rect 54486 44857 54540 44903
rect 54269 44816 54540 44857
rect 54085 44740 54540 44816
rect 54085 44724 54440 44740
rect 53585 44702 54440 44724
rect 51789 44656 51802 44702
rect 53776 44694 54440 44702
rect 54486 44694 54540 44740
rect 53776 44656 54540 44694
rect 53585 44605 54540 44656
rect 51589 44480 51657 44532
rect 54085 44577 54540 44605
rect 54085 44531 54440 44577
rect 54486 44531 54540 44577
rect 50044 44443 51657 44480
rect 51797 44478 52105 44500
rect 44282 44411 44918 44432
rect 38658 44391 39723 44405
rect 30683 44367 30855 44373
rect 30583 44327 30855 44367
rect 30901 44327 31040 44373
rect 33484 44360 34643 44389
rect 35260 44345 35273 44391
rect 35523 44345 35543 44391
rect 35626 44345 35683 44391
rect 35729 44345 35754 44391
rect 35832 44345 35889 44391
rect 35935 44345 35965 44391
rect 36038 44345 36095 44391
rect 36141 44345 36176 44391
rect 36244 44345 36301 44391
rect 36347 44345 36360 44391
rect 36438 44345 36854 44391
rect 36900 44345 36971 44391
rect 37017 44345 37088 44391
rect 37134 44345 37206 44391
rect 37252 44345 37324 44391
rect 37370 44345 37442 44391
rect 37488 44389 37909 44391
rect 37488 44345 37891 44389
rect 37955 44345 38026 44391
rect 38072 44389 38143 44391
rect 38123 44345 38143 44389
rect 38189 44345 38261 44391
rect 38307 44345 38379 44391
rect 38425 44345 38497 44391
rect 38543 44345 38556 44391
rect 38658 44345 39021 44391
rect 39067 44345 39144 44391
rect 39190 44345 39267 44391
rect 39313 44345 39641 44391
rect 39687 44345 39730 44391
rect 39809 44373 44918 44411
rect 48905 44391 49877 44431
rect 48765 44345 48778 44391
rect 48824 44345 48881 44391
rect 48927 44345 48943 44391
rect 49030 44345 49087 44391
rect 49133 44345 49154 44391
rect 49236 44345 49293 44391
rect 49339 44345 49365 44391
rect 49442 44345 49499 44391
rect 49545 44345 49576 44391
rect 49852 44345 49877 44391
rect 50044 44397 50516 44443
rect 50562 44397 50703 44443
rect 50749 44397 50890 44443
rect 50936 44397 51076 44443
rect 51122 44397 51263 44443
rect 51309 44397 51657 44443
rect 51789 44432 51802 44478
rect 53776 44432 53789 44478
rect 50044 44387 51657 44397
rect 50481 44360 51657 44387
rect 51797 44407 51835 44432
rect 51887 44407 52015 44432
rect 52067 44407 52105 44432
rect 51797 44367 52105 44407
rect 54085 44413 54540 44531
rect 54085 44373 54440 44413
rect 30583 44294 31040 44327
rect 35294 44339 35332 44345
rect 35384 44339 35543 44345
rect 35595 44339 35754 44345
rect 35806 44339 35965 44345
rect 36017 44339 36176 44345
rect 36228 44339 36266 44345
rect 34870 44294 35025 44301
rect 35294 44299 36266 44339
rect 36438 44305 36953 44345
rect 37439 44337 37891 44345
rect 37943 44337 38071 44345
rect 38123 44337 38161 44345
rect 37439 44305 38161 44337
rect 37853 44297 38161 44305
rect 27387 44201 27790 44253
rect 27842 44201 28001 44253
rect 28053 44201 28212 44253
rect 28264 44201 28423 44253
rect 28475 44201 28634 44253
rect 28686 44250 28845 44253
rect 28686 44204 28810 44250
rect 28686 44201 28845 44204
rect 28897 44201 29056 44253
rect 29108 44201 29196 44253
rect 27387 44087 29196 44201
rect 29283 44253 30365 44294
rect 29283 44250 29582 44253
rect 29283 44204 29317 44250
rect 29363 44204 29478 44250
rect 29524 44204 29582 44250
rect 29283 44201 29582 44204
rect 29634 44250 29793 44253
rect 29845 44250 30005 44253
rect 29634 44204 29638 44250
rect 29684 44204 29793 44250
rect 29845 44204 29959 44250
rect 29634 44201 29793 44204
rect 29845 44201 30005 44204
rect 30057 44250 30216 44253
rect 30057 44204 30121 44250
rect 30167 44204 30216 44250
rect 30057 44201 30216 44204
rect 30268 44250 30365 44253
rect 30268 44204 30284 44250
rect 30330 44204 30365 44250
rect 30268 44201 30365 44204
rect 29283 44161 30365 44201
rect 30583 44253 32842 44294
rect 30583 44250 30854 44253
rect 30583 44204 30637 44250
rect 30683 44204 30854 44250
rect 30583 44201 30854 44204
rect 30906 44201 31065 44253
rect 31117 44201 31276 44253
rect 31328 44201 31486 44253
rect 31538 44201 31697 44253
rect 31749 44201 31909 44253
rect 31961 44201 32120 44253
rect 32172 44201 32330 44253
rect 32382 44201 32541 44253
rect 32593 44201 32752 44253
rect 32804 44201 32842 44253
rect 29544 44160 30306 44161
rect 30583 44160 32842 44201
rect 34717 44253 35025 44294
rect 38658 44285 39723 44345
rect 48905 44339 48943 44345
rect 48995 44339 49154 44345
rect 49206 44339 49365 44345
rect 49417 44339 49576 44345
rect 49628 44339 49787 44345
rect 49839 44339 49877 44345
rect 48905 44299 49877 44339
rect 54085 44327 54223 44373
rect 54269 44367 54440 44373
rect 54486 44367 54540 44413
rect 54269 44327 54540 44367
rect 50099 44294 50255 44301
rect 54085 44294 54540 44327
rect 55927 45020 56267 45066
rect 56313 45020 57736 45066
rect 55927 44944 57736 45020
rect 55927 44898 55961 44944
rect 56007 44903 57736 44944
rect 56007 44898 56267 44903
rect 55927 44857 56267 44898
rect 56313 44857 57736 44903
rect 55927 44781 57736 44857
rect 55927 44735 55961 44781
rect 56007 44740 57736 44781
rect 56007 44735 56267 44740
rect 55927 44694 56267 44735
rect 56313 44694 57736 44740
rect 55927 44617 57736 44694
rect 55927 44571 55961 44617
rect 56007 44577 57736 44617
rect 56007 44571 56267 44577
rect 55927 44531 56267 44571
rect 56313 44531 57736 44577
rect 55927 44454 57736 44531
rect 55927 44408 55961 44454
rect 56007 44413 57736 44454
rect 56007 44408 56267 44413
rect 55927 44367 56267 44408
rect 56313 44367 57736 44413
rect 34717 44201 34755 44253
rect 34807 44250 34935 44253
rect 34807 44204 34916 44250
rect 34807 44201 34935 44204
rect 34987 44201 35025 44253
rect 34717 44160 35025 44201
rect 50099 44253 50408 44294
rect 50099 44201 50138 44253
rect 50190 44250 50318 44253
rect 50206 44204 50318 44250
rect 50190 44201 50318 44204
rect 50370 44201 50408 44253
rect 27387 44041 28810 44087
rect 28856 44044 29196 44087
rect 28856 44041 29116 44044
rect 27387 43998 29116 44041
rect 29162 43998 29196 44044
rect 27387 43923 29196 43998
rect 27387 43877 28810 43923
rect 28856 43881 29196 43923
rect 28856 43877 29116 43881
rect 27387 43835 29116 43877
rect 29162 43835 29196 43881
rect 27387 43760 29196 43835
rect 27387 43714 28810 43760
rect 28856 43717 29196 43760
rect 28856 43714 29116 43717
rect 27387 43671 29116 43714
rect 29162 43671 29196 43717
rect 27387 43597 29196 43671
rect 27387 43551 28810 43597
rect 28856 43554 29196 43597
rect 28856 43551 29116 43554
rect 27387 43508 29116 43551
rect 29162 43508 29196 43554
rect 27387 43434 29196 43508
rect 27387 43388 28810 43434
rect 28856 43388 29196 43434
rect 30583 44127 31040 44160
rect 34870 44153 35025 44160
rect 30583 44087 30855 44127
rect 30583 44041 30637 44087
rect 30683 44081 30855 44087
rect 30901 44081 31040 44127
rect 35294 44115 36266 44155
rect 37853 44149 38161 44157
rect 35294 44109 35332 44115
rect 35384 44109 35543 44115
rect 35595 44109 35754 44115
rect 35806 44109 35965 44115
rect 36017 44109 36176 44115
rect 36228 44109 36266 44115
rect 36438 44109 36953 44149
rect 37439 44117 38161 44149
rect 37439 44109 37891 44117
rect 37943 44109 38071 44117
rect 38123 44109 38161 44117
rect 38658 44109 39723 44169
rect 50099 44160 50408 44201
rect 52278 44253 54540 44294
rect 52278 44201 52316 44253
rect 52368 44201 52527 44253
rect 52579 44201 52738 44253
rect 52790 44201 52948 44253
rect 53000 44201 53159 44253
rect 53211 44201 53371 44253
rect 53423 44201 53582 44253
rect 53634 44201 53792 44253
rect 53844 44201 54003 44253
rect 54055 44201 54214 44253
rect 54266 44250 54540 44253
rect 54266 44204 54440 44250
rect 54486 44204 54540 44250
rect 54266 44201 54540 44204
rect 52278 44160 54540 44201
rect 54758 44253 55840 44294
rect 54758 44250 54855 44253
rect 54758 44204 54793 44250
rect 54839 44204 54855 44250
rect 54758 44201 54855 44204
rect 54907 44250 55066 44253
rect 54907 44204 54956 44250
rect 55002 44204 55066 44250
rect 54907 44201 55066 44204
rect 55118 44250 55278 44253
rect 55330 44250 55489 44253
rect 55164 44204 55278 44250
rect 55330 44204 55439 44250
rect 55485 44204 55489 44250
rect 55118 44201 55278 44204
rect 55330 44201 55489 44204
rect 55541 44250 55840 44253
rect 55541 44204 55599 44250
rect 55645 44204 55760 44250
rect 55806 44204 55840 44250
rect 55541 44201 55840 44204
rect 54758 44161 55840 44201
rect 55927 44253 57736 44367
rect 55927 44201 56015 44253
rect 56067 44201 56226 44253
rect 56278 44250 56437 44253
rect 56313 44204 56437 44250
rect 56278 44201 56437 44204
rect 56489 44201 56648 44253
rect 56700 44201 56859 44253
rect 56911 44201 57070 44253
rect 57122 44201 57281 44253
rect 57333 44201 57736 44253
rect 54817 44160 55579 44161
rect 48905 44115 49877 44155
rect 50099 44153 50255 44160
rect 48905 44109 48943 44115
rect 48995 44109 49154 44115
rect 49206 44109 49365 44115
rect 49417 44109 49576 44115
rect 49628 44109 49787 44115
rect 49839 44109 49877 44115
rect 30683 44041 31040 44081
rect 33484 44065 34643 44094
rect 30583 43964 31040 44041
rect 33019 44025 33327 44065
rect 33019 44022 33057 44025
rect 33109 44022 33237 44025
rect 33289 44022 33327 44025
rect 33484 44057 35082 44065
rect 35260 44063 35273 44109
rect 35523 44063 35543 44109
rect 35626 44063 35683 44109
rect 35729 44063 35754 44109
rect 35832 44063 35889 44109
rect 35935 44063 35965 44109
rect 36038 44063 36095 44109
rect 36141 44063 36176 44109
rect 36244 44063 36301 44109
rect 36347 44063 36360 44109
rect 36438 44063 36854 44109
rect 36900 44063 36971 44109
rect 37017 44063 37088 44109
rect 37134 44063 37206 44109
rect 37252 44063 37324 44109
rect 37370 44063 37442 44109
rect 37488 44065 37891 44109
rect 37488 44063 37909 44065
rect 37955 44063 38026 44109
rect 38123 44065 38143 44109
rect 38072 44063 38143 44065
rect 38189 44063 38261 44109
rect 38307 44063 38379 44109
rect 38425 44063 38497 44109
rect 38543 44063 38556 44109
rect 38658 44063 39021 44109
rect 39067 44063 39144 44109
rect 39190 44063 39267 44109
rect 39313 44063 39641 44109
rect 39687 44063 39730 44109
rect 31336 43976 31349 44022
rect 33323 43976 33336 44022
rect 33484 44011 33816 44057
rect 33862 44011 34002 44057
rect 34048 44011 34189 44057
rect 34235 44011 34376 44057
rect 34422 44011 34562 44057
rect 34608 44011 35082 44057
rect 35294 44023 36266 44063
rect 36438 44029 36953 44063
rect 37439 44029 38161 44063
rect 30583 43923 30855 43964
rect 30583 43877 30637 43923
rect 30683 43918 30855 43923
rect 30901 43918 31040 43964
rect 33019 43973 33057 43976
rect 33109 43973 33237 43976
rect 33289 43973 33327 43976
rect 33019 43932 33327 43973
rect 33484 43974 35082 44011
rect 30683 43877 31040 43918
rect 30583 43849 31040 43877
rect 33484 43892 33552 43974
rect 30583 43801 31493 43849
rect 30583 43760 30855 43801
rect 30583 43714 30637 43760
rect 30683 43755 30855 43760
rect 30901 43798 31493 43801
rect 30901 43755 31349 43798
rect 30683 43752 31349 43755
rect 33323 43752 33336 43798
rect 30683 43730 31493 43752
rect 30683 43714 31040 43730
rect 30583 43638 31040 43714
rect 30583 43597 30855 43638
rect 30583 43551 30637 43597
rect 30683 43592 30855 43597
rect 30901 43592 31040 43638
rect 30683 43551 31040 43592
rect 33019 43577 33327 43617
rect 33019 43574 33057 43577
rect 33109 43574 33237 43577
rect 33289 43574 33327 43577
rect 30583 43474 31040 43551
rect 31336 43528 31349 43574
rect 33323 43528 33336 43574
rect 33019 43525 33057 43528
rect 33109 43525 33237 43528
rect 33289 43525 33327 43528
rect 33019 43484 33327 43525
rect 30583 43434 30855 43474
rect 27387 43266 29196 43388
rect 27387 43220 28810 43266
rect 28856 43220 29196 43266
rect 29283 43353 30365 43394
rect 29283 43350 29582 43353
rect 29283 43304 29317 43350
rect 29363 43304 29478 43350
rect 29524 43304 29582 43350
rect 29283 43301 29582 43304
rect 29634 43350 29793 43353
rect 29845 43350 30005 43353
rect 29634 43304 29638 43350
rect 29684 43304 29793 43350
rect 29845 43304 29959 43350
rect 29634 43301 29793 43304
rect 29845 43301 30005 43304
rect 30057 43350 30216 43353
rect 30057 43304 30121 43350
rect 30167 43304 30216 43350
rect 30057 43301 30216 43304
rect 30268 43350 30365 43353
rect 30268 43304 30284 43350
rect 30330 43304 30365 43350
rect 30268 43301 30365 43304
rect 29283 43261 30365 43301
rect 30583 43388 30637 43434
rect 30683 43428 30855 43434
rect 30901 43428 31040 43474
rect 33484 43470 33495 43892
rect 33541 43470 33552 43892
rect 34964 43917 35082 43974
rect 36438 43929 36554 44029
rect 37853 44024 38161 44029
rect 38658 44049 39723 44063
rect 34964 43885 36360 43917
rect 34228 43815 34718 43856
rect 34228 43798 34267 43815
rect 34319 43798 34447 43815
rect 34499 43798 34627 43815
rect 33671 43752 33684 43798
rect 33730 43752 33787 43798
rect 33833 43752 33890 43798
rect 33936 43752 33993 43798
rect 34039 43752 34096 43798
rect 34142 43752 34199 43798
rect 34245 43763 34267 43798
rect 34245 43752 34302 43763
rect 34348 43752 34405 43798
rect 34499 43763 34508 43798
rect 34451 43752 34508 43763
rect 34554 43752 34612 43798
rect 34679 43763 34718 43815
rect 34964 43839 35273 43885
rect 35523 43839 35580 43885
rect 35626 43839 35683 43885
rect 35729 43839 35786 43885
rect 35832 43839 35889 43885
rect 35935 43839 35992 43885
rect 36038 43839 36095 43885
rect 36141 43839 36198 43885
rect 36244 43839 36301 43885
rect 36347 43839 36360 43885
rect 34964 43795 36360 43839
rect 34658 43752 34718 43763
rect 34228 43723 34718 43752
rect 36438 43789 36475 43929
rect 36521 43789 36554 43929
rect 35294 43661 36266 43695
rect 36438 43686 36554 43789
rect 36640 43929 36773 43949
rect 36640 43890 36697 43929
rect 36640 43838 36678 43890
rect 36640 43789 36697 43838
rect 36743 43789 36773 43929
rect 38658 43927 38726 44049
rect 39809 44043 44918 44081
rect 48765 44063 48778 44109
rect 48824 44063 48881 44109
rect 48927 44063 48943 44109
rect 49030 44063 49087 44109
rect 49133 44063 49154 44109
rect 49236 44063 49293 44109
rect 49339 44063 49365 44109
rect 49442 44063 49499 44109
rect 49545 44063 49576 44109
rect 49852 44063 49877 44109
rect 54085 44127 54540 44160
rect 50481 44067 51657 44094
rect 39809 43997 43739 44043
rect 43785 43997 43906 44043
rect 43952 43997 44071 44043
rect 44117 43997 44236 44043
rect 44282 44022 44918 44043
rect 48905 44023 49877 44063
rect 50044 44057 51657 44067
rect 44282 43997 44812 44022
rect 39809 43994 44812 43997
rect 39809 43948 39844 43994
rect 39890 43992 44812 43994
rect 39890 43948 39994 43992
rect 39809 43940 39994 43948
rect 40046 43976 44812 43992
rect 44858 43976 44925 44022
rect 44971 43976 45038 44022
rect 45084 43976 45151 44022
rect 45197 43976 45264 44022
rect 45310 43976 45323 44022
rect 48557 43977 48687 44017
rect 40046 43961 44918 43976
rect 40046 43940 40085 43961
rect 39809 43937 40085 43940
rect 36924 43917 37685 43924
rect 36923 43885 37931 43917
rect 36841 43839 36854 43885
rect 36900 43883 36971 43885
rect 36900 43839 36961 43883
rect 37017 43839 37088 43885
rect 37134 43883 37206 43885
rect 37134 43839 37172 43883
rect 37252 43839 37324 43885
rect 37370 43883 37442 43885
rect 37370 43839 37384 43883
rect 36923 43831 36961 43839
rect 37013 43831 37172 43839
rect 37224 43831 37384 43839
rect 37436 43839 37442 43883
rect 37488 43883 37909 43885
rect 37488 43839 37595 43883
rect 37436 43831 37595 43839
rect 37647 43839 37909 43883
rect 37955 43839 38026 43885
rect 38072 43839 38143 43885
rect 38189 43839 38261 43885
rect 38307 43839 38379 43885
rect 38425 43839 38497 43885
rect 38543 43839 38556 43885
rect 37647 43831 37931 43839
rect 36923 43798 37931 43831
rect 36923 43797 37685 43798
rect 36924 43791 37685 43797
rect 36640 43766 36773 43789
rect 38658 43787 38669 43927
rect 38715 43787 38726 43927
rect 39014 43885 39323 43917
rect 39492 43885 39608 43917
rect 39008 43839 39021 43885
rect 39067 43839 39144 43885
rect 39190 43839 39267 43885
rect 39313 43839 39326 43885
rect 39492 43839 39641 43885
rect 39687 43839 39730 43885
rect 38658 43776 38726 43787
rect 36438 43661 36953 43686
rect 37439 43683 37931 43686
rect 37439 43661 38161 43683
rect 35260 43615 35273 43661
rect 35523 43655 35580 43661
rect 35523 43615 35543 43655
rect 35626 43615 35683 43661
rect 35729 43655 35786 43661
rect 35729 43615 35754 43655
rect 35832 43615 35889 43661
rect 35935 43655 35992 43661
rect 35935 43615 35965 43655
rect 36038 43615 36095 43661
rect 36141 43655 36198 43661
rect 36141 43615 36176 43655
rect 36244 43615 36301 43661
rect 36347 43615 36360 43661
rect 36438 43615 36854 43661
rect 36900 43615 36971 43661
rect 37017 43615 37088 43661
rect 37134 43615 37206 43661
rect 37252 43615 37324 43661
rect 37370 43615 37442 43661
rect 37488 43643 37909 43661
rect 37488 43615 37891 43643
rect 37955 43615 38026 43661
rect 38072 43643 38143 43661
rect 38123 43615 38143 43643
rect 38189 43615 38261 43661
rect 38307 43615 38379 43661
rect 38425 43615 38497 43661
rect 38543 43615 38556 43661
rect 33781 43574 34089 43609
rect 35294 43603 35332 43615
rect 35384 43603 35543 43615
rect 35595 43603 35754 43615
rect 35806 43603 35965 43615
rect 36017 43603 36176 43615
rect 36228 43603 36266 43615
rect 33671 43528 33684 43574
rect 33730 43528 33787 43574
rect 33833 43569 33890 43574
rect 33871 43528 33890 43569
rect 33936 43528 33993 43574
rect 34039 43569 34096 43574
rect 34051 43528 34096 43569
rect 34142 43528 34199 43574
rect 34245 43528 34302 43574
rect 34348 43528 34405 43574
rect 34451 43528 34508 43574
rect 34554 43528 34612 43574
rect 34658 43528 34671 43574
rect 35294 43563 36266 43603
rect 36438 43566 36953 43615
rect 37439 43591 37891 43615
rect 37943 43591 38071 43615
rect 38123 43591 38161 43615
rect 37439 43566 38161 43591
rect 37853 43550 38161 43566
rect 33781 43517 33819 43528
rect 33871 43517 33999 43528
rect 34051 43517 34089 43528
rect 33781 43476 34089 43517
rect 33484 43459 33552 43470
rect 30683 43394 31040 43428
rect 30683 43388 32842 43394
rect 30583 43353 32842 43388
rect 34247 43387 35008 43394
rect 30583 43301 30854 43353
rect 30906 43301 31065 43353
rect 31117 43301 31276 43353
rect 31328 43350 31486 43353
rect 31538 43350 31697 43353
rect 31749 43350 31909 43353
rect 31961 43350 32120 43353
rect 32172 43350 32330 43353
rect 32382 43350 32541 43353
rect 32593 43350 32752 43353
rect 32804 43350 32842 43353
rect 34246 43353 35008 43387
rect 34246 43350 34284 43353
rect 34336 43350 34495 43353
rect 34547 43350 34707 43353
rect 31328 43304 31349 43350
rect 33323 43304 33336 43350
rect 33671 43304 33684 43350
rect 33730 43304 33787 43350
rect 33833 43304 33890 43350
rect 33936 43304 33993 43350
rect 34039 43304 34096 43350
rect 34142 43304 34199 43350
rect 34245 43304 34284 43350
rect 34348 43304 34405 43350
rect 34451 43304 34495 43350
rect 34554 43304 34612 43350
rect 34658 43304 34707 43350
rect 31328 43301 31486 43304
rect 31538 43301 31697 43304
rect 31749 43301 31909 43304
rect 31961 43301 32120 43304
rect 32172 43301 32330 43304
rect 32382 43301 32541 43304
rect 32593 43301 32752 43304
rect 32804 43301 32842 43304
rect 30583 43266 32842 43301
rect 34246 43301 34284 43304
rect 34336 43301 34495 43304
rect 34547 43301 34707 43304
rect 34759 43301 34918 43353
rect 34970 43301 35008 43353
rect 34246 43267 35008 43301
rect 29544 43260 30306 43261
rect 27387 43144 29196 43220
rect 27387 43103 29116 43144
rect 27387 43057 28810 43103
rect 28856 43098 29116 43103
rect 29162 43098 29196 43144
rect 28856 43057 29196 43098
rect 27387 42981 29196 43057
rect 27387 42940 29116 42981
rect 27387 42894 28810 42940
rect 28856 42935 29116 42940
rect 29162 42935 29196 42981
rect 28856 42894 29196 42935
rect 27387 42817 29196 42894
rect 27387 42777 29116 42817
rect 27387 42731 28810 42777
rect 28856 42771 29116 42777
rect 29162 42771 29196 42817
rect 28856 42731 29196 42771
rect 27387 42654 29196 42731
rect 27387 42613 29116 42654
rect 27387 42567 28810 42613
rect 28856 42608 29116 42613
rect 29162 42608 29196 42654
rect 28856 42567 29196 42608
rect 27387 42453 29196 42567
rect 30583 43220 30637 43266
rect 30683 43260 32842 43266
rect 34247 43260 35008 43267
rect 35182 43387 36364 43394
rect 35182 43353 36958 43387
rect 35182 43301 35220 43353
rect 35272 43301 35430 43353
rect 35482 43301 35641 43353
rect 35693 43301 35853 43353
rect 35905 43301 36064 43353
rect 36116 43301 36274 43353
rect 36326 43350 36958 43353
rect 36326 43304 36489 43350
rect 36723 43304 36958 43350
rect 36326 43301 36958 43304
rect 35182 43267 36958 43301
rect 37946 43353 38842 43394
rect 37946 43350 38330 43353
rect 38382 43350 38541 43353
rect 37946 43304 37957 43350
rect 38473 43304 38541 43350
rect 37946 43301 38330 43304
rect 38382 43301 38541 43304
rect 38593 43301 38752 43353
rect 38804 43301 38842 43353
rect 35182 43260 36364 43267
rect 37946 43260 38842 43301
rect 39014 43353 39323 43839
rect 39014 43301 39052 43353
rect 39104 43350 39232 43353
rect 39108 43304 39220 43350
rect 39104 43301 39232 43304
rect 39284 43301 39323 43353
rect 30683 43226 31040 43260
rect 30683 43220 30855 43226
rect 30583 43180 30855 43220
rect 30901 43180 31040 43226
rect 30583 43103 31040 43180
rect 33484 43184 33552 43195
rect 33019 43129 33327 43170
rect 33019 43126 33057 43129
rect 33109 43126 33237 43129
rect 33289 43126 33327 43129
rect 30583 43057 30637 43103
rect 30683 43062 31040 43103
rect 31336 43080 31349 43126
rect 33323 43080 33336 43126
rect 30683 43057 30855 43062
rect 30583 43016 30855 43057
rect 30901 43016 31040 43062
rect 33019 43077 33057 43080
rect 33109 43077 33237 43080
rect 33289 43077 33327 43080
rect 33019 43037 33327 43077
rect 30583 42940 31040 43016
rect 30583 42894 30637 42940
rect 30683 42924 31040 42940
rect 30683 42902 31493 42924
rect 30683 42899 31349 42902
rect 30683 42894 30855 42899
rect 30583 42853 30855 42894
rect 30901 42856 31349 42899
rect 33323 42856 33336 42902
rect 30901 42853 31493 42856
rect 30583 42805 31493 42853
rect 30583 42777 31040 42805
rect 30583 42731 30637 42777
rect 30683 42736 31040 42777
rect 30683 42731 30855 42736
rect 30583 42690 30855 42731
rect 30901 42690 31040 42736
rect 33484 42762 33495 43184
rect 33541 42762 33552 43184
rect 33781 43137 34089 43178
rect 33781 43126 33819 43137
rect 33871 43126 33999 43137
rect 34051 43126 34089 43137
rect 33671 43080 33684 43126
rect 33730 43080 33787 43126
rect 33871 43085 33890 43126
rect 33833 43080 33890 43085
rect 33936 43080 33993 43126
rect 34051 43085 34096 43126
rect 34039 43080 34096 43085
rect 34142 43080 34199 43126
rect 34245 43080 34302 43126
rect 34348 43080 34405 43126
rect 34451 43080 34508 43126
rect 34554 43080 34612 43126
rect 34658 43080 34671 43126
rect 33781 43045 34089 43080
rect 35294 43051 36266 43091
rect 37853 43088 38161 43104
rect 35294 43039 35332 43051
rect 35384 43039 35543 43051
rect 35595 43039 35754 43051
rect 35806 43039 35965 43051
rect 36017 43039 36176 43051
rect 36228 43039 36266 43051
rect 36438 43039 36953 43088
rect 37439 43063 38161 43088
rect 37439 43039 37891 43063
rect 37943 43039 38071 43063
rect 38123 43039 38161 43063
rect 35260 42993 35273 43039
rect 35523 42999 35543 43039
rect 35523 42993 35580 42999
rect 35626 42993 35683 43039
rect 35729 42999 35754 43039
rect 35729 42993 35786 42999
rect 35832 42993 35889 43039
rect 35935 42999 35965 43039
rect 35935 42993 35992 42999
rect 36038 42993 36095 43039
rect 36141 42999 36176 43039
rect 36141 42993 36198 42999
rect 36244 42993 36301 43039
rect 36347 42993 36360 43039
rect 36438 42993 36854 43039
rect 36900 42993 36971 43039
rect 37017 42993 37088 43039
rect 37134 42993 37206 43039
rect 37252 42993 37324 43039
rect 37370 42993 37442 43039
rect 37488 43011 37891 43039
rect 37488 42993 37909 43011
rect 37955 42993 38026 43039
rect 38123 43011 38143 43039
rect 38072 42993 38143 43011
rect 38189 42993 38261 43039
rect 38307 42993 38379 43039
rect 38425 42993 38497 43039
rect 38543 42993 38556 43039
rect 35294 42959 36266 42993
rect 36438 42968 36953 42993
rect 37439 42971 38161 42993
rect 37439 42968 37931 42971
rect 34228 42902 34718 42931
rect 33671 42856 33684 42902
rect 33730 42856 33787 42902
rect 33833 42856 33890 42902
rect 33936 42856 33993 42902
rect 34039 42856 34096 42902
rect 34142 42856 34199 42902
rect 34245 42891 34302 42902
rect 34245 42856 34267 42891
rect 34348 42856 34405 42902
rect 34451 42891 34508 42902
rect 34499 42856 34508 42891
rect 34554 42856 34612 42902
rect 34658 42891 34718 42902
rect 34228 42839 34267 42856
rect 34319 42839 34447 42856
rect 34499 42839 34627 42856
rect 34679 42839 34718 42891
rect 36438 42865 36554 42968
rect 34228 42798 34718 42839
rect 34964 42815 36360 42859
rect 30583 42613 31040 42690
rect 33019 42681 33327 42722
rect 33019 42678 33057 42681
rect 33109 42678 33237 42681
rect 33289 42678 33327 42681
rect 33484 42680 33552 42762
rect 34964 42769 35273 42815
rect 35523 42769 35580 42815
rect 35626 42769 35683 42815
rect 35729 42769 35786 42815
rect 35832 42769 35889 42815
rect 35935 42769 35992 42815
rect 36038 42769 36095 42815
rect 36141 42769 36198 42815
rect 36244 42769 36301 42815
rect 36347 42769 36360 42815
rect 34964 42737 36360 42769
rect 34964 42680 35082 42737
rect 31336 42632 31349 42678
rect 33323 42632 33336 42678
rect 33484 42643 35082 42680
rect 30583 42567 30637 42613
rect 30683 42573 31040 42613
rect 33019 42629 33057 42632
rect 33109 42629 33237 42632
rect 33289 42629 33327 42632
rect 33019 42589 33327 42629
rect 33484 42597 33816 42643
rect 33862 42597 34002 42643
rect 34048 42597 34189 42643
rect 34235 42597 34376 42643
rect 34422 42597 34562 42643
rect 34608 42597 35082 42643
rect 36438 42725 36475 42865
rect 36521 42725 36554 42865
rect 33484 42589 35082 42597
rect 35294 42591 36266 42631
rect 36438 42625 36554 42725
rect 36640 42865 36773 42888
rect 36640 42816 36697 42865
rect 36640 42764 36678 42816
rect 36640 42725 36697 42764
rect 36743 42725 36773 42865
rect 38658 42867 38726 42878
rect 36924 42857 37685 42863
rect 36923 42856 37685 42857
rect 36923 42823 37931 42856
rect 36923 42815 36961 42823
rect 37013 42815 37172 42823
rect 37224 42815 37384 42823
rect 36841 42769 36854 42815
rect 36900 42771 36961 42815
rect 36900 42769 36971 42771
rect 37017 42769 37088 42815
rect 37134 42771 37172 42815
rect 37134 42769 37206 42771
rect 37252 42769 37324 42815
rect 37370 42771 37384 42815
rect 37436 42815 37595 42823
rect 37436 42771 37442 42815
rect 37370 42769 37442 42771
rect 37488 42771 37595 42815
rect 37647 42815 37931 42823
rect 37647 42771 37909 42815
rect 37488 42769 37909 42771
rect 37955 42769 38026 42815
rect 38072 42769 38143 42815
rect 38189 42769 38261 42815
rect 38307 42769 38379 42815
rect 38425 42769 38497 42815
rect 38543 42769 38556 42815
rect 36923 42737 37931 42769
rect 36924 42730 37685 42737
rect 36640 42705 36773 42725
rect 38658 42727 38669 42867
rect 38715 42727 38726 42867
rect 39014 42815 39323 43301
rect 39492 43387 39608 43839
rect 39923 43806 40085 43937
rect 39923 43754 39994 43806
rect 40046 43754 40085 43806
rect 39923 43714 40085 43754
rect 39737 43618 39865 43631
rect 39737 43591 39866 43618
rect 39737 43574 39775 43591
rect 39827 43574 39866 43591
rect 39727 43528 39740 43574
rect 39827 43539 39862 43574
rect 39786 43528 39862 43539
rect 39908 43528 39985 43574
rect 40031 43528 40108 43574
rect 40154 43528 40167 43574
rect 40246 43563 40362 43961
rect 42229 43822 44509 43863
rect 42229 43770 43068 43822
rect 43120 43770 44509 43822
rect 42229 43730 44509 43770
rect 44341 43686 44509 43730
rect 44341 43640 44358 43686
rect 44498 43640 44509 43686
rect 39737 43499 39866 43528
rect 40246 43517 40281 43563
rect 40327 43517 40362 43563
rect 40246 43480 40362 43517
rect 40718 43591 43524 43632
rect 44341 43629 44509 43640
rect 40718 43539 41935 43591
rect 41987 43539 43524 43591
rect 40718 43498 43524 43539
rect 44605 43574 44721 43961
rect 45400 43931 48379 43972
rect 45400 43917 48241 43931
rect 45400 43871 45464 43917
rect 45604 43879 48241 43917
rect 48293 43879 48379 43931
rect 45604 43871 48379 43879
rect 44901 43815 45241 43856
rect 45400 43838 48379 43871
rect 48557 43925 48596 43977
rect 48648 43925 48687 43977
rect 48557 43902 48687 43925
rect 50044 44011 50516 44057
rect 50562 44011 50703 44057
rect 50749 44011 50890 44057
rect 50936 44011 51076 44057
rect 51122 44011 51263 44057
rect 51309 44011 51657 44057
rect 51797 44047 52105 44087
rect 51797 44022 51835 44047
rect 51887 44022 52015 44047
rect 52067 44022 52105 44047
rect 54085 44081 54223 44127
rect 54269 44087 54540 44127
rect 54269 44081 54440 44087
rect 54085 44041 54440 44081
rect 54486 44041 54540 44087
rect 50044 43974 51657 44011
rect 51789 43976 51802 44022
rect 53776 43976 53789 44022
rect 50044 43917 50160 43974
rect 44901 43798 44939 43815
rect 44991 43798 45151 43815
rect 45203 43798 45241 43815
rect 44799 43752 44812 43798
rect 44858 43752 44925 43798
rect 44991 43763 45038 43798
rect 44971 43752 45038 43763
rect 45084 43752 45151 43798
rect 45203 43763 45264 43798
rect 45197 43752 45264 43763
rect 45310 43752 45323 43798
rect 48557 43762 48622 43902
rect 48668 43762 48687 43902
rect 49820 43885 50160 43917
rect 48765 43839 48778 43885
rect 48824 43839 48881 43885
rect 48927 43839 48984 43885
rect 49030 43839 49087 43885
rect 49133 43839 49190 43885
rect 49236 43839 49293 43885
rect 49339 43839 49396 43885
rect 49442 43839 49499 43885
rect 49545 43839 49602 43885
rect 49852 43839 50160 43885
rect 51589 43922 51657 43974
rect 51797 43954 52105 43976
rect 49820 43798 50160 43839
rect 50262 43815 50812 43856
rect 48557 43759 48687 43762
rect 44901 43723 45241 43752
rect 48557 43707 48596 43759
rect 48648 43707 48687 43759
rect 50262 43763 50300 43815
rect 50352 43798 50511 43815
rect 50563 43798 50722 43815
rect 50352 43763 50467 43798
rect 50563 43763 50571 43798
rect 50262 43752 50467 43763
rect 50513 43752 50571 43763
rect 50617 43752 50674 43798
rect 50720 43763 50722 43798
rect 50774 43798 50812 43815
rect 50774 43763 50777 43798
rect 50720 43752 50777 43763
rect 50823 43752 50880 43798
rect 50926 43752 50983 43798
rect 51029 43752 51086 43798
rect 51132 43752 51189 43798
rect 51235 43752 51292 43798
rect 51338 43752 51395 43798
rect 51441 43752 51454 43798
rect 50262 43723 50812 43752
rect 48557 43666 48687 43707
rect 48905 43661 49877 43692
rect 48765 43615 48778 43661
rect 48824 43615 48881 43661
rect 48927 43652 48984 43661
rect 48927 43615 48943 43652
rect 49030 43615 49087 43661
rect 49133 43652 49190 43661
rect 49133 43615 49154 43652
rect 49236 43615 49293 43661
rect 49339 43652 49396 43661
rect 49339 43615 49365 43652
rect 49442 43615 49499 43661
rect 49545 43652 49602 43661
rect 49545 43615 49576 43652
rect 49852 43615 49877 43661
rect 48905 43600 48943 43615
rect 48995 43600 49154 43615
rect 49206 43600 49365 43615
rect 49417 43600 49576 43615
rect 49628 43600 49787 43615
rect 49839 43600 49877 43615
rect 44605 43528 44812 43574
rect 44858 43528 44925 43574
rect 44971 43528 45038 43574
rect 45084 43528 45151 43574
rect 45197 43528 45264 43574
rect 45310 43528 45323 43574
rect 48905 43560 49877 43600
rect 51035 43577 51343 43617
rect 51035 43574 51073 43577
rect 51125 43574 51253 43577
rect 51305 43574 51343 43577
rect 43362 43491 43524 43498
rect 43362 43445 43373 43491
rect 43513 43445 43524 43491
rect 43362 43434 43524 43445
rect 45584 43514 48546 43550
rect 50454 43528 50467 43574
rect 50513 43528 50571 43574
rect 50617 43528 50674 43574
rect 50720 43528 50777 43574
rect 50823 43528 50880 43574
rect 50926 43528 50983 43574
rect 51029 43528 51073 43574
rect 51132 43528 51189 43574
rect 51235 43528 51253 43574
rect 51338 43528 51395 43574
rect 51441 43528 51454 43574
rect 45584 43468 45619 43514
rect 45665 43468 45777 43514
rect 45823 43468 45935 43514
rect 45981 43468 46093 43514
rect 46139 43468 46251 43514
rect 46297 43468 46409 43514
rect 46455 43468 46568 43514
rect 46614 43468 46726 43514
rect 46772 43468 46884 43514
rect 46930 43468 47042 43514
rect 47088 43468 47200 43514
rect 47246 43468 47358 43514
rect 47404 43468 47516 43514
rect 47562 43468 47675 43514
rect 47721 43468 47833 43514
rect 47879 43468 47991 43514
rect 48037 43468 48149 43514
rect 48195 43468 48307 43514
rect 48353 43468 48465 43514
rect 48511 43468 48546 43514
rect 51035 43525 51073 43528
rect 51125 43525 51253 43528
rect 51305 43525 51343 43528
rect 51035 43484 51343 43525
rect 51589 43500 51600 43922
rect 51646 43500 51657 43922
rect 54085 43923 54540 44041
rect 54085 43877 54440 43923
rect 54486 43877 54540 43923
rect 54085 43849 54540 43877
rect 53585 43798 54540 43849
rect 51789 43752 51802 43798
rect 53776 43760 54540 43798
rect 53776 43752 54440 43760
rect 53585 43730 54440 43752
rect 54085 43714 54440 43730
rect 54486 43714 54540 43760
rect 54085 43638 54540 43714
rect 51797 43584 52105 43624
rect 51797 43574 51835 43584
rect 51887 43574 52015 43584
rect 52067 43574 52105 43584
rect 54085 43592 54223 43638
rect 54269 43597 54540 43638
rect 54269 43592 54440 43597
rect 51789 43528 51802 43574
rect 53776 43528 53789 43574
rect 54085 43551 54440 43592
rect 54486 43551 54540 43597
rect 51589 43489 51657 43500
rect 51797 43491 52105 43528
rect 40215 43387 40523 43394
rect 40788 43387 42986 43401
rect 43753 43387 44514 43394
rect 39492 43364 42986 43387
rect 43704 43364 44514 43387
rect 39492 43353 44514 43364
rect 39492 43350 40253 43353
rect 39492 43304 39740 43350
rect 39786 43304 39862 43350
rect 39908 43304 39985 43350
rect 40031 43304 40108 43350
rect 40154 43304 40253 43350
rect 39492 43301 40253 43304
rect 40305 43301 40433 43353
rect 40485 43350 43790 43353
rect 40485 43304 40836 43350
rect 40882 43304 40994 43350
rect 41040 43304 41152 43350
rect 41198 43304 41310 43350
rect 41356 43304 41469 43350
rect 41515 43304 41627 43350
rect 41673 43304 41785 43350
rect 41831 43304 41943 43350
rect 41989 43304 42101 43350
rect 42147 43304 42259 43350
rect 42305 43304 42418 43350
rect 42464 43304 42576 43350
rect 42622 43304 42734 43350
rect 42780 43304 42892 43350
rect 42938 43304 43739 43350
rect 43785 43304 43790 43350
rect 40485 43301 43790 43304
rect 43842 43350 44001 43353
rect 43842 43304 43906 43350
rect 43952 43304 44001 43350
rect 43842 43301 44001 43304
rect 44053 43350 44213 43353
rect 44265 43350 44424 43353
rect 44053 43304 44071 43350
rect 44117 43304 44213 43350
rect 44282 43304 44424 43350
rect 44053 43301 44213 43304
rect 44265 43301 44424 43304
rect 44476 43301 44514 43353
rect 39492 43290 44514 43301
rect 39492 43267 42986 43290
rect 43704 43267 44514 43290
rect 39492 42815 39608 43267
rect 40215 43260 40523 43267
rect 40788 43253 42986 43267
rect 43753 43260 44514 43267
rect 44796 43387 45346 43394
rect 45584 43387 48546 43468
rect 54085 43474 54540 43551
rect 54085 43428 54223 43474
rect 54269 43434 54540 43474
rect 54269 43428 54440 43434
rect 54085 43394 54440 43428
rect 48800 43387 49982 43394
rect 50308 43387 50859 43394
rect 44796 43353 49982 43387
rect 44796 43350 44834 43353
rect 44886 43350 45045 43353
rect 45097 43350 45256 43353
rect 45308 43350 48838 43353
rect 44796 43304 44812 43350
rect 44886 43304 44925 43350
rect 44971 43304 45038 43350
rect 45097 43304 45151 43350
rect 45197 43304 45256 43350
rect 45310 43304 45619 43350
rect 45665 43304 45777 43350
rect 45823 43304 45935 43350
rect 45981 43304 46093 43350
rect 46139 43304 46251 43350
rect 46297 43304 46409 43350
rect 46455 43304 46568 43350
rect 46614 43304 46726 43350
rect 46772 43304 46884 43350
rect 46930 43304 47042 43350
rect 47088 43304 47200 43350
rect 47246 43304 47358 43350
rect 47404 43304 47516 43350
rect 47562 43304 47675 43350
rect 47721 43304 47833 43350
rect 47879 43304 47991 43350
rect 48037 43304 48149 43350
rect 48195 43304 48307 43350
rect 48353 43304 48465 43350
rect 48511 43304 48838 43350
rect 44796 43301 44834 43304
rect 44886 43301 45045 43304
rect 45097 43301 45256 43304
rect 45308 43301 48838 43304
rect 48890 43301 49048 43353
rect 49100 43301 49259 43353
rect 49311 43301 49471 43353
rect 49523 43301 49682 43353
rect 49734 43301 49892 43353
rect 49944 43301 49982 43353
rect 44796 43267 49982 43301
rect 50307 43353 50859 43387
rect 50307 43301 50346 43353
rect 50398 43350 50557 43353
rect 50609 43350 50768 43353
rect 50820 43350 50859 43353
rect 52278 43388 54440 43394
rect 54486 43388 54540 43434
rect 55927 44087 57736 44201
rect 55927 44044 56267 44087
rect 55927 43998 55961 44044
rect 56007 44041 56267 44044
rect 56313 44041 57736 44087
rect 56007 43998 57736 44041
rect 55927 43923 57736 43998
rect 55927 43881 56267 43923
rect 55927 43835 55961 43881
rect 56007 43877 56267 43881
rect 56313 43877 57736 43923
rect 56007 43835 57736 43877
rect 55927 43760 57736 43835
rect 55927 43717 56267 43760
rect 55927 43671 55961 43717
rect 56007 43714 56267 43717
rect 56313 43714 57736 43760
rect 56007 43671 57736 43714
rect 55927 43597 57736 43671
rect 55927 43554 56267 43597
rect 55927 43508 55961 43554
rect 56007 43551 56267 43554
rect 56313 43551 57736 43597
rect 56007 43508 57736 43551
rect 55927 43434 57736 43508
rect 52278 43353 54540 43388
rect 52278 43350 52316 43353
rect 52368 43350 52527 43353
rect 52579 43350 52738 43353
rect 52790 43350 52948 43353
rect 53000 43350 53159 43353
rect 53211 43350 53371 43353
rect 53423 43350 53582 43353
rect 53634 43350 53792 43353
rect 50398 43304 50467 43350
rect 50513 43304 50557 43350
rect 50617 43304 50674 43350
rect 50720 43304 50768 43350
rect 50823 43304 50880 43350
rect 50926 43304 50983 43350
rect 51029 43304 51086 43350
rect 51132 43304 51189 43350
rect 51235 43304 51292 43350
rect 51338 43304 51395 43350
rect 51441 43304 51454 43350
rect 51789 43304 51802 43350
rect 53776 43304 53792 43350
rect 50398 43301 50557 43304
rect 50609 43301 50768 43304
rect 50820 43301 50859 43304
rect 50307 43267 50859 43301
rect 44796 43260 45346 43267
rect 43362 43209 43524 43220
rect 39737 43126 39866 43155
rect 40246 43137 40362 43174
rect 43362 43163 43373 43209
rect 43513 43163 43524 43209
rect 43362 43156 43524 43163
rect 39727 43080 39740 43126
rect 39786 43115 39862 43126
rect 39827 43080 39862 43115
rect 39908 43080 39985 43126
rect 40031 43080 40108 43126
rect 40154 43080 40167 43126
rect 40246 43091 40281 43137
rect 40327 43091 40362 43137
rect 39737 43063 39775 43080
rect 39827 43063 39866 43080
rect 39737 43036 39866 43063
rect 39737 43023 39865 43036
rect 39923 42900 40085 42940
rect 39923 42848 39994 42900
rect 40046 42848 40085 42900
rect 39008 42769 39021 42815
rect 39067 42769 39144 42815
rect 39190 42769 39267 42815
rect 39313 42769 39326 42815
rect 39492 42769 39641 42815
rect 39687 42769 39730 42815
rect 39014 42737 39323 42769
rect 39492 42737 39608 42769
rect 37853 42625 38161 42630
rect 36438 42591 36953 42625
rect 37439 42591 38161 42625
rect 38658 42605 38726 42727
rect 39923 42717 40085 42848
rect 39809 42714 40085 42717
rect 39809 42706 39994 42714
rect 39809 42660 39844 42706
rect 39890 42662 39994 42706
rect 40046 42693 40085 42714
rect 40246 42693 40362 43091
rect 40718 43115 43524 43156
rect 45584 43186 48546 43267
rect 48800 43260 49982 43267
rect 50308 43260 50859 43267
rect 52278 43301 52316 43304
rect 52368 43301 52527 43304
rect 52579 43301 52738 43304
rect 52790 43301 52948 43304
rect 53000 43301 53159 43304
rect 53211 43301 53371 43304
rect 53423 43301 53582 43304
rect 53634 43301 53792 43304
rect 53844 43301 54003 43353
rect 54055 43301 54214 43353
rect 54266 43301 54540 43353
rect 52278 43266 54540 43301
rect 52278 43260 54440 43266
rect 45584 43140 45619 43186
rect 45665 43140 45777 43186
rect 45823 43140 45935 43186
rect 45981 43140 46093 43186
rect 46139 43140 46251 43186
rect 46297 43140 46409 43186
rect 46455 43140 46568 43186
rect 46614 43140 46726 43186
rect 46772 43140 46884 43186
rect 46930 43140 47042 43186
rect 47088 43140 47200 43186
rect 47246 43140 47358 43186
rect 47404 43140 47516 43186
rect 47562 43140 47675 43186
rect 47721 43140 47833 43186
rect 47879 43140 47991 43186
rect 48037 43140 48149 43186
rect 48195 43140 48307 43186
rect 48353 43140 48465 43186
rect 48511 43140 48546 43186
rect 54085 43226 54440 43260
rect 54085 43180 54223 43226
rect 54269 43220 54440 43226
rect 54486 43220 54540 43266
rect 54758 43353 55840 43394
rect 54758 43350 54855 43353
rect 54758 43304 54793 43350
rect 54839 43304 54855 43350
rect 54758 43301 54855 43304
rect 54907 43350 55066 43353
rect 54907 43304 54956 43350
rect 55002 43304 55066 43350
rect 54907 43301 55066 43304
rect 55118 43350 55278 43353
rect 55330 43350 55489 43353
rect 55164 43304 55278 43350
rect 55330 43304 55439 43350
rect 55485 43304 55489 43350
rect 55118 43301 55278 43304
rect 55330 43301 55489 43304
rect 55541 43350 55840 43353
rect 55541 43304 55599 43350
rect 55645 43304 55760 43350
rect 55806 43304 55840 43350
rect 55541 43301 55840 43304
rect 54758 43261 55840 43301
rect 55927 43388 56267 43434
rect 56313 43388 57736 43434
rect 55927 43266 57736 43388
rect 54817 43260 55579 43261
rect 54269 43180 54540 43220
rect 40718 43063 41935 43115
rect 41987 43063 43524 43115
rect 40718 43022 43524 43063
rect 44605 43080 44812 43126
rect 44858 43080 44925 43126
rect 44971 43080 45038 43126
rect 45084 43080 45151 43126
rect 45197 43080 45264 43126
rect 45310 43080 45323 43126
rect 45584 43104 48546 43140
rect 51035 43129 51343 43170
rect 51035 43126 51073 43129
rect 51125 43126 51253 43129
rect 51305 43126 51343 43129
rect 51589 43154 51657 43165
rect 44341 43014 44509 43025
rect 44341 42968 44358 43014
rect 44498 42968 44509 43014
rect 44341 42924 44509 42968
rect 42229 42884 44509 42924
rect 42229 42832 43445 42884
rect 43497 42832 44509 42884
rect 42229 42791 44509 42832
rect 44605 42693 44721 43080
rect 48905 43054 49877 43094
rect 50454 43080 50467 43126
rect 50513 43080 50571 43126
rect 50617 43080 50674 43126
rect 50720 43080 50777 43126
rect 50823 43080 50880 43126
rect 50926 43080 50983 43126
rect 51029 43080 51073 43126
rect 51132 43080 51189 43126
rect 51235 43080 51253 43126
rect 51338 43080 51395 43126
rect 51441 43080 51454 43126
rect 48905 43039 48943 43054
rect 48995 43039 49154 43054
rect 49206 43039 49365 43054
rect 49417 43039 49576 43054
rect 49628 43039 49787 43054
rect 49839 43039 49877 43054
rect 48765 42993 48778 43039
rect 48824 42993 48881 43039
rect 48927 43002 48943 43039
rect 48927 42993 48984 43002
rect 49030 42993 49087 43039
rect 49133 43002 49154 43039
rect 49133 42993 49190 43002
rect 49236 42993 49293 43039
rect 49339 43002 49365 43039
rect 49339 42993 49396 43002
rect 49442 42993 49499 43039
rect 49545 43002 49576 43039
rect 49545 42993 49602 43002
rect 49852 42993 49877 43039
rect 51035 43077 51073 43080
rect 51125 43077 51253 43080
rect 51305 43077 51343 43080
rect 51035 43037 51343 43077
rect 48557 42947 48687 42988
rect 48905 42962 49877 42993
rect 44901 42902 45241 42931
rect 44799 42856 44812 42902
rect 44858 42856 44925 42902
rect 44971 42891 45038 42902
rect 44991 42856 45038 42891
rect 45084 42856 45151 42902
rect 45197 42891 45264 42902
rect 45203 42856 45264 42891
rect 45310 42856 45323 42902
rect 48557 42895 48596 42947
rect 48648 42895 48687 42947
rect 48557 42892 48687 42895
rect 44901 42839 44939 42856
rect 44991 42839 45151 42856
rect 45203 42839 45241 42856
rect 44901 42798 45241 42839
rect 45400 42783 48379 42816
rect 45400 42737 45464 42783
rect 45604 42775 48379 42783
rect 45400 42723 45597 42737
rect 45649 42723 48379 42775
rect 40046 42678 44918 42693
rect 45400 42682 48379 42723
rect 48557 42752 48622 42892
rect 48668 42752 48687 42892
rect 50262 42902 50812 42931
rect 50262 42891 50467 42902
rect 50513 42891 50571 42902
rect 49820 42815 50160 42856
rect 48765 42769 48778 42815
rect 48824 42769 48881 42815
rect 48927 42769 48984 42815
rect 49030 42769 49087 42815
rect 49133 42769 49190 42815
rect 49236 42769 49293 42815
rect 49339 42769 49396 42815
rect 49442 42769 49499 42815
rect 49545 42769 49602 42815
rect 49852 42769 50160 42815
rect 50262 42839 50300 42891
rect 50352 42856 50467 42891
rect 50563 42856 50571 42891
rect 50617 42856 50674 42902
rect 50720 42891 50777 42902
rect 50720 42856 50722 42891
rect 50352 42839 50511 42856
rect 50563 42839 50722 42856
rect 50774 42856 50777 42891
rect 50823 42856 50880 42902
rect 50926 42856 50983 42902
rect 51029 42856 51086 42902
rect 51132 42856 51189 42902
rect 51235 42856 51292 42902
rect 51338 42856 51395 42902
rect 51441 42856 51454 42902
rect 50774 42839 50812 42856
rect 50262 42798 50812 42839
rect 48557 42729 48687 42752
rect 49820 42737 50160 42769
rect 40046 42662 44812 42678
rect 39890 42660 44812 42662
rect 39809 42657 44812 42660
rect 39809 42611 43739 42657
rect 43785 42611 43906 42657
rect 43952 42611 44071 42657
rect 44117 42611 44236 42657
rect 44282 42632 44812 42657
rect 44858 42632 44925 42678
rect 44971 42632 45038 42678
rect 45084 42632 45151 42678
rect 45197 42632 45264 42678
rect 45310 42632 45323 42678
rect 48557 42677 48596 42729
rect 48648 42677 48687 42729
rect 48557 42637 48687 42677
rect 50044 42680 50160 42737
rect 51589 42732 51600 43154
rect 51646 42732 51657 43154
rect 51797 43126 52105 43163
rect 51789 43080 51802 43126
rect 53776 43080 53789 43126
rect 54085 43103 54540 43180
rect 51797 43070 51835 43080
rect 51887 43070 52015 43080
rect 52067 43070 52105 43080
rect 51797 43030 52105 43070
rect 54085 43062 54440 43103
rect 54085 43016 54223 43062
rect 54269 43057 54440 43062
rect 54486 43057 54540 43103
rect 54269 43016 54540 43057
rect 54085 42940 54540 43016
rect 54085 42924 54440 42940
rect 53585 42902 54440 42924
rect 51789 42856 51802 42902
rect 53776 42894 54440 42902
rect 54486 42894 54540 42940
rect 53776 42856 54540 42894
rect 53585 42805 54540 42856
rect 51589 42680 51657 42732
rect 54085 42777 54540 42805
rect 54085 42731 54440 42777
rect 54486 42731 54540 42777
rect 50044 42643 51657 42680
rect 51797 42678 52105 42700
rect 44282 42611 44918 42632
rect 38658 42591 39723 42605
rect 30683 42567 30855 42573
rect 30583 42527 30855 42567
rect 30901 42527 31040 42573
rect 33484 42560 34643 42589
rect 35260 42545 35273 42591
rect 35523 42545 35543 42591
rect 35626 42545 35683 42591
rect 35729 42545 35754 42591
rect 35832 42545 35889 42591
rect 35935 42545 35965 42591
rect 36038 42545 36095 42591
rect 36141 42545 36176 42591
rect 36244 42545 36301 42591
rect 36347 42545 36360 42591
rect 36438 42545 36854 42591
rect 36900 42545 36971 42591
rect 37017 42545 37088 42591
rect 37134 42545 37206 42591
rect 37252 42545 37324 42591
rect 37370 42545 37442 42591
rect 37488 42589 37909 42591
rect 37488 42545 37891 42589
rect 37955 42545 38026 42591
rect 38072 42589 38143 42591
rect 38123 42545 38143 42589
rect 38189 42545 38261 42591
rect 38307 42545 38379 42591
rect 38425 42545 38497 42591
rect 38543 42545 38556 42591
rect 38658 42545 39021 42591
rect 39067 42545 39144 42591
rect 39190 42545 39267 42591
rect 39313 42545 39641 42591
rect 39687 42545 39730 42591
rect 39809 42573 44918 42611
rect 48905 42591 49877 42631
rect 48765 42545 48778 42591
rect 48824 42545 48881 42591
rect 48927 42545 48943 42591
rect 49030 42545 49087 42591
rect 49133 42545 49154 42591
rect 49236 42545 49293 42591
rect 49339 42545 49365 42591
rect 49442 42545 49499 42591
rect 49545 42545 49576 42591
rect 49852 42545 49877 42591
rect 50044 42597 50516 42643
rect 50562 42597 50703 42643
rect 50749 42597 50890 42643
rect 50936 42597 51076 42643
rect 51122 42597 51263 42643
rect 51309 42597 51657 42643
rect 51789 42632 51802 42678
rect 53776 42632 53789 42678
rect 50044 42587 51657 42597
rect 50481 42560 51657 42587
rect 51797 42607 51835 42632
rect 51887 42607 52015 42632
rect 52067 42607 52105 42632
rect 51797 42567 52105 42607
rect 54085 42613 54540 42731
rect 54085 42573 54440 42613
rect 30583 42494 31040 42527
rect 35294 42539 35332 42545
rect 35384 42539 35543 42545
rect 35595 42539 35754 42545
rect 35806 42539 35965 42545
rect 36017 42539 36176 42545
rect 36228 42539 36266 42545
rect 34870 42494 35025 42501
rect 35294 42499 36266 42539
rect 36438 42505 36953 42545
rect 37439 42537 37891 42545
rect 37943 42537 38071 42545
rect 38123 42537 38161 42545
rect 37439 42505 38161 42537
rect 37853 42497 38161 42505
rect 27387 42401 27790 42453
rect 27842 42401 28001 42453
rect 28053 42401 28212 42453
rect 28264 42401 28423 42453
rect 28475 42401 28634 42453
rect 28686 42450 28845 42453
rect 28686 42404 28810 42450
rect 28686 42401 28845 42404
rect 28897 42401 29056 42453
rect 29108 42401 29196 42453
rect 27387 42287 29196 42401
rect 29283 42453 30365 42494
rect 29283 42450 29582 42453
rect 29283 42404 29317 42450
rect 29363 42404 29478 42450
rect 29524 42404 29582 42450
rect 29283 42401 29582 42404
rect 29634 42450 29793 42453
rect 29845 42450 30005 42453
rect 29634 42404 29638 42450
rect 29684 42404 29793 42450
rect 29845 42404 29959 42450
rect 29634 42401 29793 42404
rect 29845 42401 30005 42404
rect 30057 42450 30216 42453
rect 30057 42404 30121 42450
rect 30167 42404 30216 42450
rect 30057 42401 30216 42404
rect 30268 42450 30365 42453
rect 30268 42404 30284 42450
rect 30330 42404 30365 42450
rect 30268 42401 30365 42404
rect 29283 42361 30365 42401
rect 30583 42453 32842 42494
rect 30583 42450 30854 42453
rect 30583 42404 30637 42450
rect 30683 42404 30854 42450
rect 30583 42401 30854 42404
rect 30906 42401 31065 42453
rect 31117 42401 31276 42453
rect 31328 42401 31486 42453
rect 31538 42401 31697 42453
rect 31749 42401 31909 42453
rect 31961 42401 32120 42453
rect 32172 42401 32330 42453
rect 32382 42401 32541 42453
rect 32593 42401 32752 42453
rect 32804 42401 32842 42453
rect 29544 42360 30306 42361
rect 30583 42360 32842 42401
rect 34717 42453 35025 42494
rect 38658 42485 39723 42545
rect 48905 42539 48943 42545
rect 48995 42539 49154 42545
rect 49206 42539 49365 42545
rect 49417 42539 49576 42545
rect 49628 42539 49787 42545
rect 49839 42539 49877 42545
rect 48905 42499 49877 42539
rect 54085 42527 54223 42573
rect 54269 42567 54440 42573
rect 54486 42567 54540 42613
rect 54269 42527 54540 42567
rect 50099 42494 50255 42501
rect 54085 42494 54540 42527
rect 55927 43220 56267 43266
rect 56313 43220 57736 43266
rect 55927 43144 57736 43220
rect 55927 43098 55961 43144
rect 56007 43103 57736 43144
rect 56007 43098 56267 43103
rect 55927 43057 56267 43098
rect 56313 43057 57736 43103
rect 55927 42981 57736 43057
rect 55927 42935 55961 42981
rect 56007 42940 57736 42981
rect 56007 42935 56267 42940
rect 55927 42894 56267 42935
rect 56313 42894 57736 42940
rect 55927 42817 57736 42894
rect 55927 42771 55961 42817
rect 56007 42777 57736 42817
rect 56007 42771 56267 42777
rect 55927 42731 56267 42771
rect 56313 42731 57736 42777
rect 55927 42654 57736 42731
rect 55927 42608 55961 42654
rect 56007 42613 57736 42654
rect 56007 42608 56267 42613
rect 55927 42567 56267 42608
rect 56313 42567 57736 42613
rect 34717 42401 34755 42453
rect 34807 42450 34935 42453
rect 34807 42404 34916 42450
rect 34807 42401 34935 42404
rect 34987 42401 35025 42453
rect 34717 42360 35025 42401
rect 50099 42453 50408 42494
rect 50099 42401 50138 42453
rect 50190 42450 50318 42453
rect 50206 42404 50318 42450
rect 50190 42401 50318 42404
rect 50370 42401 50408 42453
rect 27387 42241 28810 42287
rect 28856 42244 29196 42287
rect 28856 42241 29116 42244
rect 27387 42198 29116 42241
rect 29162 42198 29196 42244
rect 27387 42123 29196 42198
rect 27387 42077 28810 42123
rect 28856 42081 29196 42123
rect 28856 42077 29116 42081
rect 27387 42035 29116 42077
rect 29162 42035 29196 42081
rect 27387 41960 29196 42035
rect 27387 41914 28810 41960
rect 28856 41917 29196 41960
rect 28856 41914 29116 41917
rect 27387 41871 29116 41914
rect 29162 41871 29196 41917
rect 27387 41797 29196 41871
rect 27387 41751 28810 41797
rect 28856 41754 29196 41797
rect 28856 41751 29116 41754
rect 27387 41708 29116 41751
rect 29162 41708 29196 41754
rect 27387 41634 29196 41708
rect 27387 41588 28810 41634
rect 28856 41588 29196 41634
rect 30583 42327 31040 42360
rect 34870 42353 35025 42360
rect 30583 42287 30855 42327
rect 30583 42241 30637 42287
rect 30683 42281 30855 42287
rect 30901 42281 31040 42327
rect 35294 42315 36266 42355
rect 37853 42349 38161 42357
rect 35294 42309 35332 42315
rect 35384 42309 35543 42315
rect 35595 42309 35754 42315
rect 35806 42309 35965 42315
rect 36017 42309 36176 42315
rect 36228 42309 36266 42315
rect 36438 42309 36953 42349
rect 37439 42317 38161 42349
rect 37439 42309 37891 42317
rect 37943 42309 38071 42317
rect 38123 42309 38161 42317
rect 38658 42309 39723 42369
rect 50099 42360 50408 42401
rect 52278 42453 54540 42494
rect 52278 42401 52316 42453
rect 52368 42401 52527 42453
rect 52579 42401 52738 42453
rect 52790 42401 52948 42453
rect 53000 42401 53159 42453
rect 53211 42401 53371 42453
rect 53423 42401 53582 42453
rect 53634 42401 53792 42453
rect 53844 42401 54003 42453
rect 54055 42401 54214 42453
rect 54266 42450 54540 42453
rect 54266 42404 54440 42450
rect 54486 42404 54540 42450
rect 54266 42401 54540 42404
rect 52278 42360 54540 42401
rect 54758 42453 55840 42494
rect 54758 42450 54855 42453
rect 54758 42404 54793 42450
rect 54839 42404 54855 42450
rect 54758 42401 54855 42404
rect 54907 42450 55066 42453
rect 54907 42404 54956 42450
rect 55002 42404 55066 42450
rect 54907 42401 55066 42404
rect 55118 42450 55278 42453
rect 55330 42450 55489 42453
rect 55164 42404 55278 42450
rect 55330 42404 55439 42450
rect 55485 42404 55489 42450
rect 55118 42401 55278 42404
rect 55330 42401 55489 42404
rect 55541 42450 55840 42453
rect 55541 42404 55599 42450
rect 55645 42404 55760 42450
rect 55806 42404 55840 42450
rect 55541 42401 55840 42404
rect 54758 42361 55840 42401
rect 55927 42453 57736 42567
rect 55927 42401 56015 42453
rect 56067 42401 56226 42453
rect 56278 42450 56437 42453
rect 56313 42404 56437 42450
rect 56278 42401 56437 42404
rect 56489 42401 56648 42453
rect 56700 42401 56859 42453
rect 56911 42401 57070 42453
rect 57122 42401 57281 42453
rect 57333 42401 57736 42453
rect 54817 42360 55579 42361
rect 48905 42315 49877 42355
rect 50099 42353 50255 42360
rect 48905 42309 48943 42315
rect 48995 42309 49154 42315
rect 49206 42309 49365 42315
rect 49417 42309 49576 42315
rect 49628 42309 49787 42315
rect 49839 42309 49877 42315
rect 30683 42241 31040 42281
rect 33484 42265 34643 42294
rect 30583 42164 31040 42241
rect 33019 42225 33327 42265
rect 33019 42222 33057 42225
rect 33109 42222 33237 42225
rect 33289 42222 33327 42225
rect 33484 42257 35082 42265
rect 35260 42263 35273 42309
rect 35523 42263 35543 42309
rect 35626 42263 35683 42309
rect 35729 42263 35754 42309
rect 35832 42263 35889 42309
rect 35935 42263 35965 42309
rect 36038 42263 36095 42309
rect 36141 42263 36176 42309
rect 36244 42263 36301 42309
rect 36347 42263 36360 42309
rect 36438 42263 36854 42309
rect 36900 42263 36971 42309
rect 37017 42263 37088 42309
rect 37134 42263 37206 42309
rect 37252 42263 37324 42309
rect 37370 42263 37442 42309
rect 37488 42265 37891 42309
rect 37488 42263 37909 42265
rect 37955 42263 38026 42309
rect 38123 42265 38143 42309
rect 38072 42263 38143 42265
rect 38189 42263 38261 42309
rect 38307 42263 38379 42309
rect 38425 42263 38497 42309
rect 38543 42263 38556 42309
rect 38658 42263 39021 42309
rect 39067 42263 39144 42309
rect 39190 42263 39267 42309
rect 39313 42263 39641 42309
rect 39687 42263 39730 42309
rect 31336 42176 31349 42222
rect 33323 42176 33336 42222
rect 33484 42211 33816 42257
rect 33862 42211 34002 42257
rect 34048 42211 34189 42257
rect 34235 42211 34376 42257
rect 34422 42211 34562 42257
rect 34608 42211 35082 42257
rect 35294 42223 36266 42263
rect 36438 42229 36953 42263
rect 37439 42229 38161 42263
rect 30583 42123 30855 42164
rect 30583 42077 30637 42123
rect 30683 42118 30855 42123
rect 30901 42118 31040 42164
rect 33019 42173 33057 42176
rect 33109 42173 33237 42176
rect 33289 42173 33327 42176
rect 33019 42132 33327 42173
rect 33484 42174 35082 42211
rect 30683 42077 31040 42118
rect 30583 42049 31040 42077
rect 33484 42092 33552 42174
rect 30583 42001 31493 42049
rect 30583 41960 30855 42001
rect 30583 41914 30637 41960
rect 30683 41955 30855 41960
rect 30901 41998 31493 42001
rect 30901 41955 31349 41998
rect 30683 41952 31349 41955
rect 33323 41952 33336 41998
rect 30683 41930 31493 41952
rect 30683 41914 31040 41930
rect 30583 41838 31040 41914
rect 30583 41797 30855 41838
rect 30583 41751 30637 41797
rect 30683 41792 30855 41797
rect 30901 41792 31040 41838
rect 30683 41751 31040 41792
rect 33019 41777 33327 41817
rect 33019 41774 33057 41777
rect 33109 41774 33237 41777
rect 33289 41774 33327 41777
rect 30583 41674 31040 41751
rect 31336 41728 31349 41774
rect 33323 41728 33336 41774
rect 33019 41725 33057 41728
rect 33109 41725 33237 41728
rect 33289 41725 33327 41728
rect 33019 41684 33327 41725
rect 30583 41634 30855 41674
rect 27387 41466 29196 41588
rect 27387 41420 28810 41466
rect 28856 41420 29196 41466
rect 29283 41553 30365 41594
rect 29283 41550 29582 41553
rect 29283 41504 29317 41550
rect 29363 41504 29478 41550
rect 29524 41504 29582 41550
rect 29283 41501 29582 41504
rect 29634 41550 29793 41553
rect 29845 41550 30005 41553
rect 29634 41504 29638 41550
rect 29684 41504 29793 41550
rect 29845 41504 29959 41550
rect 29634 41501 29793 41504
rect 29845 41501 30005 41504
rect 30057 41550 30216 41553
rect 30057 41504 30121 41550
rect 30167 41504 30216 41550
rect 30057 41501 30216 41504
rect 30268 41550 30365 41553
rect 30268 41504 30284 41550
rect 30330 41504 30365 41550
rect 30268 41501 30365 41504
rect 29283 41461 30365 41501
rect 30583 41588 30637 41634
rect 30683 41628 30855 41634
rect 30901 41628 31040 41674
rect 33484 41670 33495 42092
rect 33541 41670 33552 42092
rect 34964 42117 35082 42174
rect 36438 42129 36554 42229
rect 37853 42224 38161 42229
rect 38658 42249 39723 42263
rect 34964 42085 36360 42117
rect 34228 42015 34718 42056
rect 34228 41998 34267 42015
rect 34319 41998 34447 42015
rect 34499 41998 34627 42015
rect 33671 41952 33684 41998
rect 33730 41952 33787 41998
rect 33833 41952 33890 41998
rect 33936 41952 33993 41998
rect 34039 41952 34096 41998
rect 34142 41952 34199 41998
rect 34245 41963 34267 41998
rect 34245 41952 34302 41963
rect 34348 41952 34405 41998
rect 34499 41963 34508 41998
rect 34451 41952 34508 41963
rect 34554 41952 34612 41998
rect 34679 41963 34718 42015
rect 34964 42039 35273 42085
rect 35523 42039 35580 42085
rect 35626 42039 35683 42085
rect 35729 42039 35786 42085
rect 35832 42039 35889 42085
rect 35935 42039 35992 42085
rect 36038 42039 36095 42085
rect 36141 42039 36198 42085
rect 36244 42039 36301 42085
rect 36347 42039 36360 42085
rect 34964 41995 36360 42039
rect 34658 41952 34718 41963
rect 34228 41923 34718 41952
rect 36438 41989 36475 42129
rect 36521 41989 36554 42129
rect 35294 41861 36266 41895
rect 36438 41886 36554 41989
rect 36640 42129 36773 42149
rect 36640 42090 36697 42129
rect 36640 42038 36678 42090
rect 36640 41989 36697 42038
rect 36743 41989 36773 42129
rect 38658 42127 38726 42249
rect 39809 42243 44918 42281
rect 48765 42263 48778 42309
rect 48824 42263 48881 42309
rect 48927 42263 48943 42309
rect 49030 42263 49087 42309
rect 49133 42263 49154 42309
rect 49236 42263 49293 42309
rect 49339 42263 49365 42309
rect 49442 42263 49499 42309
rect 49545 42263 49576 42309
rect 49852 42263 49877 42309
rect 54085 42327 54540 42360
rect 50481 42267 51657 42294
rect 39809 42197 43739 42243
rect 43785 42197 43906 42243
rect 43952 42197 44071 42243
rect 44117 42197 44236 42243
rect 44282 42222 44918 42243
rect 48905 42223 49877 42263
rect 50044 42257 51657 42267
rect 44282 42197 44812 42222
rect 39809 42194 44812 42197
rect 39809 42148 39844 42194
rect 39890 42192 44812 42194
rect 39890 42148 39994 42192
rect 39809 42140 39994 42148
rect 40046 42176 44812 42192
rect 44858 42176 44925 42222
rect 44971 42176 45038 42222
rect 45084 42176 45151 42222
rect 45197 42176 45264 42222
rect 45310 42176 45323 42222
rect 48557 42177 48687 42217
rect 40046 42161 44918 42176
rect 40046 42140 40085 42161
rect 39809 42137 40085 42140
rect 36924 42117 37685 42124
rect 36923 42085 37931 42117
rect 36841 42039 36854 42085
rect 36900 42083 36971 42085
rect 36900 42039 36961 42083
rect 37017 42039 37088 42085
rect 37134 42083 37206 42085
rect 37134 42039 37172 42083
rect 37252 42039 37324 42085
rect 37370 42083 37442 42085
rect 37370 42039 37384 42083
rect 36923 42031 36961 42039
rect 37013 42031 37172 42039
rect 37224 42031 37384 42039
rect 37436 42039 37442 42083
rect 37488 42083 37909 42085
rect 37488 42039 37595 42083
rect 37436 42031 37595 42039
rect 37647 42039 37909 42083
rect 37955 42039 38026 42085
rect 38072 42039 38143 42085
rect 38189 42039 38261 42085
rect 38307 42039 38379 42085
rect 38425 42039 38497 42085
rect 38543 42039 38556 42085
rect 37647 42031 37931 42039
rect 36923 41998 37931 42031
rect 36923 41997 37685 41998
rect 36924 41991 37685 41997
rect 36640 41966 36773 41989
rect 38658 41987 38669 42127
rect 38715 41987 38726 42127
rect 39014 42085 39323 42117
rect 39492 42085 39608 42117
rect 39008 42039 39021 42085
rect 39067 42039 39144 42085
rect 39190 42039 39267 42085
rect 39313 42039 39326 42085
rect 39492 42039 39641 42085
rect 39687 42039 39730 42085
rect 38658 41976 38726 41987
rect 36438 41861 36953 41886
rect 37439 41883 37931 41886
rect 37439 41861 38161 41883
rect 35260 41815 35273 41861
rect 35523 41855 35580 41861
rect 35523 41815 35543 41855
rect 35626 41815 35683 41861
rect 35729 41855 35786 41861
rect 35729 41815 35754 41855
rect 35832 41815 35889 41861
rect 35935 41855 35992 41861
rect 35935 41815 35965 41855
rect 36038 41815 36095 41861
rect 36141 41855 36198 41861
rect 36141 41815 36176 41855
rect 36244 41815 36301 41861
rect 36347 41815 36360 41861
rect 36438 41815 36854 41861
rect 36900 41815 36971 41861
rect 37017 41815 37088 41861
rect 37134 41815 37206 41861
rect 37252 41815 37324 41861
rect 37370 41815 37442 41861
rect 37488 41843 37909 41861
rect 37488 41815 37891 41843
rect 37955 41815 38026 41861
rect 38072 41843 38143 41861
rect 38123 41815 38143 41843
rect 38189 41815 38261 41861
rect 38307 41815 38379 41861
rect 38425 41815 38497 41861
rect 38543 41815 38556 41861
rect 33781 41774 34089 41809
rect 35294 41803 35332 41815
rect 35384 41803 35543 41815
rect 35595 41803 35754 41815
rect 35806 41803 35965 41815
rect 36017 41803 36176 41815
rect 36228 41803 36266 41815
rect 33671 41728 33684 41774
rect 33730 41728 33787 41774
rect 33833 41769 33890 41774
rect 33871 41728 33890 41769
rect 33936 41728 33993 41774
rect 34039 41769 34096 41774
rect 34051 41728 34096 41769
rect 34142 41728 34199 41774
rect 34245 41728 34302 41774
rect 34348 41728 34405 41774
rect 34451 41728 34508 41774
rect 34554 41728 34612 41774
rect 34658 41728 34671 41774
rect 35294 41763 36266 41803
rect 36438 41766 36953 41815
rect 37439 41791 37891 41815
rect 37943 41791 38071 41815
rect 38123 41791 38161 41815
rect 37439 41766 38161 41791
rect 37853 41750 38161 41766
rect 33781 41717 33819 41728
rect 33871 41717 33999 41728
rect 34051 41717 34089 41728
rect 33781 41676 34089 41717
rect 33484 41659 33552 41670
rect 30683 41594 31040 41628
rect 30683 41588 32842 41594
rect 30583 41553 32842 41588
rect 34247 41587 35008 41594
rect 30583 41501 30854 41553
rect 30906 41501 31065 41553
rect 31117 41501 31276 41553
rect 31328 41550 31486 41553
rect 31538 41550 31697 41553
rect 31749 41550 31909 41553
rect 31961 41550 32120 41553
rect 32172 41550 32330 41553
rect 32382 41550 32541 41553
rect 32593 41550 32752 41553
rect 32804 41550 32842 41553
rect 34246 41553 35008 41587
rect 34246 41550 34284 41553
rect 34336 41550 34495 41553
rect 34547 41550 34707 41553
rect 31328 41504 31349 41550
rect 33323 41504 33336 41550
rect 33671 41504 33684 41550
rect 33730 41504 33787 41550
rect 33833 41504 33890 41550
rect 33936 41504 33993 41550
rect 34039 41504 34096 41550
rect 34142 41504 34199 41550
rect 34245 41504 34284 41550
rect 34348 41504 34405 41550
rect 34451 41504 34495 41550
rect 34554 41504 34612 41550
rect 34658 41504 34707 41550
rect 31328 41501 31486 41504
rect 31538 41501 31697 41504
rect 31749 41501 31909 41504
rect 31961 41501 32120 41504
rect 32172 41501 32330 41504
rect 32382 41501 32541 41504
rect 32593 41501 32752 41504
rect 32804 41501 32842 41504
rect 30583 41466 32842 41501
rect 34246 41501 34284 41504
rect 34336 41501 34495 41504
rect 34547 41501 34707 41504
rect 34759 41501 34918 41553
rect 34970 41501 35008 41553
rect 34246 41467 35008 41501
rect 29544 41460 30306 41461
rect 27387 41344 29196 41420
rect 27387 41303 29116 41344
rect 27387 41257 28810 41303
rect 28856 41298 29116 41303
rect 29162 41298 29196 41344
rect 28856 41257 29196 41298
rect 27387 41181 29196 41257
rect 27387 41140 29116 41181
rect 27387 41094 28810 41140
rect 28856 41135 29116 41140
rect 29162 41135 29196 41181
rect 28856 41094 29196 41135
rect 27387 41017 29196 41094
rect 27387 40977 29116 41017
rect 27387 40931 28810 40977
rect 28856 40971 29116 40977
rect 29162 40971 29196 41017
rect 28856 40931 29196 40971
rect 27387 40854 29196 40931
rect 27387 40813 29116 40854
rect 27387 40767 28810 40813
rect 28856 40808 29116 40813
rect 29162 40808 29196 40854
rect 28856 40767 29196 40808
rect 27387 40653 29196 40767
rect 30583 41420 30637 41466
rect 30683 41460 32842 41466
rect 34247 41460 35008 41467
rect 35182 41587 36364 41594
rect 35182 41553 36958 41587
rect 35182 41501 35220 41553
rect 35272 41501 35430 41553
rect 35482 41501 35641 41553
rect 35693 41501 35853 41553
rect 35905 41501 36064 41553
rect 36116 41501 36274 41553
rect 36326 41550 36958 41553
rect 36326 41504 36489 41550
rect 36723 41504 36958 41550
rect 36326 41501 36958 41504
rect 35182 41467 36958 41501
rect 37946 41553 38842 41594
rect 37946 41550 38330 41553
rect 38382 41550 38541 41553
rect 37946 41504 37957 41550
rect 38473 41504 38541 41550
rect 37946 41501 38330 41504
rect 38382 41501 38541 41504
rect 38593 41501 38752 41553
rect 38804 41501 38842 41553
rect 35182 41460 36364 41467
rect 37946 41460 38842 41501
rect 39014 41553 39323 42039
rect 39014 41501 39052 41553
rect 39104 41550 39232 41553
rect 39108 41504 39220 41550
rect 39104 41501 39232 41504
rect 39284 41501 39323 41553
rect 30683 41426 31040 41460
rect 30683 41420 30855 41426
rect 30583 41380 30855 41420
rect 30901 41380 31040 41426
rect 30583 41303 31040 41380
rect 33484 41384 33552 41395
rect 33019 41329 33327 41370
rect 33019 41326 33057 41329
rect 33109 41326 33237 41329
rect 33289 41326 33327 41329
rect 30583 41257 30637 41303
rect 30683 41262 31040 41303
rect 31336 41280 31349 41326
rect 33323 41280 33336 41326
rect 30683 41257 30855 41262
rect 30583 41216 30855 41257
rect 30901 41216 31040 41262
rect 33019 41277 33057 41280
rect 33109 41277 33237 41280
rect 33289 41277 33327 41280
rect 33019 41237 33327 41277
rect 30583 41140 31040 41216
rect 30583 41094 30637 41140
rect 30683 41124 31040 41140
rect 30683 41102 31493 41124
rect 30683 41099 31349 41102
rect 30683 41094 30855 41099
rect 30583 41053 30855 41094
rect 30901 41056 31349 41099
rect 33323 41056 33336 41102
rect 30901 41053 31493 41056
rect 30583 41005 31493 41053
rect 30583 40977 31040 41005
rect 30583 40931 30637 40977
rect 30683 40936 31040 40977
rect 30683 40931 30855 40936
rect 30583 40890 30855 40931
rect 30901 40890 31040 40936
rect 33484 40962 33495 41384
rect 33541 40962 33552 41384
rect 33781 41337 34089 41378
rect 33781 41326 33819 41337
rect 33871 41326 33999 41337
rect 34051 41326 34089 41337
rect 33671 41280 33684 41326
rect 33730 41280 33787 41326
rect 33871 41285 33890 41326
rect 33833 41280 33890 41285
rect 33936 41280 33993 41326
rect 34051 41285 34096 41326
rect 34039 41280 34096 41285
rect 34142 41280 34199 41326
rect 34245 41280 34302 41326
rect 34348 41280 34405 41326
rect 34451 41280 34508 41326
rect 34554 41280 34612 41326
rect 34658 41280 34671 41326
rect 33781 41245 34089 41280
rect 35294 41251 36266 41291
rect 37853 41288 38161 41304
rect 35294 41239 35332 41251
rect 35384 41239 35543 41251
rect 35595 41239 35754 41251
rect 35806 41239 35965 41251
rect 36017 41239 36176 41251
rect 36228 41239 36266 41251
rect 36438 41239 36953 41288
rect 37439 41263 38161 41288
rect 37439 41239 37891 41263
rect 37943 41239 38071 41263
rect 38123 41239 38161 41263
rect 35260 41193 35273 41239
rect 35523 41199 35543 41239
rect 35523 41193 35580 41199
rect 35626 41193 35683 41239
rect 35729 41199 35754 41239
rect 35729 41193 35786 41199
rect 35832 41193 35889 41239
rect 35935 41199 35965 41239
rect 35935 41193 35992 41199
rect 36038 41193 36095 41239
rect 36141 41199 36176 41239
rect 36141 41193 36198 41199
rect 36244 41193 36301 41239
rect 36347 41193 36360 41239
rect 36438 41193 36854 41239
rect 36900 41193 36971 41239
rect 37017 41193 37088 41239
rect 37134 41193 37206 41239
rect 37252 41193 37324 41239
rect 37370 41193 37442 41239
rect 37488 41211 37891 41239
rect 37488 41193 37909 41211
rect 37955 41193 38026 41239
rect 38123 41211 38143 41239
rect 38072 41193 38143 41211
rect 38189 41193 38261 41239
rect 38307 41193 38379 41239
rect 38425 41193 38497 41239
rect 38543 41193 38556 41239
rect 35294 41159 36266 41193
rect 36438 41168 36953 41193
rect 37439 41171 38161 41193
rect 37439 41168 37931 41171
rect 34228 41102 34718 41131
rect 33671 41056 33684 41102
rect 33730 41056 33787 41102
rect 33833 41056 33890 41102
rect 33936 41056 33993 41102
rect 34039 41056 34096 41102
rect 34142 41056 34199 41102
rect 34245 41091 34302 41102
rect 34245 41056 34267 41091
rect 34348 41056 34405 41102
rect 34451 41091 34508 41102
rect 34499 41056 34508 41091
rect 34554 41056 34612 41102
rect 34658 41091 34718 41102
rect 34228 41039 34267 41056
rect 34319 41039 34447 41056
rect 34499 41039 34627 41056
rect 34679 41039 34718 41091
rect 36438 41065 36554 41168
rect 34228 40998 34718 41039
rect 34964 41015 36360 41059
rect 30583 40813 31040 40890
rect 33019 40881 33327 40922
rect 33019 40878 33057 40881
rect 33109 40878 33237 40881
rect 33289 40878 33327 40881
rect 33484 40880 33552 40962
rect 34964 40969 35273 41015
rect 35523 40969 35580 41015
rect 35626 40969 35683 41015
rect 35729 40969 35786 41015
rect 35832 40969 35889 41015
rect 35935 40969 35992 41015
rect 36038 40969 36095 41015
rect 36141 40969 36198 41015
rect 36244 40969 36301 41015
rect 36347 40969 36360 41015
rect 34964 40937 36360 40969
rect 34964 40880 35082 40937
rect 31336 40832 31349 40878
rect 33323 40832 33336 40878
rect 33484 40843 35082 40880
rect 30583 40767 30637 40813
rect 30683 40773 31040 40813
rect 33019 40829 33057 40832
rect 33109 40829 33237 40832
rect 33289 40829 33327 40832
rect 33019 40789 33327 40829
rect 33484 40797 33816 40843
rect 33862 40797 34002 40843
rect 34048 40797 34189 40843
rect 34235 40797 34376 40843
rect 34422 40797 34562 40843
rect 34608 40797 35082 40843
rect 36438 40925 36475 41065
rect 36521 40925 36554 41065
rect 33484 40789 35082 40797
rect 35294 40791 36266 40831
rect 36438 40825 36554 40925
rect 36640 41065 36773 41088
rect 36640 41016 36697 41065
rect 36640 40964 36678 41016
rect 36640 40925 36697 40964
rect 36743 40925 36773 41065
rect 38658 41067 38726 41078
rect 36924 41057 37685 41063
rect 36923 41056 37685 41057
rect 36923 41023 37931 41056
rect 36923 41015 36961 41023
rect 37013 41015 37172 41023
rect 37224 41015 37384 41023
rect 36841 40969 36854 41015
rect 36900 40971 36961 41015
rect 36900 40969 36971 40971
rect 37017 40969 37088 41015
rect 37134 40971 37172 41015
rect 37134 40969 37206 40971
rect 37252 40969 37324 41015
rect 37370 40971 37384 41015
rect 37436 41015 37595 41023
rect 37436 40971 37442 41015
rect 37370 40969 37442 40971
rect 37488 40971 37595 41015
rect 37647 41015 37931 41023
rect 37647 40971 37909 41015
rect 37488 40969 37909 40971
rect 37955 40969 38026 41015
rect 38072 40969 38143 41015
rect 38189 40969 38261 41015
rect 38307 40969 38379 41015
rect 38425 40969 38497 41015
rect 38543 40969 38556 41015
rect 36923 40937 37931 40969
rect 36924 40930 37685 40937
rect 36640 40905 36773 40925
rect 38658 40927 38669 41067
rect 38715 40927 38726 41067
rect 39014 41015 39323 41501
rect 39492 41587 39608 42039
rect 39923 42006 40085 42137
rect 39923 41954 39994 42006
rect 40046 41954 40085 42006
rect 39923 41914 40085 41954
rect 39737 41818 39865 41831
rect 39737 41791 39866 41818
rect 39737 41774 39775 41791
rect 39827 41774 39866 41791
rect 39727 41728 39740 41774
rect 39827 41739 39862 41774
rect 39786 41728 39862 41739
rect 39908 41728 39985 41774
rect 40031 41728 40108 41774
rect 40154 41728 40167 41774
rect 40246 41763 40362 42161
rect 42229 42022 44509 42063
rect 42229 41970 43445 42022
rect 43497 41970 44509 42022
rect 42229 41930 44509 41970
rect 44341 41886 44509 41930
rect 44341 41840 44358 41886
rect 44498 41840 44509 41886
rect 39737 41699 39866 41728
rect 40246 41717 40281 41763
rect 40327 41717 40362 41763
rect 40246 41680 40362 41717
rect 40718 41791 43524 41832
rect 44341 41829 44509 41840
rect 40718 41739 41935 41791
rect 41987 41739 43524 41791
rect 40718 41698 43524 41739
rect 44605 41774 44721 42161
rect 45400 42131 48379 42172
rect 45400 42117 45975 42131
rect 45400 42071 45464 42117
rect 45604 42079 45975 42117
rect 46027 42079 48379 42131
rect 45604 42071 48379 42079
rect 44901 42015 45241 42056
rect 45400 42038 48379 42071
rect 48557 42125 48596 42177
rect 48648 42125 48687 42177
rect 48557 42102 48687 42125
rect 50044 42211 50516 42257
rect 50562 42211 50703 42257
rect 50749 42211 50890 42257
rect 50936 42211 51076 42257
rect 51122 42211 51263 42257
rect 51309 42211 51657 42257
rect 51797 42247 52105 42287
rect 51797 42222 51835 42247
rect 51887 42222 52015 42247
rect 52067 42222 52105 42247
rect 54085 42281 54223 42327
rect 54269 42287 54540 42327
rect 54269 42281 54440 42287
rect 54085 42241 54440 42281
rect 54486 42241 54540 42287
rect 50044 42174 51657 42211
rect 51789 42176 51802 42222
rect 53776 42176 53789 42222
rect 50044 42117 50160 42174
rect 44901 41998 44939 42015
rect 44991 41998 45151 42015
rect 45203 41998 45241 42015
rect 44799 41952 44812 41998
rect 44858 41952 44925 41998
rect 44991 41963 45038 41998
rect 44971 41952 45038 41963
rect 45084 41952 45151 41998
rect 45203 41963 45264 41998
rect 45197 41952 45264 41963
rect 45310 41952 45323 41998
rect 48557 41962 48622 42102
rect 48668 41962 48687 42102
rect 49820 42085 50160 42117
rect 48765 42039 48778 42085
rect 48824 42039 48881 42085
rect 48927 42039 48984 42085
rect 49030 42039 49087 42085
rect 49133 42039 49190 42085
rect 49236 42039 49293 42085
rect 49339 42039 49396 42085
rect 49442 42039 49499 42085
rect 49545 42039 49602 42085
rect 49852 42039 50160 42085
rect 51589 42122 51657 42174
rect 51797 42154 52105 42176
rect 49820 41998 50160 42039
rect 50262 42015 50812 42056
rect 48557 41959 48687 41962
rect 44901 41923 45241 41952
rect 48557 41907 48596 41959
rect 48648 41907 48687 41959
rect 50262 41963 50300 42015
rect 50352 41998 50511 42015
rect 50563 41998 50722 42015
rect 50352 41963 50467 41998
rect 50563 41963 50571 41998
rect 50262 41952 50467 41963
rect 50513 41952 50571 41963
rect 50617 41952 50674 41998
rect 50720 41963 50722 41998
rect 50774 41998 50812 42015
rect 50774 41963 50777 41998
rect 50720 41952 50777 41963
rect 50823 41952 50880 41998
rect 50926 41952 50983 41998
rect 51029 41952 51086 41998
rect 51132 41952 51189 41998
rect 51235 41952 51292 41998
rect 51338 41952 51395 41998
rect 51441 41952 51454 41998
rect 50262 41923 50812 41952
rect 48557 41866 48687 41907
rect 48905 41861 49877 41892
rect 48765 41815 48778 41861
rect 48824 41815 48881 41861
rect 48927 41852 48984 41861
rect 48927 41815 48943 41852
rect 49030 41815 49087 41861
rect 49133 41852 49190 41861
rect 49133 41815 49154 41852
rect 49236 41815 49293 41861
rect 49339 41852 49396 41861
rect 49339 41815 49365 41852
rect 49442 41815 49499 41861
rect 49545 41852 49602 41861
rect 49545 41815 49576 41852
rect 49852 41815 49877 41861
rect 48905 41800 48943 41815
rect 48995 41800 49154 41815
rect 49206 41800 49365 41815
rect 49417 41800 49576 41815
rect 49628 41800 49787 41815
rect 49839 41800 49877 41815
rect 44605 41728 44812 41774
rect 44858 41728 44925 41774
rect 44971 41728 45038 41774
rect 45084 41728 45151 41774
rect 45197 41728 45264 41774
rect 45310 41728 45323 41774
rect 48905 41760 49877 41800
rect 51035 41777 51343 41817
rect 51035 41774 51073 41777
rect 51125 41774 51253 41777
rect 51305 41774 51343 41777
rect 43362 41691 43524 41698
rect 43362 41645 43373 41691
rect 43513 41645 43524 41691
rect 43362 41634 43524 41645
rect 45584 41714 48546 41750
rect 50454 41728 50467 41774
rect 50513 41728 50571 41774
rect 50617 41728 50674 41774
rect 50720 41728 50777 41774
rect 50823 41728 50880 41774
rect 50926 41728 50983 41774
rect 51029 41728 51073 41774
rect 51132 41728 51189 41774
rect 51235 41728 51253 41774
rect 51338 41728 51395 41774
rect 51441 41728 51454 41774
rect 45584 41668 45619 41714
rect 45665 41668 45777 41714
rect 45823 41668 45935 41714
rect 45981 41668 46093 41714
rect 46139 41668 46251 41714
rect 46297 41668 46409 41714
rect 46455 41668 46568 41714
rect 46614 41668 46726 41714
rect 46772 41668 46884 41714
rect 46930 41668 47042 41714
rect 47088 41668 47200 41714
rect 47246 41668 47358 41714
rect 47404 41668 47516 41714
rect 47562 41668 47675 41714
rect 47721 41668 47833 41714
rect 47879 41668 47991 41714
rect 48037 41668 48149 41714
rect 48195 41668 48307 41714
rect 48353 41668 48465 41714
rect 48511 41668 48546 41714
rect 51035 41725 51073 41728
rect 51125 41725 51253 41728
rect 51305 41725 51343 41728
rect 51035 41684 51343 41725
rect 51589 41700 51600 42122
rect 51646 41700 51657 42122
rect 54085 42123 54540 42241
rect 54085 42077 54440 42123
rect 54486 42077 54540 42123
rect 54085 42049 54540 42077
rect 53585 41998 54540 42049
rect 51789 41952 51802 41998
rect 53776 41960 54540 41998
rect 53776 41952 54440 41960
rect 53585 41930 54440 41952
rect 54085 41914 54440 41930
rect 54486 41914 54540 41960
rect 54085 41838 54540 41914
rect 51797 41784 52105 41824
rect 51797 41774 51835 41784
rect 51887 41774 52015 41784
rect 52067 41774 52105 41784
rect 54085 41792 54223 41838
rect 54269 41797 54540 41838
rect 54269 41792 54440 41797
rect 51789 41728 51802 41774
rect 53776 41728 53789 41774
rect 54085 41751 54440 41792
rect 54486 41751 54540 41797
rect 51589 41689 51657 41700
rect 51797 41691 52105 41728
rect 40215 41587 40523 41594
rect 40788 41587 42986 41601
rect 43753 41587 44514 41594
rect 39492 41564 42986 41587
rect 43704 41564 44514 41587
rect 39492 41553 44514 41564
rect 39492 41550 40253 41553
rect 39492 41504 39740 41550
rect 39786 41504 39862 41550
rect 39908 41504 39985 41550
rect 40031 41504 40108 41550
rect 40154 41504 40253 41550
rect 39492 41501 40253 41504
rect 40305 41501 40433 41553
rect 40485 41550 43790 41553
rect 40485 41504 40836 41550
rect 40882 41504 40994 41550
rect 41040 41504 41152 41550
rect 41198 41504 41310 41550
rect 41356 41504 41469 41550
rect 41515 41504 41627 41550
rect 41673 41504 41785 41550
rect 41831 41504 41943 41550
rect 41989 41504 42101 41550
rect 42147 41504 42259 41550
rect 42305 41504 42418 41550
rect 42464 41504 42576 41550
rect 42622 41504 42734 41550
rect 42780 41504 42892 41550
rect 42938 41504 43739 41550
rect 43785 41504 43790 41550
rect 40485 41501 43790 41504
rect 43842 41550 44001 41553
rect 43842 41504 43906 41550
rect 43952 41504 44001 41550
rect 43842 41501 44001 41504
rect 44053 41550 44213 41553
rect 44265 41550 44424 41553
rect 44053 41504 44071 41550
rect 44117 41504 44213 41550
rect 44282 41504 44424 41550
rect 44053 41501 44213 41504
rect 44265 41501 44424 41504
rect 44476 41501 44514 41553
rect 39492 41490 44514 41501
rect 39492 41467 42986 41490
rect 43704 41467 44514 41490
rect 39492 41015 39608 41467
rect 40215 41460 40523 41467
rect 40788 41453 42986 41467
rect 43753 41460 44514 41467
rect 44796 41587 45346 41594
rect 45584 41587 48546 41668
rect 54085 41674 54540 41751
rect 54085 41628 54223 41674
rect 54269 41634 54540 41674
rect 54269 41628 54440 41634
rect 54085 41594 54440 41628
rect 48800 41587 49982 41594
rect 50308 41587 50859 41594
rect 44796 41553 49982 41587
rect 44796 41550 44834 41553
rect 44886 41550 45045 41553
rect 45097 41550 45256 41553
rect 45308 41550 48838 41553
rect 44796 41504 44812 41550
rect 44886 41504 44925 41550
rect 44971 41504 45038 41550
rect 45097 41504 45151 41550
rect 45197 41504 45256 41550
rect 45310 41504 45619 41550
rect 45665 41504 45777 41550
rect 45823 41504 45935 41550
rect 45981 41504 46093 41550
rect 46139 41504 46251 41550
rect 46297 41504 46409 41550
rect 46455 41504 46568 41550
rect 46614 41504 46726 41550
rect 46772 41504 46884 41550
rect 46930 41504 47042 41550
rect 47088 41504 47200 41550
rect 47246 41504 47358 41550
rect 47404 41504 47516 41550
rect 47562 41504 47675 41550
rect 47721 41504 47833 41550
rect 47879 41504 47991 41550
rect 48037 41504 48149 41550
rect 48195 41504 48307 41550
rect 48353 41504 48465 41550
rect 48511 41504 48838 41550
rect 44796 41501 44834 41504
rect 44886 41501 45045 41504
rect 45097 41501 45256 41504
rect 45308 41501 48838 41504
rect 48890 41501 49048 41553
rect 49100 41501 49259 41553
rect 49311 41501 49471 41553
rect 49523 41501 49682 41553
rect 49734 41501 49892 41553
rect 49944 41501 49982 41553
rect 44796 41467 49982 41501
rect 50307 41553 50859 41587
rect 50307 41501 50346 41553
rect 50398 41550 50557 41553
rect 50609 41550 50768 41553
rect 50820 41550 50859 41553
rect 52278 41588 54440 41594
rect 54486 41588 54540 41634
rect 55927 42287 57736 42401
rect 55927 42244 56267 42287
rect 55927 42198 55961 42244
rect 56007 42241 56267 42244
rect 56313 42241 57736 42287
rect 56007 42198 57736 42241
rect 55927 42123 57736 42198
rect 55927 42081 56267 42123
rect 55927 42035 55961 42081
rect 56007 42077 56267 42081
rect 56313 42077 57736 42123
rect 56007 42035 57736 42077
rect 55927 41960 57736 42035
rect 55927 41917 56267 41960
rect 55927 41871 55961 41917
rect 56007 41914 56267 41917
rect 56313 41914 57736 41960
rect 56007 41871 57736 41914
rect 55927 41797 57736 41871
rect 55927 41754 56267 41797
rect 55927 41708 55961 41754
rect 56007 41751 56267 41754
rect 56313 41751 57736 41797
rect 56007 41708 57736 41751
rect 55927 41634 57736 41708
rect 52278 41553 54540 41588
rect 52278 41550 52316 41553
rect 52368 41550 52527 41553
rect 52579 41550 52738 41553
rect 52790 41550 52948 41553
rect 53000 41550 53159 41553
rect 53211 41550 53371 41553
rect 53423 41550 53582 41553
rect 53634 41550 53792 41553
rect 50398 41504 50467 41550
rect 50513 41504 50557 41550
rect 50617 41504 50674 41550
rect 50720 41504 50768 41550
rect 50823 41504 50880 41550
rect 50926 41504 50983 41550
rect 51029 41504 51086 41550
rect 51132 41504 51189 41550
rect 51235 41504 51292 41550
rect 51338 41504 51395 41550
rect 51441 41504 51454 41550
rect 51789 41504 51802 41550
rect 53776 41504 53792 41550
rect 50398 41501 50557 41504
rect 50609 41501 50768 41504
rect 50820 41501 50859 41504
rect 50307 41467 50859 41501
rect 44796 41460 45346 41467
rect 43362 41409 43524 41420
rect 39737 41326 39866 41355
rect 40246 41337 40362 41374
rect 43362 41363 43373 41409
rect 43513 41363 43524 41409
rect 43362 41356 43524 41363
rect 39727 41280 39740 41326
rect 39786 41315 39862 41326
rect 39827 41280 39862 41315
rect 39908 41280 39985 41326
rect 40031 41280 40108 41326
rect 40154 41280 40167 41326
rect 40246 41291 40281 41337
rect 40327 41291 40362 41337
rect 39737 41263 39775 41280
rect 39827 41263 39866 41280
rect 39737 41236 39866 41263
rect 39737 41223 39865 41236
rect 39923 41100 40085 41140
rect 39923 41048 39994 41100
rect 40046 41048 40085 41100
rect 39008 40969 39021 41015
rect 39067 40969 39144 41015
rect 39190 40969 39267 41015
rect 39313 40969 39326 41015
rect 39492 40969 39641 41015
rect 39687 40969 39730 41015
rect 39014 40937 39323 40969
rect 39492 40937 39608 40969
rect 37853 40825 38161 40830
rect 36438 40791 36953 40825
rect 37439 40791 38161 40825
rect 38658 40805 38726 40927
rect 39923 40917 40085 41048
rect 39809 40914 40085 40917
rect 39809 40906 39994 40914
rect 39809 40860 39844 40906
rect 39890 40862 39994 40906
rect 40046 40893 40085 40914
rect 40246 40893 40362 41291
rect 40718 41315 43524 41356
rect 45584 41386 48546 41467
rect 48800 41460 49982 41467
rect 50308 41460 50859 41467
rect 52278 41501 52316 41504
rect 52368 41501 52527 41504
rect 52579 41501 52738 41504
rect 52790 41501 52948 41504
rect 53000 41501 53159 41504
rect 53211 41501 53371 41504
rect 53423 41501 53582 41504
rect 53634 41501 53792 41504
rect 53844 41501 54003 41553
rect 54055 41501 54214 41553
rect 54266 41501 54540 41553
rect 52278 41466 54540 41501
rect 52278 41460 54440 41466
rect 45584 41340 45619 41386
rect 45665 41340 45777 41386
rect 45823 41340 45935 41386
rect 45981 41340 46093 41386
rect 46139 41340 46251 41386
rect 46297 41340 46409 41386
rect 46455 41340 46568 41386
rect 46614 41340 46726 41386
rect 46772 41340 46884 41386
rect 46930 41340 47042 41386
rect 47088 41340 47200 41386
rect 47246 41340 47358 41386
rect 47404 41340 47516 41386
rect 47562 41340 47675 41386
rect 47721 41340 47833 41386
rect 47879 41340 47991 41386
rect 48037 41340 48149 41386
rect 48195 41340 48307 41386
rect 48353 41340 48465 41386
rect 48511 41340 48546 41386
rect 54085 41426 54440 41460
rect 54085 41380 54223 41426
rect 54269 41420 54440 41426
rect 54486 41420 54540 41466
rect 54758 41553 55840 41594
rect 54758 41550 54855 41553
rect 54758 41504 54793 41550
rect 54839 41504 54855 41550
rect 54758 41501 54855 41504
rect 54907 41550 55066 41553
rect 54907 41504 54956 41550
rect 55002 41504 55066 41550
rect 54907 41501 55066 41504
rect 55118 41550 55278 41553
rect 55330 41550 55489 41553
rect 55164 41504 55278 41550
rect 55330 41504 55439 41550
rect 55485 41504 55489 41550
rect 55118 41501 55278 41504
rect 55330 41501 55489 41504
rect 55541 41550 55840 41553
rect 55541 41504 55599 41550
rect 55645 41504 55760 41550
rect 55806 41504 55840 41550
rect 55541 41501 55840 41504
rect 54758 41461 55840 41501
rect 55927 41588 56267 41634
rect 56313 41588 57736 41634
rect 55927 41466 57736 41588
rect 54817 41460 55579 41461
rect 54269 41380 54540 41420
rect 40718 41263 41935 41315
rect 41987 41263 43524 41315
rect 40718 41222 43524 41263
rect 44605 41280 44812 41326
rect 44858 41280 44925 41326
rect 44971 41280 45038 41326
rect 45084 41280 45151 41326
rect 45197 41280 45264 41326
rect 45310 41280 45323 41326
rect 45584 41304 48546 41340
rect 51035 41329 51343 41370
rect 51035 41326 51073 41329
rect 51125 41326 51253 41329
rect 51305 41326 51343 41329
rect 51589 41354 51657 41365
rect 44341 41214 44509 41225
rect 44341 41168 44358 41214
rect 44498 41168 44509 41214
rect 44341 41124 44509 41168
rect 42229 41084 44509 41124
rect 42229 41032 43445 41084
rect 43497 41032 44509 41084
rect 42229 40991 44509 41032
rect 44605 40893 44721 41280
rect 48905 41254 49877 41294
rect 50454 41280 50467 41326
rect 50513 41280 50571 41326
rect 50617 41280 50674 41326
rect 50720 41280 50777 41326
rect 50823 41280 50880 41326
rect 50926 41280 50983 41326
rect 51029 41280 51073 41326
rect 51132 41280 51189 41326
rect 51235 41280 51253 41326
rect 51338 41280 51395 41326
rect 51441 41280 51454 41326
rect 48905 41239 48943 41254
rect 48995 41239 49154 41254
rect 49206 41239 49365 41254
rect 49417 41239 49576 41254
rect 49628 41239 49787 41254
rect 49839 41239 49877 41254
rect 48765 41193 48778 41239
rect 48824 41193 48881 41239
rect 48927 41202 48943 41239
rect 48927 41193 48984 41202
rect 49030 41193 49087 41239
rect 49133 41202 49154 41239
rect 49133 41193 49190 41202
rect 49236 41193 49293 41239
rect 49339 41202 49365 41239
rect 49339 41193 49396 41202
rect 49442 41193 49499 41239
rect 49545 41202 49576 41239
rect 49545 41193 49602 41202
rect 49852 41193 49877 41239
rect 51035 41277 51073 41280
rect 51125 41277 51253 41280
rect 51305 41277 51343 41280
rect 51035 41237 51343 41277
rect 48557 41147 48687 41188
rect 48905 41162 49877 41193
rect 44901 41102 45241 41131
rect 44799 41056 44812 41102
rect 44858 41056 44925 41102
rect 44971 41091 45038 41102
rect 44991 41056 45038 41091
rect 45084 41056 45151 41102
rect 45197 41091 45264 41102
rect 45203 41056 45264 41091
rect 45310 41056 45323 41102
rect 48557 41095 48596 41147
rect 48648 41095 48687 41147
rect 48557 41092 48687 41095
rect 44901 41039 44939 41056
rect 44991 41039 45151 41056
rect 45203 41039 45241 41056
rect 44901 40998 45241 41039
rect 45400 40983 48379 41016
rect 45400 40937 45464 40983
rect 45604 40975 48379 40983
rect 45604 40937 46353 40975
rect 45400 40923 46353 40937
rect 46405 40923 48379 40975
rect 40046 40878 44918 40893
rect 45400 40882 48379 40923
rect 48557 40952 48622 41092
rect 48668 40952 48687 41092
rect 50262 41102 50812 41131
rect 50262 41091 50467 41102
rect 50513 41091 50571 41102
rect 49820 41015 50160 41056
rect 48765 40969 48778 41015
rect 48824 40969 48881 41015
rect 48927 40969 48984 41015
rect 49030 40969 49087 41015
rect 49133 40969 49190 41015
rect 49236 40969 49293 41015
rect 49339 40969 49396 41015
rect 49442 40969 49499 41015
rect 49545 40969 49602 41015
rect 49852 40969 50160 41015
rect 50262 41039 50300 41091
rect 50352 41056 50467 41091
rect 50563 41056 50571 41091
rect 50617 41056 50674 41102
rect 50720 41091 50777 41102
rect 50720 41056 50722 41091
rect 50352 41039 50511 41056
rect 50563 41039 50722 41056
rect 50774 41056 50777 41091
rect 50823 41056 50880 41102
rect 50926 41056 50983 41102
rect 51029 41056 51086 41102
rect 51132 41056 51189 41102
rect 51235 41056 51292 41102
rect 51338 41056 51395 41102
rect 51441 41056 51454 41102
rect 50774 41039 50812 41056
rect 50262 40998 50812 41039
rect 48557 40929 48687 40952
rect 49820 40937 50160 40969
rect 40046 40862 44812 40878
rect 39890 40860 44812 40862
rect 39809 40857 44812 40860
rect 39809 40811 43739 40857
rect 43785 40811 43906 40857
rect 43952 40811 44071 40857
rect 44117 40811 44236 40857
rect 44282 40832 44812 40857
rect 44858 40832 44925 40878
rect 44971 40832 45038 40878
rect 45084 40832 45151 40878
rect 45197 40832 45264 40878
rect 45310 40832 45323 40878
rect 48557 40877 48596 40929
rect 48648 40877 48687 40929
rect 48557 40837 48687 40877
rect 50044 40880 50160 40937
rect 51589 40932 51600 41354
rect 51646 40932 51657 41354
rect 51797 41326 52105 41363
rect 51789 41280 51802 41326
rect 53776 41280 53789 41326
rect 54085 41303 54540 41380
rect 51797 41270 51835 41280
rect 51887 41270 52015 41280
rect 52067 41270 52105 41280
rect 51797 41230 52105 41270
rect 54085 41262 54440 41303
rect 54085 41216 54223 41262
rect 54269 41257 54440 41262
rect 54486 41257 54540 41303
rect 54269 41216 54540 41257
rect 54085 41140 54540 41216
rect 54085 41124 54440 41140
rect 53585 41102 54440 41124
rect 51789 41056 51802 41102
rect 53776 41094 54440 41102
rect 54486 41094 54540 41140
rect 53776 41056 54540 41094
rect 53585 41005 54540 41056
rect 51589 40880 51657 40932
rect 54085 40977 54540 41005
rect 54085 40931 54440 40977
rect 54486 40931 54540 40977
rect 50044 40843 51657 40880
rect 51797 40878 52105 40900
rect 44282 40811 44918 40832
rect 38658 40791 39723 40805
rect 30683 40767 30855 40773
rect 30583 40727 30855 40767
rect 30901 40727 31040 40773
rect 33484 40760 34643 40789
rect 35260 40745 35273 40791
rect 35523 40745 35543 40791
rect 35626 40745 35683 40791
rect 35729 40745 35754 40791
rect 35832 40745 35889 40791
rect 35935 40745 35965 40791
rect 36038 40745 36095 40791
rect 36141 40745 36176 40791
rect 36244 40745 36301 40791
rect 36347 40745 36360 40791
rect 36438 40745 36854 40791
rect 36900 40745 36971 40791
rect 37017 40745 37088 40791
rect 37134 40745 37206 40791
rect 37252 40745 37324 40791
rect 37370 40745 37442 40791
rect 37488 40789 37909 40791
rect 37488 40745 37891 40789
rect 37955 40745 38026 40791
rect 38072 40789 38143 40791
rect 38123 40745 38143 40789
rect 38189 40745 38261 40791
rect 38307 40745 38379 40791
rect 38425 40745 38497 40791
rect 38543 40745 38556 40791
rect 38658 40745 39021 40791
rect 39067 40745 39144 40791
rect 39190 40745 39267 40791
rect 39313 40745 39641 40791
rect 39687 40745 39730 40791
rect 39809 40773 44918 40811
rect 48905 40791 49877 40831
rect 48765 40745 48778 40791
rect 48824 40745 48881 40791
rect 48927 40745 48943 40791
rect 49030 40745 49087 40791
rect 49133 40745 49154 40791
rect 49236 40745 49293 40791
rect 49339 40745 49365 40791
rect 49442 40745 49499 40791
rect 49545 40745 49576 40791
rect 49852 40745 49877 40791
rect 50044 40797 50516 40843
rect 50562 40797 50703 40843
rect 50749 40797 50890 40843
rect 50936 40797 51076 40843
rect 51122 40797 51263 40843
rect 51309 40797 51657 40843
rect 51789 40832 51802 40878
rect 53776 40832 53789 40878
rect 50044 40787 51657 40797
rect 50481 40760 51657 40787
rect 51797 40807 51835 40832
rect 51887 40807 52015 40832
rect 52067 40807 52105 40832
rect 51797 40767 52105 40807
rect 54085 40813 54540 40931
rect 54085 40773 54440 40813
rect 30583 40694 31040 40727
rect 35294 40739 35332 40745
rect 35384 40739 35543 40745
rect 35595 40739 35754 40745
rect 35806 40739 35965 40745
rect 36017 40739 36176 40745
rect 36228 40739 36266 40745
rect 34870 40694 35025 40701
rect 35294 40699 36266 40739
rect 36438 40705 36953 40745
rect 37439 40737 37891 40745
rect 37943 40737 38071 40745
rect 38123 40737 38161 40745
rect 37439 40705 38161 40737
rect 37853 40697 38161 40705
rect 27387 40601 27790 40653
rect 27842 40601 28001 40653
rect 28053 40601 28212 40653
rect 28264 40601 28423 40653
rect 28475 40601 28634 40653
rect 28686 40650 28845 40653
rect 28686 40604 28810 40650
rect 28686 40601 28845 40604
rect 28897 40601 29056 40653
rect 29108 40601 29196 40653
rect 27387 40487 29196 40601
rect 29283 40653 30365 40694
rect 29283 40650 29582 40653
rect 29283 40604 29317 40650
rect 29363 40604 29478 40650
rect 29524 40604 29582 40650
rect 29283 40601 29582 40604
rect 29634 40650 29793 40653
rect 29845 40650 30005 40653
rect 29634 40604 29638 40650
rect 29684 40604 29793 40650
rect 29845 40604 29959 40650
rect 29634 40601 29793 40604
rect 29845 40601 30005 40604
rect 30057 40650 30216 40653
rect 30057 40604 30121 40650
rect 30167 40604 30216 40650
rect 30057 40601 30216 40604
rect 30268 40650 30365 40653
rect 30268 40604 30284 40650
rect 30330 40604 30365 40650
rect 30268 40601 30365 40604
rect 29283 40561 30365 40601
rect 30583 40653 32842 40694
rect 30583 40650 30854 40653
rect 30583 40604 30637 40650
rect 30683 40604 30854 40650
rect 30583 40601 30854 40604
rect 30906 40601 31065 40653
rect 31117 40601 31276 40653
rect 31328 40601 31486 40653
rect 31538 40601 31697 40653
rect 31749 40601 31909 40653
rect 31961 40601 32120 40653
rect 32172 40601 32330 40653
rect 32382 40601 32541 40653
rect 32593 40601 32752 40653
rect 32804 40601 32842 40653
rect 29544 40560 30306 40561
rect 30583 40560 32842 40601
rect 34717 40653 35025 40694
rect 38658 40685 39723 40745
rect 48905 40739 48943 40745
rect 48995 40739 49154 40745
rect 49206 40739 49365 40745
rect 49417 40739 49576 40745
rect 49628 40739 49787 40745
rect 49839 40739 49877 40745
rect 48905 40699 49877 40739
rect 54085 40727 54223 40773
rect 54269 40767 54440 40773
rect 54486 40767 54540 40813
rect 54269 40727 54540 40767
rect 50099 40694 50255 40701
rect 54085 40694 54540 40727
rect 55927 41420 56267 41466
rect 56313 41420 57736 41466
rect 55927 41344 57736 41420
rect 55927 41298 55961 41344
rect 56007 41303 57736 41344
rect 56007 41298 56267 41303
rect 55927 41257 56267 41298
rect 56313 41257 57736 41303
rect 55927 41181 57736 41257
rect 55927 41135 55961 41181
rect 56007 41140 57736 41181
rect 56007 41135 56267 41140
rect 55927 41094 56267 41135
rect 56313 41094 57736 41140
rect 55927 41017 57736 41094
rect 55927 40971 55961 41017
rect 56007 40977 57736 41017
rect 56007 40971 56267 40977
rect 55927 40931 56267 40971
rect 56313 40931 57736 40977
rect 55927 40854 57736 40931
rect 55927 40808 55961 40854
rect 56007 40813 57736 40854
rect 56007 40808 56267 40813
rect 55927 40767 56267 40808
rect 56313 40767 57736 40813
rect 34717 40601 34755 40653
rect 34807 40650 34935 40653
rect 34807 40604 34916 40650
rect 34807 40601 34935 40604
rect 34987 40601 35025 40653
rect 34717 40560 35025 40601
rect 50099 40653 50408 40694
rect 50099 40601 50138 40653
rect 50190 40650 50318 40653
rect 50206 40604 50318 40650
rect 50190 40601 50318 40604
rect 50370 40601 50408 40653
rect 27387 40441 28810 40487
rect 28856 40444 29196 40487
rect 28856 40441 29116 40444
rect 27387 40398 29116 40441
rect 29162 40398 29196 40444
rect 27387 40323 29196 40398
rect 27387 40277 28810 40323
rect 28856 40281 29196 40323
rect 28856 40277 29116 40281
rect 27387 40235 29116 40277
rect 29162 40235 29196 40281
rect 27387 40160 29196 40235
rect 27387 40114 28810 40160
rect 28856 40117 29196 40160
rect 28856 40114 29116 40117
rect 27387 40071 29116 40114
rect 29162 40071 29196 40117
rect 27387 39997 29196 40071
rect 27387 39951 28810 39997
rect 28856 39954 29196 39997
rect 28856 39951 29116 39954
rect 27387 39908 29116 39951
rect 29162 39908 29196 39954
rect 27387 39834 29196 39908
rect 27387 39788 28810 39834
rect 28856 39788 29196 39834
rect 30583 40527 31040 40560
rect 34870 40553 35025 40560
rect 30583 40487 30855 40527
rect 30583 40441 30637 40487
rect 30683 40481 30855 40487
rect 30901 40481 31040 40527
rect 35294 40515 36266 40555
rect 37853 40549 38161 40557
rect 35294 40509 35332 40515
rect 35384 40509 35543 40515
rect 35595 40509 35754 40515
rect 35806 40509 35965 40515
rect 36017 40509 36176 40515
rect 36228 40509 36266 40515
rect 36438 40509 36953 40549
rect 37439 40517 38161 40549
rect 37439 40509 37891 40517
rect 37943 40509 38071 40517
rect 38123 40509 38161 40517
rect 38658 40509 39723 40569
rect 50099 40560 50408 40601
rect 52278 40653 54540 40694
rect 52278 40601 52316 40653
rect 52368 40601 52527 40653
rect 52579 40601 52738 40653
rect 52790 40601 52948 40653
rect 53000 40601 53159 40653
rect 53211 40601 53371 40653
rect 53423 40601 53582 40653
rect 53634 40601 53792 40653
rect 53844 40601 54003 40653
rect 54055 40601 54214 40653
rect 54266 40650 54540 40653
rect 54266 40604 54440 40650
rect 54486 40604 54540 40650
rect 54266 40601 54540 40604
rect 52278 40560 54540 40601
rect 54758 40653 55840 40694
rect 54758 40650 54855 40653
rect 54758 40604 54793 40650
rect 54839 40604 54855 40650
rect 54758 40601 54855 40604
rect 54907 40650 55066 40653
rect 54907 40604 54956 40650
rect 55002 40604 55066 40650
rect 54907 40601 55066 40604
rect 55118 40650 55278 40653
rect 55330 40650 55489 40653
rect 55164 40604 55278 40650
rect 55330 40604 55439 40650
rect 55485 40604 55489 40650
rect 55118 40601 55278 40604
rect 55330 40601 55489 40604
rect 55541 40650 55840 40653
rect 55541 40604 55599 40650
rect 55645 40604 55760 40650
rect 55806 40604 55840 40650
rect 55541 40601 55840 40604
rect 54758 40561 55840 40601
rect 55927 40653 57736 40767
rect 55927 40601 56015 40653
rect 56067 40601 56226 40653
rect 56278 40650 56437 40653
rect 56313 40604 56437 40650
rect 56278 40601 56437 40604
rect 56489 40601 56648 40653
rect 56700 40601 56859 40653
rect 56911 40601 57070 40653
rect 57122 40601 57281 40653
rect 57333 40601 57736 40653
rect 54817 40560 55579 40561
rect 48905 40515 49877 40555
rect 50099 40553 50255 40560
rect 48905 40509 48943 40515
rect 48995 40509 49154 40515
rect 49206 40509 49365 40515
rect 49417 40509 49576 40515
rect 49628 40509 49787 40515
rect 49839 40509 49877 40515
rect 30683 40441 31040 40481
rect 33484 40465 34643 40494
rect 30583 40364 31040 40441
rect 33019 40425 33327 40465
rect 33019 40422 33057 40425
rect 33109 40422 33237 40425
rect 33289 40422 33327 40425
rect 33484 40457 35082 40465
rect 35260 40463 35273 40509
rect 35523 40463 35543 40509
rect 35626 40463 35683 40509
rect 35729 40463 35754 40509
rect 35832 40463 35889 40509
rect 35935 40463 35965 40509
rect 36038 40463 36095 40509
rect 36141 40463 36176 40509
rect 36244 40463 36301 40509
rect 36347 40463 36360 40509
rect 36438 40463 36854 40509
rect 36900 40463 36971 40509
rect 37017 40463 37088 40509
rect 37134 40463 37206 40509
rect 37252 40463 37324 40509
rect 37370 40463 37442 40509
rect 37488 40465 37891 40509
rect 37488 40463 37909 40465
rect 37955 40463 38026 40509
rect 38123 40465 38143 40509
rect 38072 40463 38143 40465
rect 38189 40463 38261 40509
rect 38307 40463 38379 40509
rect 38425 40463 38497 40509
rect 38543 40463 38556 40509
rect 38658 40463 39021 40509
rect 39067 40463 39144 40509
rect 39190 40463 39267 40509
rect 39313 40463 39641 40509
rect 39687 40463 39730 40509
rect 31336 40376 31349 40422
rect 33323 40376 33336 40422
rect 33484 40411 33816 40457
rect 33862 40411 34002 40457
rect 34048 40411 34189 40457
rect 34235 40411 34376 40457
rect 34422 40411 34562 40457
rect 34608 40411 35082 40457
rect 35294 40423 36266 40463
rect 36438 40429 36953 40463
rect 37439 40429 38161 40463
rect 30583 40323 30855 40364
rect 30583 40277 30637 40323
rect 30683 40318 30855 40323
rect 30901 40318 31040 40364
rect 33019 40373 33057 40376
rect 33109 40373 33237 40376
rect 33289 40373 33327 40376
rect 33019 40332 33327 40373
rect 33484 40374 35082 40411
rect 30683 40277 31040 40318
rect 30583 40249 31040 40277
rect 33484 40292 33552 40374
rect 30583 40201 31493 40249
rect 30583 40160 30855 40201
rect 30583 40114 30637 40160
rect 30683 40155 30855 40160
rect 30901 40198 31493 40201
rect 30901 40155 31349 40198
rect 30683 40152 31349 40155
rect 33323 40152 33336 40198
rect 30683 40130 31493 40152
rect 30683 40114 31040 40130
rect 30583 40038 31040 40114
rect 30583 39997 30855 40038
rect 30583 39951 30637 39997
rect 30683 39992 30855 39997
rect 30901 39992 31040 40038
rect 30683 39951 31040 39992
rect 33019 39977 33327 40017
rect 33019 39974 33057 39977
rect 33109 39974 33237 39977
rect 33289 39974 33327 39977
rect 30583 39874 31040 39951
rect 31336 39928 31349 39974
rect 33323 39928 33336 39974
rect 33019 39925 33057 39928
rect 33109 39925 33237 39928
rect 33289 39925 33327 39928
rect 33019 39884 33327 39925
rect 30583 39834 30855 39874
rect 27387 39666 29196 39788
rect 27387 39620 28810 39666
rect 28856 39620 29196 39666
rect 29283 39753 30365 39794
rect 29283 39750 29582 39753
rect 29283 39704 29317 39750
rect 29363 39704 29478 39750
rect 29524 39704 29582 39750
rect 29283 39701 29582 39704
rect 29634 39750 29793 39753
rect 29845 39750 30005 39753
rect 29634 39704 29638 39750
rect 29684 39704 29793 39750
rect 29845 39704 29959 39750
rect 29634 39701 29793 39704
rect 29845 39701 30005 39704
rect 30057 39750 30216 39753
rect 30057 39704 30121 39750
rect 30167 39704 30216 39750
rect 30057 39701 30216 39704
rect 30268 39750 30365 39753
rect 30268 39704 30284 39750
rect 30330 39704 30365 39750
rect 30268 39701 30365 39704
rect 29283 39661 30365 39701
rect 30583 39788 30637 39834
rect 30683 39828 30855 39834
rect 30901 39828 31040 39874
rect 33484 39870 33495 40292
rect 33541 39870 33552 40292
rect 34964 40317 35082 40374
rect 36438 40329 36554 40429
rect 37853 40424 38161 40429
rect 38658 40449 39723 40463
rect 34964 40285 36360 40317
rect 34228 40215 34718 40256
rect 34228 40198 34267 40215
rect 34319 40198 34447 40215
rect 34499 40198 34627 40215
rect 33671 40152 33684 40198
rect 33730 40152 33787 40198
rect 33833 40152 33890 40198
rect 33936 40152 33993 40198
rect 34039 40152 34096 40198
rect 34142 40152 34199 40198
rect 34245 40163 34267 40198
rect 34245 40152 34302 40163
rect 34348 40152 34405 40198
rect 34499 40163 34508 40198
rect 34451 40152 34508 40163
rect 34554 40152 34612 40198
rect 34679 40163 34718 40215
rect 34964 40239 35273 40285
rect 35523 40239 35580 40285
rect 35626 40239 35683 40285
rect 35729 40239 35786 40285
rect 35832 40239 35889 40285
rect 35935 40239 35992 40285
rect 36038 40239 36095 40285
rect 36141 40239 36198 40285
rect 36244 40239 36301 40285
rect 36347 40239 36360 40285
rect 34964 40195 36360 40239
rect 34658 40152 34718 40163
rect 34228 40123 34718 40152
rect 36438 40189 36475 40329
rect 36521 40189 36554 40329
rect 35294 40061 36266 40095
rect 36438 40086 36554 40189
rect 36640 40329 36773 40349
rect 36640 40290 36697 40329
rect 36640 40238 36678 40290
rect 36640 40189 36697 40238
rect 36743 40189 36773 40329
rect 38658 40327 38726 40449
rect 39809 40443 44918 40481
rect 48765 40463 48778 40509
rect 48824 40463 48881 40509
rect 48927 40463 48943 40509
rect 49030 40463 49087 40509
rect 49133 40463 49154 40509
rect 49236 40463 49293 40509
rect 49339 40463 49365 40509
rect 49442 40463 49499 40509
rect 49545 40463 49576 40509
rect 49852 40463 49877 40509
rect 54085 40527 54540 40560
rect 50481 40467 51657 40494
rect 39809 40397 43739 40443
rect 43785 40397 43906 40443
rect 43952 40397 44071 40443
rect 44117 40397 44236 40443
rect 44282 40422 44918 40443
rect 48905 40423 49877 40463
rect 50044 40457 51657 40467
rect 44282 40397 44812 40422
rect 39809 40394 44812 40397
rect 39809 40348 39844 40394
rect 39890 40392 44812 40394
rect 39890 40348 39994 40392
rect 39809 40340 39994 40348
rect 40046 40376 44812 40392
rect 44858 40376 44925 40422
rect 44971 40376 45038 40422
rect 45084 40376 45151 40422
rect 45197 40376 45264 40422
rect 45310 40376 45323 40422
rect 48557 40377 48687 40417
rect 40046 40361 44918 40376
rect 40046 40340 40085 40361
rect 39809 40337 40085 40340
rect 36924 40317 37685 40324
rect 36923 40285 37931 40317
rect 36841 40239 36854 40285
rect 36900 40283 36971 40285
rect 36900 40239 36961 40283
rect 37017 40239 37088 40285
rect 37134 40283 37206 40285
rect 37134 40239 37172 40283
rect 37252 40239 37324 40285
rect 37370 40283 37442 40285
rect 37370 40239 37384 40283
rect 36923 40231 36961 40239
rect 37013 40231 37172 40239
rect 37224 40231 37384 40239
rect 37436 40239 37442 40283
rect 37488 40283 37909 40285
rect 37488 40239 37595 40283
rect 37436 40231 37595 40239
rect 37647 40239 37909 40283
rect 37955 40239 38026 40285
rect 38072 40239 38143 40285
rect 38189 40239 38261 40285
rect 38307 40239 38379 40285
rect 38425 40239 38497 40285
rect 38543 40239 38556 40285
rect 37647 40231 37931 40239
rect 36923 40198 37931 40231
rect 36923 40197 37685 40198
rect 36924 40191 37685 40197
rect 36640 40166 36773 40189
rect 38658 40187 38669 40327
rect 38715 40187 38726 40327
rect 39014 40285 39323 40317
rect 39492 40285 39608 40317
rect 39008 40239 39021 40285
rect 39067 40239 39144 40285
rect 39190 40239 39267 40285
rect 39313 40239 39326 40285
rect 39492 40239 39641 40285
rect 39687 40239 39730 40285
rect 38658 40176 38726 40187
rect 36438 40061 36953 40086
rect 37439 40083 37931 40086
rect 37439 40061 38161 40083
rect 35260 40015 35273 40061
rect 35523 40055 35580 40061
rect 35523 40015 35543 40055
rect 35626 40015 35683 40061
rect 35729 40055 35786 40061
rect 35729 40015 35754 40055
rect 35832 40015 35889 40061
rect 35935 40055 35992 40061
rect 35935 40015 35965 40055
rect 36038 40015 36095 40061
rect 36141 40055 36198 40061
rect 36141 40015 36176 40055
rect 36244 40015 36301 40061
rect 36347 40015 36360 40061
rect 36438 40015 36854 40061
rect 36900 40015 36971 40061
rect 37017 40015 37088 40061
rect 37134 40015 37206 40061
rect 37252 40015 37324 40061
rect 37370 40015 37442 40061
rect 37488 40043 37909 40061
rect 37488 40015 37891 40043
rect 37955 40015 38026 40061
rect 38072 40043 38143 40061
rect 38123 40015 38143 40043
rect 38189 40015 38261 40061
rect 38307 40015 38379 40061
rect 38425 40015 38497 40061
rect 38543 40015 38556 40061
rect 33781 39974 34089 40009
rect 35294 40003 35332 40015
rect 35384 40003 35543 40015
rect 35595 40003 35754 40015
rect 35806 40003 35965 40015
rect 36017 40003 36176 40015
rect 36228 40003 36266 40015
rect 33671 39928 33684 39974
rect 33730 39928 33787 39974
rect 33833 39969 33890 39974
rect 33871 39928 33890 39969
rect 33936 39928 33993 39974
rect 34039 39969 34096 39974
rect 34051 39928 34096 39969
rect 34142 39928 34199 39974
rect 34245 39928 34302 39974
rect 34348 39928 34405 39974
rect 34451 39928 34508 39974
rect 34554 39928 34612 39974
rect 34658 39928 34671 39974
rect 35294 39963 36266 40003
rect 36438 39966 36953 40015
rect 37439 39991 37891 40015
rect 37943 39991 38071 40015
rect 38123 39991 38161 40015
rect 37439 39966 38161 39991
rect 37853 39950 38161 39966
rect 33781 39917 33819 39928
rect 33871 39917 33999 39928
rect 34051 39917 34089 39928
rect 33781 39876 34089 39917
rect 33484 39859 33552 39870
rect 30683 39794 31040 39828
rect 30683 39788 32842 39794
rect 30583 39753 32842 39788
rect 34247 39787 35008 39794
rect 30583 39701 30854 39753
rect 30906 39701 31065 39753
rect 31117 39701 31276 39753
rect 31328 39750 31486 39753
rect 31538 39750 31697 39753
rect 31749 39750 31909 39753
rect 31961 39750 32120 39753
rect 32172 39750 32330 39753
rect 32382 39750 32541 39753
rect 32593 39750 32752 39753
rect 32804 39750 32842 39753
rect 34246 39753 35008 39787
rect 34246 39750 34284 39753
rect 34336 39750 34495 39753
rect 34547 39750 34707 39753
rect 31328 39704 31349 39750
rect 33323 39704 33336 39750
rect 33671 39704 33684 39750
rect 33730 39704 33787 39750
rect 33833 39704 33890 39750
rect 33936 39704 33993 39750
rect 34039 39704 34096 39750
rect 34142 39704 34199 39750
rect 34245 39704 34284 39750
rect 34348 39704 34405 39750
rect 34451 39704 34495 39750
rect 34554 39704 34612 39750
rect 34658 39704 34707 39750
rect 31328 39701 31486 39704
rect 31538 39701 31697 39704
rect 31749 39701 31909 39704
rect 31961 39701 32120 39704
rect 32172 39701 32330 39704
rect 32382 39701 32541 39704
rect 32593 39701 32752 39704
rect 32804 39701 32842 39704
rect 30583 39666 32842 39701
rect 34246 39701 34284 39704
rect 34336 39701 34495 39704
rect 34547 39701 34707 39704
rect 34759 39701 34918 39753
rect 34970 39701 35008 39753
rect 34246 39667 35008 39701
rect 29544 39660 30306 39661
rect 27387 39544 29196 39620
rect 27387 39503 29116 39544
rect 27387 39457 28810 39503
rect 28856 39498 29116 39503
rect 29162 39498 29196 39544
rect 28856 39457 29196 39498
rect 27387 39381 29196 39457
rect 27387 39340 29116 39381
rect 27387 39294 28810 39340
rect 28856 39335 29116 39340
rect 29162 39335 29196 39381
rect 28856 39294 29196 39335
rect 27387 39217 29196 39294
rect 27387 39177 29116 39217
rect 27387 39131 28810 39177
rect 28856 39171 29116 39177
rect 29162 39171 29196 39217
rect 28856 39131 29196 39171
rect 27387 39054 29196 39131
rect 27387 39013 29116 39054
rect 27387 38967 28810 39013
rect 28856 39008 29116 39013
rect 29162 39008 29196 39054
rect 28856 38967 29196 39008
rect 27387 38853 29196 38967
rect 30583 39620 30637 39666
rect 30683 39660 32842 39666
rect 34247 39660 35008 39667
rect 35182 39787 36364 39794
rect 35182 39753 36958 39787
rect 35182 39701 35220 39753
rect 35272 39701 35430 39753
rect 35482 39701 35641 39753
rect 35693 39701 35853 39753
rect 35905 39701 36064 39753
rect 36116 39701 36274 39753
rect 36326 39750 36958 39753
rect 36326 39704 36489 39750
rect 36723 39704 36958 39750
rect 36326 39701 36958 39704
rect 35182 39667 36958 39701
rect 37946 39753 38842 39794
rect 37946 39750 38330 39753
rect 38382 39750 38541 39753
rect 37946 39704 37957 39750
rect 38473 39704 38541 39750
rect 37946 39701 38330 39704
rect 38382 39701 38541 39704
rect 38593 39701 38752 39753
rect 38804 39701 38842 39753
rect 35182 39660 36364 39667
rect 37946 39660 38842 39701
rect 39014 39753 39323 40239
rect 39014 39701 39052 39753
rect 39104 39750 39232 39753
rect 39108 39704 39220 39750
rect 39104 39701 39232 39704
rect 39284 39701 39323 39753
rect 30683 39626 31040 39660
rect 30683 39620 30855 39626
rect 30583 39580 30855 39620
rect 30901 39580 31040 39626
rect 30583 39503 31040 39580
rect 33484 39584 33552 39595
rect 33019 39529 33327 39570
rect 33019 39526 33057 39529
rect 33109 39526 33237 39529
rect 33289 39526 33327 39529
rect 30583 39457 30637 39503
rect 30683 39462 31040 39503
rect 31336 39480 31349 39526
rect 33323 39480 33336 39526
rect 30683 39457 30855 39462
rect 30583 39416 30855 39457
rect 30901 39416 31040 39462
rect 33019 39477 33057 39480
rect 33109 39477 33237 39480
rect 33289 39477 33327 39480
rect 33019 39437 33327 39477
rect 30583 39340 31040 39416
rect 30583 39294 30637 39340
rect 30683 39324 31040 39340
rect 30683 39302 31493 39324
rect 30683 39299 31349 39302
rect 30683 39294 30855 39299
rect 30583 39253 30855 39294
rect 30901 39256 31349 39299
rect 33323 39256 33336 39302
rect 30901 39253 31493 39256
rect 30583 39205 31493 39253
rect 30583 39177 31040 39205
rect 30583 39131 30637 39177
rect 30683 39136 31040 39177
rect 30683 39131 30855 39136
rect 30583 39090 30855 39131
rect 30901 39090 31040 39136
rect 33484 39162 33495 39584
rect 33541 39162 33552 39584
rect 33781 39537 34089 39578
rect 33781 39526 33819 39537
rect 33871 39526 33999 39537
rect 34051 39526 34089 39537
rect 33671 39480 33684 39526
rect 33730 39480 33787 39526
rect 33871 39485 33890 39526
rect 33833 39480 33890 39485
rect 33936 39480 33993 39526
rect 34051 39485 34096 39526
rect 34039 39480 34096 39485
rect 34142 39480 34199 39526
rect 34245 39480 34302 39526
rect 34348 39480 34405 39526
rect 34451 39480 34508 39526
rect 34554 39480 34612 39526
rect 34658 39480 34671 39526
rect 33781 39445 34089 39480
rect 35294 39451 36266 39491
rect 37853 39488 38161 39504
rect 35294 39439 35332 39451
rect 35384 39439 35543 39451
rect 35595 39439 35754 39451
rect 35806 39439 35965 39451
rect 36017 39439 36176 39451
rect 36228 39439 36266 39451
rect 36438 39439 36953 39488
rect 37439 39463 38161 39488
rect 37439 39439 37891 39463
rect 37943 39439 38071 39463
rect 38123 39439 38161 39463
rect 35260 39393 35273 39439
rect 35523 39399 35543 39439
rect 35523 39393 35580 39399
rect 35626 39393 35683 39439
rect 35729 39399 35754 39439
rect 35729 39393 35786 39399
rect 35832 39393 35889 39439
rect 35935 39399 35965 39439
rect 35935 39393 35992 39399
rect 36038 39393 36095 39439
rect 36141 39399 36176 39439
rect 36141 39393 36198 39399
rect 36244 39393 36301 39439
rect 36347 39393 36360 39439
rect 36438 39393 36854 39439
rect 36900 39393 36971 39439
rect 37017 39393 37088 39439
rect 37134 39393 37206 39439
rect 37252 39393 37324 39439
rect 37370 39393 37442 39439
rect 37488 39411 37891 39439
rect 37488 39393 37909 39411
rect 37955 39393 38026 39439
rect 38123 39411 38143 39439
rect 38072 39393 38143 39411
rect 38189 39393 38261 39439
rect 38307 39393 38379 39439
rect 38425 39393 38497 39439
rect 38543 39393 38556 39439
rect 35294 39359 36266 39393
rect 36438 39368 36953 39393
rect 37439 39371 38161 39393
rect 37439 39368 37931 39371
rect 34228 39302 34718 39331
rect 33671 39256 33684 39302
rect 33730 39256 33787 39302
rect 33833 39256 33890 39302
rect 33936 39256 33993 39302
rect 34039 39256 34096 39302
rect 34142 39256 34199 39302
rect 34245 39291 34302 39302
rect 34245 39256 34267 39291
rect 34348 39256 34405 39302
rect 34451 39291 34508 39302
rect 34499 39256 34508 39291
rect 34554 39256 34612 39302
rect 34658 39291 34718 39302
rect 34228 39239 34267 39256
rect 34319 39239 34447 39256
rect 34499 39239 34627 39256
rect 34679 39239 34718 39291
rect 36438 39265 36554 39368
rect 34228 39198 34718 39239
rect 34964 39215 36360 39259
rect 30583 39013 31040 39090
rect 33019 39081 33327 39122
rect 33019 39078 33057 39081
rect 33109 39078 33237 39081
rect 33289 39078 33327 39081
rect 33484 39080 33552 39162
rect 34964 39169 35273 39215
rect 35523 39169 35580 39215
rect 35626 39169 35683 39215
rect 35729 39169 35786 39215
rect 35832 39169 35889 39215
rect 35935 39169 35992 39215
rect 36038 39169 36095 39215
rect 36141 39169 36198 39215
rect 36244 39169 36301 39215
rect 36347 39169 36360 39215
rect 34964 39137 36360 39169
rect 34964 39080 35082 39137
rect 31336 39032 31349 39078
rect 33323 39032 33336 39078
rect 33484 39043 35082 39080
rect 30583 38967 30637 39013
rect 30683 38973 31040 39013
rect 33019 39029 33057 39032
rect 33109 39029 33237 39032
rect 33289 39029 33327 39032
rect 33019 38989 33327 39029
rect 33484 38997 33816 39043
rect 33862 38997 34002 39043
rect 34048 38997 34189 39043
rect 34235 38997 34376 39043
rect 34422 38997 34562 39043
rect 34608 38997 35082 39043
rect 36438 39125 36475 39265
rect 36521 39125 36554 39265
rect 33484 38989 35082 38997
rect 35294 38991 36266 39031
rect 36438 39025 36554 39125
rect 36640 39265 36773 39288
rect 36640 39216 36697 39265
rect 36640 39164 36678 39216
rect 36640 39125 36697 39164
rect 36743 39125 36773 39265
rect 38658 39267 38726 39278
rect 36924 39257 37685 39263
rect 36923 39256 37685 39257
rect 36923 39223 37931 39256
rect 36923 39215 36961 39223
rect 37013 39215 37172 39223
rect 37224 39215 37384 39223
rect 36841 39169 36854 39215
rect 36900 39171 36961 39215
rect 36900 39169 36971 39171
rect 37017 39169 37088 39215
rect 37134 39171 37172 39215
rect 37134 39169 37206 39171
rect 37252 39169 37324 39215
rect 37370 39171 37384 39215
rect 37436 39215 37595 39223
rect 37436 39171 37442 39215
rect 37370 39169 37442 39171
rect 37488 39171 37595 39215
rect 37647 39215 37931 39223
rect 37647 39171 37909 39215
rect 37488 39169 37909 39171
rect 37955 39169 38026 39215
rect 38072 39169 38143 39215
rect 38189 39169 38261 39215
rect 38307 39169 38379 39215
rect 38425 39169 38497 39215
rect 38543 39169 38556 39215
rect 36923 39137 37931 39169
rect 36924 39130 37685 39137
rect 36640 39105 36773 39125
rect 38658 39127 38669 39267
rect 38715 39127 38726 39267
rect 39014 39215 39323 39701
rect 39492 39787 39608 40239
rect 39923 40206 40085 40337
rect 39923 40154 39994 40206
rect 40046 40154 40085 40206
rect 39923 40114 40085 40154
rect 39737 40018 39865 40031
rect 39737 39991 39866 40018
rect 39737 39974 39775 39991
rect 39827 39974 39866 39991
rect 39727 39928 39740 39974
rect 39827 39939 39862 39974
rect 39786 39928 39862 39939
rect 39908 39928 39985 39974
rect 40031 39928 40108 39974
rect 40154 39928 40167 39974
rect 40246 39963 40362 40361
rect 42229 40222 44509 40263
rect 42229 40170 43445 40222
rect 43497 40170 44509 40222
rect 42229 40130 44509 40170
rect 44341 40086 44509 40130
rect 44341 40040 44358 40086
rect 44498 40040 44509 40086
rect 39737 39899 39866 39928
rect 40246 39917 40281 39963
rect 40327 39917 40362 39963
rect 40246 39880 40362 39917
rect 40718 39991 43524 40032
rect 44341 40029 44509 40040
rect 40718 39939 41935 39991
rect 41987 39939 43524 39991
rect 40718 39898 43524 39939
rect 44605 39974 44721 40361
rect 45400 40331 48379 40372
rect 45400 40317 46731 40331
rect 45400 40271 45464 40317
rect 45604 40279 46731 40317
rect 46783 40279 48379 40331
rect 45604 40271 48379 40279
rect 44901 40215 45241 40256
rect 45400 40238 48379 40271
rect 48557 40325 48596 40377
rect 48648 40325 48687 40377
rect 48557 40302 48687 40325
rect 50044 40411 50516 40457
rect 50562 40411 50703 40457
rect 50749 40411 50890 40457
rect 50936 40411 51076 40457
rect 51122 40411 51263 40457
rect 51309 40411 51657 40457
rect 51797 40447 52105 40487
rect 51797 40422 51835 40447
rect 51887 40422 52015 40447
rect 52067 40422 52105 40447
rect 54085 40481 54223 40527
rect 54269 40487 54540 40527
rect 54269 40481 54440 40487
rect 54085 40441 54440 40481
rect 54486 40441 54540 40487
rect 50044 40374 51657 40411
rect 51789 40376 51802 40422
rect 53776 40376 53789 40422
rect 50044 40317 50160 40374
rect 44901 40198 44939 40215
rect 44991 40198 45151 40215
rect 45203 40198 45241 40215
rect 44799 40152 44812 40198
rect 44858 40152 44925 40198
rect 44991 40163 45038 40198
rect 44971 40152 45038 40163
rect 45084 40152 45151 40198
rect 45203 40163 45264 40198
rect 45197 40152 45264 40163
rect 45310 40152 45323 40198
rect 48557 40162 48622 40302
rect 48668 40162 48687 40302
rect 49820 40285 50160 40317
rect 48765 40239 48778 40285
rect 48824 40239 48881 40285
rect 48927 40239 48984 40285
rect 49030 40239 49087 40285
rect 49133 40239 49190 40285
rect 49236 40239 49293 40285
rect 49339 40239 49396 40285
rect 49442 40239 49499 40285
rect 49545 40239 49602 40285
rect 49852 40239 50160 40285
rect 51589 40322 51657 40374
rect 51797 40354 52105 40376
rect 49820 40198 50160 40239
rect 50262 40215 50812 40256
rect 48557 40159 48687 40162
rect 44901 40123 45241 40152
rect 48557 40107 48596 40159
rect 48648 40107 48687 40159
rect 50262 40163 50300 40215
rect 50352 40198 50511 40215
rect 50563 40198 50722 40215
rect 50352 40163 50467 40198
rect 50563 40163 50571 40198
rect 50262 40152 50467 40163
rect 50513 40152 50571 40163
rect 50617 40152 50674 40198
rect 50720 40163 50722 40198
rect 50774 40198 50812 40215
rect 50774 40163 50777 40198
rect 50720 40152 50777 40163
rect 50823 40152 50880 40198
rect 50926 40152 50983 40198
rect 51029 40152 51086 40198
rect 51132 40152 51189 40198
rect 51235 40152 51292 40198
rect 51338 40152 51395 40198
rect 51441 40152 51454 40198
rect 50262 40123 50812 40152
rect 48557 40066 48687 40107
rect 48905 40061 49877 40092
rect 48765 40015 48778 40061
rect 48824 40015 48881 40061
rect 48927 40052 48984 40061
rect 48927 40015 48943 40052
rect 49030 40015 49087 40061
rect 49133 40052 49190 40061
rect 49133 40015 49154 40052
rect 49236 40015 49293 40061
rect 49339 40052 49396 40061
rect 49339 40015 49365 40052
rect 49442 40015 49499 40061
rect 49545 40052 49602 40061
rect 49545 40015 49576 40052
rect 49852 40015 49877 40061
rect 48905 40000 48943 40015
rect 48995 40000 49154 40015
rect 49206 40000 49365 40015
rect 49417 40000 49576 40015
rect 49628 40000 49787 40015
rect 49839 40000 49877 40015
rect 44605 39928 44812 39974
rect 44858 39928 44925 39974
rect 44971 39928 45038 39974
rect 45084 39928 45151 39974
rect 45197 39928 45264 39974
rect 45310 39928 45323 39974
rect 48905 39960 49877 40000
rect 51035 39977 51343 40017
rect 51035 39974 51073 39977
rect 51125 39974 51253 39977
rect 51305 39974 51343 39977
rect 43362 39891 43524 39898
rect 43362 39845 43373 39891
rect 43513 39845 43524 39891
rect 43362 39834 43524 39845
rect 45584 39914 48546 39950
rect 50454 39928 50467 39974
rect 50513 39928 50571 39974
rect 50617 39928 50674 39974
rect 50720 39928 50777 39974
rect 50823 39928 50880 39974
rect 50926 39928 50983 39974
rect 51029 39928 51073 39974
rect 51132 39928 51189 39974
rect 51235 39928 51253 39974
rect 51338 39928 51395 39974
rect 51441 39928 51454 39974
rect 45584 39868 45619 39914
rect 45665 39868 45777 39914
rect 45823 39868 45935 39914
rect 45981 39868 46093 39914
rect 46139 39868 46251 39914
rect 46297 39868 46409 39914
rect 46455 39868 46568 39914
rect 46614 39868 46726 39914
rect 46772 39868 46884 39914
rect 46930 39868 47042 39914
rect 47088 39868 47200 39914
rect 47246 39868 47358 39914
rect 47404 39868 47516 39914
rect 47562 39868 47675 39914
rect 47721 39868 47833 39914
rect 47879 39868 47991 39914
rect 48037 39868 48149 39914
rect 48195 39868 48307 39914
rect 48353 39868 48465 39914
rect 48511 39868 48546 39914
rect 51035 39925 51073 39928
rect 51125 39925 51253 39928
rect 51305 39925 51343 39928
rect 51035 39884 51343 39925
rect 51589 39900 51600 40322
rect 51646 39900 51657 40322
rect 54085 40323 54540 40441
rect 54085 40277 54440 40323
rect 54486 40277 54540 40323
rect 54085 40249 54540 40277
rect 53585 40198 54540 40249
rect 51789 40152 51802 40198
rect 53776 40160 54540 40198
rect 53776 40152 54440 40160
rect 53585 40130 54440 40152
rect 54085 40114 54440 40130
rect 54486 40114 54540 40160
rect 54085 40038 54540 40114
rect 51797 39984 52105 40024
rect 51797 39974 51835 39984
rect 51887 39974 52015 39984
rect 52067 39974 52105 39984
rect 54085 39992 54223 40038
rect 54269 39997 54540 40038
rect 54269 39992 54440 39997
rect 51789 39928 51802 39974
rect 53776 39928 53789 39974
rect 54085 39951 54440 39992
rect 54486 39951 54540 39997
rect 51589 39889 51657 39900
rect 51797 39891 52105 39928
rect 40215 39787 40523 39794
rect 40788 39787 42986 39801
rect 43753 39787 44514 39794
rect 39492 39764 42986 39787
rect 43704 39764 44514 39787
rect 39492 39753 44514 39764
rect 39492 39750 40253 39753
rect 39492 39704 39740 39750
rect 39786 39704 39862 39750
rect 39908 39704 39985 39750
rect 40031 39704 40108 39750
rect 40154 39704 40253 39750
rect 39492 39701 40253 39704
rect 40305 39701 40433 39753
rect 40485 39750 43790 39753
rect 40485 39704 40836 39750
rect 40882 39704 40994 39750
rect 41040 39704 41152 39750
rect 41198 39704 41310 39750
rect 41356 39704 41469 39750
rect 41515 39704 41627 39750
rect 41673 39704 41785 39750
rect 41831 39704 41943 39750
rect 41989 39704 42101 39750
rect 42147 39704 42259 39750
rect 42305 39704 42418 39750
rect 42464 39704 42576 39750
rect 42622 39704 42734 39750
rect 42780 39704 42892 39750
rect 42938 39704 43739 39750
rect 43785 39704 43790 39750
rect 40485 39701 43790 39704
rect 43842 39750 44001 39753
rect 43842 39704 43906 39750
rect 43952 39704 44001 39750
rect 43842 39701 44001 39704
rect 44053 39750 44213 39753
rect 44265 39750 44424 39753
rect 44053 39704 44071 39750
rect 44117 39704 44213 39750
rect 44282 39704 44424 39750
rect 44053 39701 44213 39704
rect 44265 39701 44424 39704
rect 44476 39701 44514 39753
rect 39492 39690 44514 39701
rect 39492 39667 42986 39690
rect 43704 39667 44514 39690
rect 39492 39215 39608 39667
rect 40215 39660 40523 39667
rect 40788 39653 42986 39667
rect 43753 39660 44514 39667
rect 44796 39787 45346 39794
rect 45584 39787 48546 39868
rect 54085 39874 54540 39951
rect 54085 39828 54223 39874
rect 54269 39834 54540 39874
rect 54269 39828 54440 39834
rect 54085 39794 54440 39828
rect 48800 39787 49982 39794
rect 50308 39787 50859 39794
rect 44796 39753 49982 39787
rect 44796 39750 44834 39753
rect 44886 39750 45045 39753
rect 45097 39750 45256 39753
rect 45308 39750 48838 39753
rect 44796 39704 44812 39750
rect 44886 39704 44925 39750
rect 44971 39704 45038 39750
rect 45097 39704 45151 39750
rect 45197 39704 45256 39750
rect 45310 39704 45619 39750
rect 45665 39704 45777 39750
rect 45823 39704 45935 39750
rect 45981 39704 46093 39750
rect 46139 39704 46251 39750
rect 46297 39704 46409 39750
rect 46455 39704 46568 39750
rect 46614 39704 46726 39750
rect 46772 39704 46884 39750
rect 46930 39704 47042 39750
rect 47088 39704 47200 39750
rect 47246 39704 47358 39750
rect 47404 39704 47516 39750
rect 47562 39704 47675 39750
rect 47721 39704 47833 39750
rect 47879 39704 47991 39750
rect 48037 39704 48149 39750
rect 48195 39704 48307 39750
rect 48353 39704 48465 39750
rect 48511 39704 48838 39750
rect 44796 39701 44834 39704
rect 44886 39701 45045 39704
rect 45097 39701 45256 39704
rect 45308 39701 48838 39704
rect 48890 39701 49048 39753
rect 49100 39701 49259 39753
rect 49311 39701 49471 39753
rect 49523 39701 49682 39753
rect 49734 39701 49892 39753
rect 49944 39701 49982 39753
rect 44796 39667 49982 39701
rect 50307 39753 50859 39787
rect 50307 39701 50346 39753
rect 50398 39750 50557 39753
rect 50609 39750 50768 39753
rect 50820 39750 50859 39753
rect 52278 39788 54440 39794
rect 54486 39788 54540 39834
rect 55927 40487 57736 40601
rect 55927 40444 56267 40487
rect 55927 40398 55961 40444
rect 56007 40441 56267 40444
rect 56313 40441 57736 40487
rect 56007 40398 57736 40441
rect 55927 40323 57736 40398
rect 55927 40281 56267 40323
rect 55927 40235 55961 40281
rect 56007 40277 56267 40281
rect 56313 40277 57736 40323
rect 56007 40235 57736 40277
rect 55927 40160 57736 40235
rect 55927 40117 56267 40160
rect 55927 40071 55961 40117
rect 56007 40114 56267 40117
rect 56313 40114 57736 40160
rect 56007 40071 57736 40114
rect 55927 39997 57736 40071
rect 55927 39954 56267 39997
rect 55927 39908 55961 39954
rect 56007 39951 56267 39954
rect 56313 39951 57736 39997
rect 56007 39908 57736 39951
rect 55927 39834 57736 39908
rect 52278 39753 54540 39788
rect 52278 39750 52316 39753
rect 52368 39750 52527 39753
rect 52579 39750 52738 39753
rect 52790 39750 52948 39753
rect 53000 39750 53159 39753
rect 53211 39750 53371 39753
rect 53423 39750 53582 39753
rect 53634 39750 53792 39753
rect 50398 39704 50467 39750
rect 50513 39704 50557 39750
rect 50617 39704 50674 39750
rect 50720 39704 50768 39750
rect 50823 39704 50880 39750
rect 50926 39704 50983 39750
rect 51029 39704 51086 39750
rect 51132 39704 51189 39750
rect 51235 39704 51292 39750
rect 51338 39704 51395 39750
rect 51441 39704 51454 39750
rect 51789 39704 51802 39750
rect 53776 39704 53792 39750
rect 50398 39701 50557 39704
rect 50609 39701 50768 39704
rect 50820 39701 50859 39704
rect 50307 39667 50859 39701
rect 44796 39660 45346 39667
rect 43362 39609 43524 39620
rect 39737 39526 39866 39555
rect 40246 39537 40362 39574
rect 43362 39563 43373 39609
rect 43513 39563 43524 39609
rect 43362 39556 43524 39563
rect 39727 39480 39740 39526
rect 39786 39515 39862 39526
rect 39827 39480 39862 39515
rect 39908 39480 39985 39526
rect 40031 39480 40108 39526
rect 40154 39480 40167 39526
rect 40246 39491 40281 39537
rect 40327 39491 40362 39537
rect 39737 39463 39775 39480
rect 39827 39463 39866 39480
rect 39737 39436 39866 39463
rect 39737 39423 39865 39436
rect 39923 39300 40085 39340
rect 39923 39248 39994 39300
rect 40046 39248 40085 39300
rect 39008 39169 39021 39215
rect 39067 39169 39144 39215
rect 39190 39169 39267 39215
rect 39313 39169 39326 39215
rect 39492 39169 39641 39215
rect 39687 39169 39730 39215
rect 39014 39137 39323 39169
rect 39492 39137 39608 39169
rect 37853 39025 38161 39030
rect 36438 38991 36953 39025
rect 37439 38991 38161 39025
rect 38658 39005 38726 39127
rect 39923 39117 40085 39248
rect 39809 39114 40085 39117
rect 39809 39106 39994 39114
rect 39809 39060 39844 39106
rect 39890 39062 39994 39106
rect 40046 39093 40085 39114
rect 40246 39093 40362 39491
rect 40718 39515 43524 39556
rect 45584 39586 48546 39667
rect 48800 39660 49982 39667
rect 50308 39660 50859 39667
rect 52278 39701 52316 39704
rect 52368 39701 52527 39704
rect 52579 39701 52738 39704
rect 52790 39701 52948 39704
rect 53000 39701 53159 39704
rect 53211 39701 53371 39704
rect 53423 39701 53582 39704
rect 53634 39701 53792 39704
rect 53844 39701 54003 39753
rect 54055 39701 54214 39753
rect 54266 39701 54540 39753
rect 52278 39666 54540 39701
rect 52278 39660 54440 39666
rect 45584 39540 45619 39586
rect 45665 39540 45777 39586
rect 45823 39540 45935 39586
rect 45981 39540 46093 39586
rect 46139 39540 46251 39586
rect 46297 39540 46409 39586
rect 46455 39540 46568 39586
rect 46614 39540 46726 39586
rect 46772 39540 46884 39586
rect 46930 39540 47042 39586
rect 47088 39540 47200 39586
rect 47246 39540 47358 39586
rect 47404 39540 47516 39586
rect 47562 39540 47675 39586
rect 47721 39540 47833 39586
rect 47879 39540 47991 39586
rect 48037 39540 48149 39586
rect 48195 39540 48307 39586
rect 48353 39540 48465 39586
rect 48511 39540 48546 39586
rect 54085 39626 54440 39660
rect 54085 39580 54223 39626
rect 54269 39620 54440 39626
rect 54486 39620 54540 39666
rect 54758 39753 55840 39794
rect 54758 39750 54855 39753
rect 54758 39704 54793 39750
rect 54839 39704 54855 39750
rect 54758 39701 54855 39704
rect 54907 39750 55066 39753
rect 54907 39704 54956 39750
rect 55002 39704 55066 39750
rect 54907 39701 55066 39704
rect 55118 39750 55278 39753
rect 55330 39750 55489 39753
rect 55164 39704 55278 39750
rect 55330 39704 55439 39750
rect 55485 39704 55489 39750
rect 55118 39701 55278 39704
rect 55330 39701 55489 39704
rect 55541 39750 55840 39753
rect 55541 39704 55599 39750
rect 55645 39704 55760 39750
rect 55806 39704 55840 39750
rect 55541 39701 55840 39704
rect 54758 39661 55840 39701
rect 55927 39788 56267 39834
rect 56313 39788 57736 39834
rect 55927 39666 57736 39788
rect 54817 39660 55579 39661
rect 54269 39580 54540 39620
rect 40718 39463 41935 39515
rect 41987 39463 43524 39515
rect 40718 39422 43524 39463
rect 44605 39480 44812 39526
rect 44858 39480 44925 39526
rect 44971 39480 45038 39526
rect 45084 39480 45151 39526
rect 45197 39480 45264 39526
rect 45310 39480 45323 39526
rect 45584 39504 48546 39540
rect 51035 39529 51343 39570
rect 51035 39526 51073 39529
rect 51125 39526 51253 39529
rect 51305 39526 51343 39529
rect 51589 39554 51657 39565
rect 44341 39414 44509 39425
rect 44341 39368 44358 39414
rect 44498 39368 44509 39414
rect 44341 39324 44509 39368
rect 42229 39284 44509 39324
rect 42229 39232 43445 39284
rect 43497 39232 44509 39284
rect 42229 39191 44509 39232
rect 44605 39093 44721 39480
rect 48905 39454 49877 39494
rect 50454 39480 50467 39526
rect 50513 39480 50571 39526
rect 50617 39480 50674 39526
rect 50720 39480 50777 39526
rect 50823 39480 50880 39526
rect 50926 39480 50983 39526
rect 51029 39480 51073 39526
rect 51132 39480 51189 39526
rect 51235 39480 51253 39526
rect 51338 39480 51395 39526
rect 51441 39480 51454 39526
rect 48905 39439 48943 39454
rect 48995 39439 49154 39454
rect 49206 39439 49365 39454
rect 49417 39439 49576 39454
rect 49628 39439 49787 39454
rect 49839 39439 49877 39454
rect 48765 39393 48778 39439
rect 48824 39393 48881 39439
rect 48927 39402 48943 39439
rect 48927 39393 48984 39402
rect 49030 39393 49087 39439
rect 49133 39402 49154 39439
rect 49133 39393 49190 39402
rect 49236 39393 49293 39439
rect 49339 39402 49365 39439
rect 49339 39393 49396 39402
rect 49442 39393 49499 39439
rect 49545 39402 49576 39439
rect 49545 39393 49602 39402
rect 49852 39393 49877 39439
rect 51035 39477 51073 39480
rect 51125 39477 51253 39480
rect 51305 39477 51343 39480
rect 51035 39437 51343 39477
rect 48557 39347 48687 39388
rect 48905 39362 49877 39393
rect 44901 39302 45241 39331
rect 44799 39256 44812 39302
rect 44858 39256 44925 39302
rect 44971 39291 45038 39302
rect 44991 39256 45038 39291
rect 45084 39256 45151 39302
rect 45197 39291 45264 39302
rect 45203 39256 45264 39291
rect 45310 39256 45323 39302
rect 48557 39295 48596 39347
rect 48648 39295 48687 39347
rect 48557 39292 48687 39295
rect 44901 39239 44939 39256
rect 44991 39239 45151 39256
rect 45203 39239 45241 39256
rect 44901 39198 45241 39239
rect 45400 39183 48379 39216
rect 45400 39137 45464 39183
rect 45604 39175 48379 39183
rect 45604 39137 47108 39175
rect 45400 39123 47108 39137
rect 47160 39123 48379 39175
rect 40046 39078 44918 39093
rect 45400 39082 48379 39123
rect 48557 39152 48622 39292
rect 48668 39152 48687 39292
rect 50262 39302 50812 39331
rect 50262 39291 50467 39302
rect 50513 39291 50571 39302
rect 49820 39215 50160 39256
rect 48765 39169 48778 39215
rect 48824 39169 48881 39215
rect 48927 39169 48984 39215
rect 49030 39169 49087 39215
rect 49133 39169 49190 39215
rect 49236 39169 49293 39215
rect 49339 39169 49396 39215
rect 49442 39169 49499 39215
rect 49545 39169 49602 39215
rect 49852 39169 50160 39215
rect 50262 39239 50300 39291
rect 50352 39256 50467 39291
rect 50563 39256 50571 39291
rect 50617 39256 50674 39302
rect 50720 39291 50777 39302
rect 50720 39256 50722 39291
rect 50352 39239 50511 39256
rect 50563 39239 50722 39256
rect 50774 39256 50777 39291
rect 50823 39256 50880 39302
rect 50926 39256 50983 39302
rect 51029 39256 51086 39302
rect 51132 39256 51189 39302
rect 51235 39256 51292 39302
rect 51338 39256 51395 39302
rect 51441 39256 51454 39302
rect 50774 39239 50812 39256
rect 50262 39198 50812 39239
rect 48557 39129 48687 39152
rect 49820 39137 50160 39169
rect 40046 39062 44812 39078
rect 39890 39060 44812 39062
rect 39809 39057 44812 39060
rect 39809 39011 43739 39057
rect 43785 39011 43906 39057
rect 43952 39011 44071 39057
rect 44117 39011 44236 39057
rect 44282 39032 44812 39057
rect 44858 39032 44925 39078
rect 44971 39032 45038 39078
rect 45084 39032 45151 39078
rect 45197 39032 45264 39078
rect 45310 39032 45323 39078
rect 48557 39077 48596 39129
rect 48648 39077 48687 39129
rect 48557 39037 48687 39077
rect 50044 39080 50160 39137
rect 51589 39132 51600 39554
rect 51646 39132 51657 39554
rect 51797 39526 52105 39563
rect 51789 39480 51802 39526
rect 53776 39480 53789 39526
rect 54085 39503 54540 39580
rect 51797 39470 51835 39480
rect 51887 39470 52015 39480
rect 52067 39470 52105 39480
rect 51797 39430 52105 39470
rect 54085 39462 54440 39503
rect 54085 39416 54223 39462
rect 54269 39457 54440 39462
rect 54486 39457 54540 39503
rect 54269 39416 54540 39457
rect 54085 39340 54540 39416
rect 54085 39324 54440 39340
rect 53585 39302 54440 39324
rect 51789 39256 51802 39302
rect 53776 39294 54440 39302
rect 54486 39294 54540 39340
rect 53776 39256 54540 39294
rect 53585 39205 54540 39256
rect 51589 39080 51657 39132
rect 54085 39177 54540 39205
rect 54085 39131 54440 39177
rect 54486 39131 54540 39177
rect 50044 39043 51657 39080
rect 51797 39078 52105 39100
rect 44282 39011 44918 39032
rect 38658 38991 39723 39005
rect 30683 38967 30855 38973
rect 30583 38927 30855 38967
rect 30901 38927 31040 38973
rect 33484 38960 34643 38989
rect 35260 38945 35273 38991
rect 35523 38945 35543 38991
rect 35626 38945 35683 38991
rect 35729 38945 35754 38991
rect 35832 38945 35889 38991
rect 35935 38945 35965 38991
rect 36038 38945 36095 38991
rect 36141 38945 36176 38991
rect 36244 38945 36301 38991
rect 36347 38945 36360 38991
rect 36438 38945 36854 38991
rect 36900 38945 36971 38991
rect 37017 38945 37088 38991
rect 37134 38945 37206 38991
rect 37252 38945 37324 38991
rect 37370 38945 37442 38991
rect 37488 38989 37909 38991
rect 37488 38945 37891 38989
rect 37955 38945 38026 38991
rect 38072 38989 38143 38991
rect 38123 38945 38143 38989
rect 38189 38945 38261 38991
rect 38307 38945 38379 38991
rect 38425 38945 38497 38991
rect 38543 38945 38556 38991
rect 38658 38945 39021 38991
rect 39067 38945 39144 38991
rect 39190 38945 39267 38991
rect 39313 38945 39641 38991
rect 39687 38945 39730 38991
rect 39809 38973 44918 39011
rect 48905 38991 49877 39031
rect 48765 38945 48778 38991
rect 48824 38945 48881 38991
rect 48927 38945 48943 38991
rect 49030 38945 49087 38991
rect 49133 38945 49154 38991
rect 49236 38945 49293 38991
rect 49339 38945 49365 38991
rect 49442 38945 49499 38991
rect 49545 38945 49576 38991
rect 49852 38945 49877 38991
rect 50044 38997 50516 39043
rect 50562 38997 50703 39043
rect 50749 38997 50890 39043
rect 50936 38997 51076 39043
rect 51122 38997 51263 39043
rect 51309 38997 51657 39043
rect 51789 39032 51802 39078
rect 53776 39032 53789 39078
rect 50044 38987 51657 38997
rect 50481 38960 51657 38987
rect 51797 39007 51835 39032
rect 51887 39007 52015 39032
rect 52067 39007 52105 39032
rect 51797 38967 52105 39007
rect 54085 39013 54540 39131
rect 54085 38973 54440 39013
rect 30583 38894 31040 38927
rect 35294 38939 35332 38945
rect 35384 38939 35543 38945
rect 35595 38939 35754 38945
rect 35806 38939 35965 38945
rect 36017 38939 36176 38945
rect 36228 38939 36266 38945
rect 34870 38894 35025 38901
rect 35294 38899 36266 38939
rect 36438 38905 36953 38945
rect 37439 38937 37891 38945
rect 37943 38937 38071 38945
rect 38123 38937 38161 38945
rect 37439 38905 38161 38937
rect 37853 38897 38161 38905
rect 27387 38801 27790 38853
rect 27842 38801 28001 38853
rect 28053 38801 28212 38853
rect 28264 38801 28423 38853
rect 28475 38801 28634 38853
rect 28686 38850 28845 38853
rect 28686 38804 28810 38850
rect 28686 38801 28845 38804
rect 28897 38801 29056 38853
rect 29108 38801 29196 38853
rect 27387 38687 29196 38801
rect 29283 38853 30365 38894
rect 29283 38850 29582 38853
rect 29283 38804 29317 38850
rect 29363 38804 29478 38850
rect 29524 38804 29582 38850
rect 29283 38801 29582 38804
rect 29634 38850 29793 38853
rect 29845 38850 30005 38853
rect 29634 38804 29638 38850
rect 29684 38804 29793 38850
rect 29845 38804 29959 38850
rect 29634 38801 29793 38804
rect 29845 38801 30005 38804
rect 30057 38850 30216 38853
rect 30057 38804 30121 38850
rect 30167 38804 30216 38850
rect 30057 38801 30216 38804
rect 30268 38850 30365 38853
rect 30268 38804 30284 38850
rect 30330 38804 30365 38850
rect 30268 38801 30365 38804
rect 29283 38761 30365 38801
rect 30583 38853 32842 38894
rect 30583 38850 30854 38853
rect 30583 38804 30637 38850
rect 30683 38804 30854 38850
rect 30583 38801 30854 38804
rect 30906 38801 31065 38853
rect 31117 38801 31276 38853
rect 31328 38801 31486 38853
rect 31538 38801 31697 38853
rect 31749 38801 31909 38853
rect 31961 38801 32120 38853
rect 32172 38801 32330 38853
rect 32382 38801 32541 38853
rect 32593 38801 32752 38853
rect 32804 38801 32842 38853
rect 29544 38760 30306 38761
rect 30583 38760 32842 38801
rect 34717 38853 35025 38894
rect 38658 38885 39723 38945
rect 48905 38939 48943 38945
rect 48995 38939 49154 38945
rect 49206 38939 49365 38945
rect 49417 38939 49576 38945
rect 49628 38939 49787 38945
rect 49839 38939 49877 38945
rect 48905 38899 49877 38939
rect 54085 38927 54223 38973
rect 54269 38967 54440 38973
rect 54486 38967 54540 39013
rect 54269 38927 54540 38967
rect 50099 38894 50255 38901
rect 54085 38894 54540 38927
rect 55927 39620 56267 39666
rect 56313 39620 57736 39666
rect 55927 39544 57736 39620
rect 55927 39498 55961 39544
rect 56007 39503 57736 39544
rect 56007 39498 56267 39503
rect 55927 39457 56267 39498
rect 56313 39457 57736 39503
rect 55927 39381 57736 39457
rect 55927 39335 55961 39381
rect 56007 39340 57736 39381
rect 56007 39335 56267 39340
rect 55927 39294 56267 39335
rect 56313 39294 57736 39340
rect 55927 39217 57736 39294
rect 55927 39171 55961 39217
rect 56007 39177 57736 39217
rect 56007 39171 56267 39177
rect 55927 39131 56267 39171
rect 56313 39131 57736 39177
rect 55927 39054 57736 39131
rect 55927 39008 55961 39054
rect 56007 39013 57736 39054
rect 56007 39008 56267 39013
rect 55927 38967 56267 39008
rect 56313 38967 57736 39013
rect 34717 38801 34755 38853
rect 34807 38850 34935 38853
rect 34807 38804 34916 38850
rect 34807 38801 34935 38804
rect 34987 38801 35025 38853
rect 34717 38760 35025 38801
rect 50099 38853 50408 38894
rect 50099 38801 50138 38853
rect 50190 38850 50318 38853
rect 50206 38804 50318 38850
rect 50190 38801 50318 38804
rect 50370 38801 50408 38853
rect 27387 38641 28810 38687
rect 28856 38644 29196 38687
rect 28856 38641 29116 38644
rect 27387 38598 29116 38641
rect 29162 38598 29196 38644
rect 27387 38523 29196 38598
rect 27387 38477 28810 38523
rect 28856 38481 29196 38523
rect 28856 38477 29116 38481
rect 27387 38435 29116 38477
rect 29162 38435 29196 38481
rect 27387 38360 29196 38435
rect 27387 38314 28810 38360
rect 28856 38317 29196 38360
rect 28856 38314 29116 38317
rect 27387 38271 29116 38314
rect 29162 38271 29196 38317
rect 27387 38197 29196 38271
rect 27387 38151 28810 38197
rect 28856 38154 29196 38197
rect 28856 38151 29116 38154
rect 27387 38108 29116 38151
rect 29162 38108 29196 38154
rect 27387 38034 29196 38108
rect 27387 37988 28810 38034
rect 28856 37988 29196 38034
rect 30583 38727 31040 38760
rect 34870 38753 35025 38760
rect 30583 38687 30855 38727
rect 30583 38641 30637 38687
rect 30683 38681 30855 38687
rect 30901 38681 31040 38727
rect 35294 38715 36266 38755
rect 37853 38749 38161 38757
rect 35294 38709 35332 38715
rect 35384 38709 35543 38715
rect 35595 38709 35754 38715
rect 35806 38709 35965 38715
rect 36017 38709 36176 38715
rect 36228 38709 36266 38715
rect 36438 38709 36953 38749
rect 37439 38717 38161 38749
rect 37439 38709 37891 38717
rect 37943 38709 38071 38717
rect 38123 38709 38161 38717
rect 38658 38709 39723 38769
rect 50099 38760 50408 38801
rect 52278 38853 54540 38894
rect 52278 38801 52316 38853
rect 52368 38801 52527 38853
rect 52579 38801 52738 38853
rect 52790 38801 52948 38853
rect 53000 38801 53159 38853
rect 53211 38801 53371 38853
rect 53423 38801 53582 38853
rect 53634 38801 53792 38853
rect 53844 38801 54003 38853
rect 54055 38801 54214 38853
rect 54266 38850 54540 38853
rect 54266 38804 54440 38850
rect 54486 38804 54540 38850
rect 54266 38801 54540 38804
rect 52278 38760 54540 38801
rect 54758 38853 55840 38894
rect 54758 38850 54855 38853
rect 54758 38804 54793 38850
rect 54839 38804 54855 38850
rect 54758 38801 54855 38804
rect 54907 38850 55066 38853
rect 54907 38804 54956 38850
rect 55002 38804 55066 38850
rect 54907 38801 55066 38804
rect 55118 38850 55278 38853
rect 55330 38850 55489 38853
rect 55164 38804 55278 38850
rect 55330 38804 55439 38850
rect 55485 38804 55489 38850
rect 55118 38801 55278 38804
rect 55330 38801 55489 38804
rect 55541 38850 55840 38853
rect 55541 38804 55599 38850
rect 55645 38804 55760 38850
rect 55806 38804 55840 38850
rect 55541 38801 55840 38804
rect 54758 38761 55840 38801
rect 55927 38853 57736 38967
rect 55927 38801 56015 38853
rect 56067 38801 56226 38853
rect 56278 38850 56437 38853
rect 56313 38804 56437 38850
rect 56278 38801 56437 38804
rect 56489 38801 56648 38853
rect 56700 38801 56859 38853
rect 56911 38801 57070 38853
rect 57122 38801 57281 38853
rect 57333 38801 57736 38853
rect 54817 38760 55579 38761
rect 48905 38715 49877 38755
rect 50099 38753 50255 38760
rect 48905 38709 48943 38715
rect 48995 38709 49154 38715
rect 49206 38709 49365 38715
rect 49417 38709 49576 38715
rect 49628 38709 49787 38715
rect 49839 38709 49877 38715
rect 30683 38641 31040 38681
rect 33484 38665 34643 38694
rect 30583 38564 31040 38641
rect 33019 38625 33327 38665
rect 33019 38622 33057 38625
rect 33109 38622 33237 38625
rect 33289 38622 33327 38625
rect 33484 38657 35082 38665
rect 35260 38663 35273 38709
rect 35523 38663 35543 38709
rect 35626 38663 35683 38709
rect 35729 38663 35754 38709
rect 35832 38663 35889 38709
rect 35935 38663 35965 38709
rect 36038 38663 36095 38709
rect 36141 38663 36176 38709
rect 36244 38663 36301 38709
rect 36347 38663 36360 38709
rect 36438 38663 36854 38709
rect 36900 38663 36971 38709
rect 37017 38663 37088 38709
rect 37134 38663 37206 38709
rect 37252 38663 37324 38709
rect 37370 38663 37442 38709
rect 37488 38665 37891 38709
rect 37488 38663 37909 38665
rect 37955 38663 38026 38709
rect 38123 38665 38143 38709
rect 38072 38663 38143 38665
rect 38189 38663 38261 38709
rect 38307 38663 38379 38709
rect 38425 38663 38497 38709
rect 38543 38663 38556 38709
rect 38658 38663 39021 38709
rect 39067 38663 39144 38709
rect 39190 38663 39267 38709
rect 39313 38663 39641 38709
rect 39687 38663 39730 38709
rect 31336 38576 31349 38622
rect 33323 38576 33336 38622
rect 33484 38611 33816 38657
rect 33862 38611 34002 38657
rect 34048 38611 34189 38657
rect 34235 38611 34376 38657
rect 34422 38611 34562 38657
rect 34608 38611 35082 38657
rect 35294 38623 36266 38663
rect 36438 38629 36953 38663
rect 37439 38629 38161 38663
rect 30583 38523 30855 38564
rect 30583 38477 30637 38523
rect 30683 38518 30855 38523
rect 30901 38518 31040 38564
rect 33019 38573 33057 38576
rect 33109 38573 33237 38576
rect 33289 38573 33327 38576
rect 33019 38532 33327 38573
rect 33484 38574 35082 38611
rect 30683 38477 31040 38518
rect 30583 38449 31040 38477
rect 33484 38492 33552 38574
rect 30583 38401 31493 38449
rect 30583 38360 30855 38401
rect 30583 38314 30637 38360
rect 30683 38355 30855 38360
rect 30901 38398 31493 38401
rect 30901 38355 31349 38398
rect 30683 38352 31349 38355
rect 33323 38352 33336 38398
rect 30683 38330 31493 38352
rect 30683 38314 31040 38330
rect 30583 38238 31040 38314
rect 30583 38197 30855 38238
rect 30583 38151 30637 38197
rect 30683 38192 30855 38197
rect 30901 38192 31040 38238
rect 30683 38151 31040 38192
rect 33019 38177 33327 38217
rect 33019 38174 33057 38177
rect 33109 38174 33237 38177
rect 33289 38174 33327 38177
rect 30583 38074 31040 38151
rect 31336 38128 31349 38174
rect 33323 38128 33336 38174
rect 33019 38125 33057 38128
rect 33109 38125 33237 38128
rect 33289 38125 33327 38128
rect 33019 38084 33327 38125
rect 30583 38034 30855 38074
rect 27387 37866 29196 37988
rect 27387 37820 28810 37866
rect 28856 37820 29196 37866
rect 29283 37953 30365 37994
rect 29283 37950 29582 37953
rect 29283 37904 29317 37950
rect 29363 37904 29478 37950
rect 29524 37904 29582 37950
rect 29283 37901 29582 37904
rect 29634 37950 29793 37953
rect 29845 37950 30005 37953
rect 29634 37904 29638 37950
rect 29684 37904 29793 37950
rect 29845 37904 29959 37950
rect 29634 37901 29793 37904
rect 29845 37901 30005 37904
rect 30057 37950 30216 37953
rect 30057 37904 30121 37950
rect 30167 37904 30216 37950
rect 30057 37901 30216 37904
rect 30268 37950 30365 37953
rect 30268 37904 30284 37950
rect 30330 37904 30365 37950
rect 30268 37901 30365 37904
rect 29283 37861 30365 37901
rect 30583 37988 30637 38034
rect 30683 38028 30855 38034
rect 30901 38028 31040 38074
rect 33484 38070 33495 38492
rect 33541 38070 33552 38492
rect 34964 38517 35082 38574
rect 36438 38529 36554 38629
rect 37853 38624 38161 38629
rect 38658 38649 39723 38663
rect 34964 38485 36360 38517
rect 34228 38415 34718 38456
rect 34228 38398 34267 38415
rect 34319 38398 34447 38415
rect 34499 38398 34627 38415
rect 33671 38352 33684 38398
rect 33730 38352 33787 38398
rect 33833 38352 33890 38398
rect 33936 38352 33993 38398
rect 34039 38352 34096 38398
rect 34142 38352 34199 38398
rect 34245 38363 34267 38398
rect 34245 38352 34302 38363
rect 34348 38352 34405 38398
rect 34499 38363 34508 38398
rect 34451 38352 34508 38363
rect 34554 38352 34612 38398
rect 34679 38363 34718 38415
rect 34964 38439 35273 38485
rect 35523 38439 35580 38485
rect 35626 38439 35683 38485
rect 35729 38439 35786 38485
rect 35832 38439 35889 38485
rect 35935 38439 35992 38485
rect 36038 38439 36095 38485
rect 36141 38439 36198 38485
rect 36244 38439 36301 38485
rect 36347 38439 36360 38485
rect 34964 38395 36360 38439
rect 34658 38352 34718 38363
rect 34228 38323 34718 38352
rect 36438 38389 36475 38529
rect 36521 38389 36554 38529
rect 35294 38261 36266 38295
rect 36438 38286 36554 38389
rect 36640 38529 36773 38549
rect 36640 38490 36697 38529
rect 36640 38438 36678 38490
rect 36640 38389 36697 38438
rect 36743 38389 36773 38529
rect 38658 38527 38726 38649
rect 39809 38643 44918 38681
rect 48765 38663 48778 38709
rect 48824 38663 48881 38709
rect 48927 38663 48943 38709
rect 49030 38663 49087 38709
rect 49133 38663 49154 38709
rect 49236 38663 49293 38709
rect 49339 38663 49365 38709
rect 49442 38663 49499 38709
rect 49545 38663 49576 38709
rect 49852 38663 49877 38709
rect 54085 38727 54540 38760
rect 50481 38667 51657 38694
rect 39809 38597 43739 38643
rect 43785 38597 43906 38643
rect 43952 38597 44071 38643
rect 44117 38597 44236 38643
rect 44282 38622 44918 38643
rect 48905 38623 49877 38663
rect 50044 38657 51657 38667
rect 44282 38597 44812 38622
rect 39809 38594 44812 38597
rect 39809 38548 39844 38594
rect 39890 38592 44812 38594
rect 39890 38548 39994 38592
rect 39809 38540 39994 38548
rect 40046 38576 44812 38592
rect 44858 38576 44925 38622
rect 44971 38576 45038 38622
rect 45084 38576 45151 38622
rect 45197 38576 45264 38622
rect 45310 38576 45323 38622
rect 48557 38577 48687 38617
rect 40046 38561 44918 38576
rect 40046 38540 40085 38561
rect 39809 38537 40085 38540
rect 36924 38517 37685 38524
rect 36923 38485 37931 38517
rect 36841 38439 36854 38485
rect 36900 38483 36971 38485
rect 36900 38439 36961 38483
rect 37017 38439 37088 38485
rect 37134 38483 37206 38485
rect 37134 38439 37172 38483
rect 37252 38439 37324 38485
rect 37370 38483 37442 38485
rect 37370 38439 37384 38483
rect 36923 38431 36961 38439
rect 37013 38431 37172 38439
rect 37224 38431 37384 38439
rect 37436 38439 37442 38483
rect 37488 38483 37909 38485
rect 37488 38439 37595 38483
rect 37436 38431 37595 38439
rect 37647 38439 37909 38483
rect 37955 38439 38026 38485
rect 38072 38439 38143 38485
rect 38189 38439 38261 38485
rect 38307 38439 38379 38485
rect 38425 38439 38497 38485
rect 38543 38439 38556 38485
rect 37647 38431 37931 38439
rect 36923 38398 37931 38431
rect 36923 38397 37685 38398
rect 36924 38391 37685 38397
rect 36640 38366 36773 38389
rect 38658 38387 38669 38527
rect 38715 38387 38726 38527
rect 39014 38485 39323 38517
rect 39492 38485 39608 38517
rect 39008 38439 39021 38485
rect 39067 38439 39144 38485
rect 39190 38439 39267 38485
rect 39313 38439 39326 38485
rect 39492 38439 39641 38485
rect 39687 38439 39730 38485
rect 38658 38376 38726 38387
rect 36438 38261 36953 38286
rect 37439 38283 37931 38286
rect 37439 38261 38161 38283
rect 35260 38215 35273 38261
rect 35523 38255 35580 38261
rect 35523 38215 35543 38255
rect 35626 38215 35683 38261
rect 35729 38255 35786 38261
rect 35729 38215 35754 38255
rect 35832 38215 35889 38261
rect 35935 38255 35992 38261
rect 35935 38215 35965 38255
rect 36038 38215 36095 38261
rect 36141 38255 36198 38261
rect 36141 38215 36176 38255
rect 36244 38215 36301 38261
rect 36347 38215 36360 38261
rect 36438 38215 36854 38261
rect 36900 38215 36971 38261
rect 37017 38215 37088 38261
rect 37134 38215 37206 38261
rect 37252 38215 37324 38261
rect 37370 38215 37442 38261
rect 37488 38243 37909 38261
rect 37488 38215 37891 38243
rect 37955 38215 38026 38261
rect 38072 38243 38143 38261
rect 38123 38215 38143 38243
rect 38189 38215 38261 38261
rect 38307 38215 38379 38261
rect 38425 38215 38497 38261
rect 38543 38215 38556 38261
rect 33781 38174 34089 38209
rect 35294 38203 35332 38215
rect 35384 38203 35543 38215
rect 35595 38203 35754 38215
rect 35806 38203 35965 38215
rect 36017 38203 36176 38215
rect 36228 38203 36266 38215
rect 33671 38128 33684 38174
rect 33730 38128 33787 38174
rect 33833 38169 33890 38174
rect 33871 38128 33890 38169
rect 33936 38128 33993 38174
rect 34039 38169 34096 38174
rect 34051 38128 34096 38169
rect 34142 38128 34199 38174
rect 34245 38128 34302 38174
rect 34348 38128 34405 38174
rect 34451 38128 34508 38174
rect 34554 38128 34612 38174
rect 34658 38128 34671 38174
rect 35294 38163 36266 38203
rect 36438 38166 36953 38215
rect 37439 38191 37891 38215
rect 37943 38191 38071 38215
rect 38123 38191 38161 38215
rect 37439 38166 38161 38191
rect 37853 38150 38161 38166
rect 33781 38117 33819 38128
rect 33871 38117 33999 38128
rect 34051 38117 34089 38128
rect 33781 38076 34089 38117
rect 33484 38059 33552 38070
rect 30683 37994 31040 38028
rect 30683 37988 32842 37994
rect 30583 37953 32842 37988
rect 34247 37987 35008 37994
rect 30583 37901 30854 37953
rect 30906 37901 31065 37953
rect 31117 37901 31276 37953
rect 31328 37950 31486 37953
rect 31538 37950 31697 37953
rect 31749 37950 31909 37953
rect 31961 37950 32120 37953
rect 32172 37950 32330 37953
rect 32382 37950 32541 37953
rect 32593 37950 32752 37953
rect 32804 37950 32842 37953
rect 34246 37953 35008 37987
rect 34246 37950 34284 37953
rect 34336 37950 34495 37953
rect 34547 37950 34707 37953
rect 31328 37904 31349 37950
rect 33323 37904 33336 37950
rect 33671 37904 33684 37950
rect 33730 37904 33787 37950
rect 33833 37904 33890 37950
rect 33936 37904 33993 37950
rect 34039 37904 34096 37950
rect 34142 37904 34199 37950
rect 34245 37904 34284 37950
rect 34348 37904 34405 37950
rect 34451 37904 34495 37950
rect 34554 37904 34612 37950
rect 34658 37904 34707 37950
rect 31328 37901 31486 37904
rect 31538 37901 31697 37904
rect 31749 37901 31909 37904
rect 31961 37901 32120 37904
rect 32172 37901 32330 37904
rect 32382 37901 32541 37904
rect 32593 37901 32752 37904
rect 32804 37901 32842 37904
rect 30583 37866 32842 37901
rect 34246 37901 34284 37904
rect 34336 37901 34495 37904
rect 34547 37901 34707 37904
rect 34759 37901 34918 37953
rect 34970 37901 35008 37953
rect 34246 37867 35008 37901
rect 29544 37860 30306 37861
rect 27387 37744 29196 37820
rect 27387 37703 29116 37744
rect 27387 37657 28810 37703
rect 28856 37698 29116 37703
rect 29162 37698 29196 37744
rect 28856 37657 29196 37698
rect 27387 37581 29196 37657
rect 27387 37540 29116 37581
rect 27387 37494 28810 37540
rect 28856 37535 29116 37540
rect 29162 37535 29196 37581
rect 28856 37494 29196 37535
rect 27387 37417 29196 37494
rect 27387 37377 29116 37417
rect 27387 37331 28810 37377
rect 28856 37371 29116 37377
rect 29162 37371 29196 37417
rect 28856 37331 29196 37371
rect 27387 37254 29196 37331
rect 27387 37213 29116 37254
rect 27387 37167 28810 37213
rect 28856 37208 29116 37213
rect 29162 37208 29196 37254
rect 28856 37167 29196 37208
rect 27387 37053 29196 37167
rect 30583 37820 30637 37866
rect 30683 37860 32842 37866
rect 34247 37860 35008 37867
rect 35182 37987 36364 37994
rect 35182 37953 36958 37987
rect 35182 37901 35220 37953
rect 35272 37901 35430 37953
rect 35482 37901 35641 37953
rect 35693 37901 35853 37953
rect 35905 37901 36064 37953
rect 36116 37901 36274 37953
rect 36326 37950 36958 37953
rect 36326 37904 36489 37950
rect 36723 37904 36958 37950
rect 36326 37901 36958 37904
rect 35182 37867 36958 37901
rect 37946 37953 38842 37994
rect 37946 37950 38330 37953
rect 38382 37950 38541 37953
rect 37946 37904 37957 37950
rect 38473 37904 38541 37950
rect 37946 37901 38330 37904
rect 38382 37901 38541 37904
rect 38593 37901 38752 37953
rect 38804 37901 38842 37953
rect 35182 37860 36364 37867
rect 37946 37860 38842 37901
rect 39014 37953 39323 38439
rect 39014 37901 39052 37953
rect 39104 37950 39232 37953
rect 39108 37904 39220 37950
rect 39104 37901 39232 37904
rect 39284 37901 39323 37953
rect 30683 37826 31040 37860
rect 30683 37820 30855 37826
rect 30583 37780 30855 37820
rect 30901 37780 31040 37826
rect 30583 37703 31040 37780
rect 33484 37784 33552 37795
rect 33019 37729 33327 37770
rect 33019 37726 33057 37729
rect 33109 37726 33237 37729
rect 33289 37726 33327 37729
rect 30583 37657 30637 37703
rect 30683 37662 31040 37703
rect 31336 37680 31349 37726
rect 33323 37680 33336 37726
rect 30683 37657 30855 37662
rect 30583 37616 30855 37657
rect 30901 37616 31040 37662
rect 33019 37677 33057 37680
rect 33109 37677 33237 37680
rect 33289 37677 33327 37680
rect 33019 37637 33327 37677
rect 30583 37540 31040 37616
rect 30583 37494 30637 37540
rect 30683 37524 31040 37540
rect 30683 37502 31493 37524
rect 30683 37499 31349 37502
rect 30683 37494 30855 37499
rect 30583 37453 30855 37494
rect 30901 37456 31349 37499
rect 33323 37456 33336 37502
rect 30901 37453 31493 37456
rect 30583 37405 31493 37453
rect 30583 37377 31040 37405
rect 30583 37331 30637 37377
rect 30683 37336 31040 37377
rect 30683 37331 30855 37336
rect 30583 37290 30855 37331
rect 30901 37290 31040 37336
rect 33484 37362 33495 37784
rect 33541 37362 33552 37784
rect 33781 37737 34089 37778
rect 33781 37726 33819 37737
rect 33871 37726 33999 37737
rect 34051 37726 34089 37737
rect 33671 37680 33684 37726
rect 33730 37680 33787 37726
rect 33871 37685 33890 37726
rect 33833 37680 33890 37685
rect 33936 37680 33993 37726
rect 34051 37685 34096 37726
rect 34039 37680 34096 37685
rect 34142 37680 34199 37726
rect 34245 37680 34302 37726
rect 34348 37680 34405 37726
rect 34451 37680 34508 37726
rect 34554 37680 34612 37726
rect 34658 37680 34671 37726
rect 33781 37645 34089 37680
rect 35294 37651 36266 37691
rect 37853 37688 38161 37704
rect 35294 37639 35332 37651
rect 35384 37639 35543 37651
rect 35595 37639 35754 37651
rect 35806 37639 35965 37651
rect 36017 37639 36176 37651
rect 36228 37639 36266 37651
rect 36438 37639 36953 37688
rect 37439 37663 38161 37688
rect 37439 37639 37891 37663
rect 37943 37639 38071 37663
rect 38123 37639 38161 37663
rect 35260 37593 35273 37639
rect 35523 37599 35543 37639
rect 35523 37593 35580 37599
rect 35626 37593 35683 37639
rect 35729 37599 35754 37639
rect 35729 37593 35786 37599
rect 35832 37593 35889 37639
rect 35935 37599 35965 37639
rect 35935 37593 35992 37599
rect 36038 37593 36095 37639
rect 36141 37599 36176 37639
rect 36141 37593 36198 37599
rect 36244 37593 36301 37639
rect 36347 37593 36360 37639
rect 36438 37593 36854 37639
rect 36900 37593 36971 37639
rect 37017 37593 37088 37639
rect 37134 37593 37206 37639
rect 37252 37593 37324 37639
rect 37370 37593 37442 37639
rect 37488 37611 37891 37639
rect 37488 37593 37909 37611
rect 37955 37593 38026 37639
rect 38123 37611 38143 37639
rect 38072 37593 38143 37611
rect 38189 37593 38261 37639
rect 38307 37593 38379 37639
rect 38425 37593 38497 37639
rect 38543 37593 38556 37639
rect 35294 37559 36266 37593
rect 36438 37568 36953 37593
rect 37439 37571 38161 37593
rect 37439 37568 37931 37571
rect 34228 37502 34718 37531
rect 33671 37456 33684 37502
rect 33730 37456 33787 37502
rect 33833 37456 33890 37502
rect 33936 37456 33993 37502
rect 34039 37456 34096 37502
rect 34142 37456 34199 37502
rect 34245 37491 34302 37502
rect 34245 37456 34267 37491
rect 34348 37456 34405 37502
rect 34451 37491 34508 37502
rect 34499 37456 34508 37491
rect 34554 37456 34612 37502
rect 34658 37491 34718 37502
rect 34228 37439 34267 37456
rect 34319 37439 34447 37456
rect 34499 37439 34627 37456
rect 34679 37439 34718 37491
rect 36438 37465 36554 37568
rect 34228 37398 34718 37439
rect 34964 37415 36360 37459
rect 30583 37213 31040 37290
rect 33019 37281 33327 37322
rect 33019 37278 33057 37281
rect 33109 37278 33237 37281
rect 33289 37278 33327 37281
rect 33484 37280 33552 37362
rect 34964 37369 35273 37415
rect 35523 37369 35580 37415
rect 35626 37369 35683 37415
rect 35729 37369 35786 37415
rect 35832 37369 35889 37415
rect 35935 37369 35992 37415
rect 36038 37369 36095 37415
rect 36141 37369 36198 37415
rect 36244 37369 36301 37415
rect 36347 37369 36360 37415
rect 34964 37337 36360 37369
rect 34964 37280 35082 37337
rect 31336 37232 31349 37278
rect 33323 37232 33336 37278
rect 33484 37243 35082 37280
rect 30583 37167 30637 37213
rect 30683 37173 31040 37213
rect 33019 37229 33057 37232
rect 33109 37229 33237 37232
rect 33289 37229 33327 37232
rect 33019 37189 33327 37229
rect 33484 37197 33816 37243
rect 33862 37197 34002 37243
rect 34048 37197 34189 37243
rect 34235 37197 34376 37243
rect 34422 37197 34562 37243
rect 34608 37197 35082 37243
rect 36438 37325 36475 37465
rect 36521 37325 36554 37465
rect 33484 37189 35082 37197
rect 35294 37191 36266 37231
rect 36438 37225 36554 37325
rect 36640 37465 36773 37488
rect 36640 37416 36697 37465
rect 36640 37364 36678 37416
rect 36640 37325 36697 37364
rect 36743 37325 36773 37465
rect 38658 37467 38726 37478
rect 36924 37457 37685 37463
rect 36923 37456 37685 37457
rect 36923 37423 37931 37456
rect 36923 37415 36961 37423
rect 37013 37415 37172 37423
rect 37224 37415 37384 37423
rect 36841 37369 36854 37415
rect 36900 37371 36961 37415
rect 36900 37369 36971 37371
rect 37017 37369 37088 37415
rect 37134 37371 37172 37415
rect 37134 37369 37206 37371
rect 37252 37369 37324 37415
rect 37370 37371 37384 37415
rect 37436 37415 37595 37423
rect 37436 37371 37442 37415
rect 37370 37369 37442 37371
rect 37488 37371 37595 37415
rect 37647 37415 37931 37423
rect 37647 37371 37909 37415
rect 37488 37369 37909 37371
rect 37955 37369 38026 37415
rect 38072 37369 38143 37415
rect 38189 37369 38261 37415
rect 38307 37369 38379 37415
rect 38425 37369 38497 37415
rect 38543 37369 38556 37415
rect 36923 37337 37931 37369
rect 36924 37330 37685 37337
rect 36640 37305 36773 37325
rect 38658 37327 38669 37467
rect 38715 37327 38726 37467
rect 39014 37415 39323 37901
rect 39492 37987 39608 38439
rect 39923 38406 40085 38537
rect 39923 38354 39994 38406
rect 40046 38354 40085 38406
rect 39923 38314 40085 38354
rect 39737 38218 39865 38231
rect 39737 38191 39866 38218
rect 39737 38174 39775 38191
rect 39827 38174 39866 38191
rect 39727 38128 39740 38174
rect 39827 38139 39862 38174
rect 39786 38128 39862 38139
rect 39908 38128 39985 38174
rect 40031 38128 40108 38174
rect 40154 38128 40167 38174
rect 40246 38163 40362 38561
rect 42229 38422 44509 38463
rect 42229 38370 43445 38422
rect 43497 38370 44509 38422
rect 42229 38330 44509 38370
rect 44341 38286 44509 38330
rect 44341 38240 44358 38286
rect 44498 38240 44509 38286
rect 39737 38099 39866 38128
rect 40246 38117 40281 38163
rect 40327 38117 40362 38163
rect 40246 38080 40362 38117
rect 40718 38191 43524 38232
rect 44341 38229 44509 38240
rect 40718 38139 41935 38191
rect 41987 38139 43524 38191
rect 40718 38098 43524 38139
rect 44605 38174 44721 38561
rect 45400 38531 48379 38572
rect 45400 38517 47486 38531
rect 45400 38471 45464 38517
rect 45604 38479 47486 38517
rect 47538 38479 48379 38531
rect 45604 38471 48379 38479
rect 44901 38415 45241 38456
rect 45400 38438 48379 38471
rect 48557 38525 48596 38577
rect 48648 38525 48687 38577
rect 48557 38502 48687 38525
rect 50044 38611 50516 38657
rect 50562 38611 50703 38657
rect 50749 38611 50890 38657
rect 50936 38611 51076 38657
rect 51122 38611 51263 38657
rect 51309 38611 51657 38657
rect 51797 38647 52105 38687
rect 51797 38622 51835 38647
rect 51887 38622 52015 38647
rect 52067 38622 52105 38647
rect 54085 38681 54223 38727
rect 54269 38687 54540 38727
rect 54269 38681 54440 38687
rect 54085 38641 54440 38681
rect 54486 38641 54540 38687
rect 50044 38574 51657 38611
rect 51789 38576 51802 38622
rect 53776 38576 53789 38622
rect 50044 38517 50160 38574
rect 44901 38398 44939 38415
rect 44991 38398 45151 38415
rect 45203 38398 45241 38415
rect 44799 38352 44812 38398
rect 44858 38352 44925 38398
rect 44991 38363 45038 38398
rect 44971 38352 45038 38363
rect 45084 38352 45151 38398
rect 45203 38363 45264 38398
rect 45197 38352 45264 38363
rect 45310 38352 45323 38398
rect 48557 38362 48622 38502
rect 48668 38362 48687 38502
rect 49820 38485 50160 38517
rect 48765 38439 48778 38485
rect 48824 38439 48881 38485
rect 48927 38439 48984 38485
rect 49030 38439 49087 38485
rect 49133 38439 49190 38485
rect 49236 38439 49293 38485
rect 49339 38439 49396 38485
rect 49442 38439 49499 38485
rect 49545 38439 49602 38485
rect 49852 38439 50160 38485
rect 51589 38522 51657 38574
rect 51797 38554 52105 38576
rect 49820 38398 50160 38439
rect 50262 38415 50812 38456
rect 48557 38359 48687 38362
rect 44901 38323 45241 38352
rect 48557 38307 48596 38359
rect 48648 38307 48687 38359
rect 50262 38363 50300 38415
rect 50352 38398 50511 38415
rect 50563 38398 50722 38415
rect 50352 38363 50467 38398
rect 50563 38363 50571 38398
rect 50262 38352 50467 38363
rect 50513 38352 50571 38363
rect 50617 38352 50674 38398
rect 50720 38363 50722 38398
rect 50774 38398 50812 38415
rect 50774 38363 50777 38398
rect 50720 38352 50777 38363
rect 50823 38352 50880 38398
rect 50926 38352 50983 38398
rect 51029 38352 51086 38398
rect 51132 38352 51189 38398
rect 51235 38352 51292 38398
rect 51338 38352 51395 38398
rect 51441 38352 51454 38398
rect 50262 38323 50812 38352
rect 48557 38266 48687 38307
rect 48905 38261 49877 38292
rect 48765 38215 48778 38261
rect 48824 38215 48881 38261
rect 48927 38252 48984 38261
rect 48927 38215 48943 38252
rect 49030 38215 49087 38261
rect 49133 38252 49190 38261
rect 49133 38215 49154 38252
rect 49236 38215 49293 38261
rect 49339 38252 49396 38261
rect 49339 38215 49365 38252
rect 49442 38215 49499 38261
rect 49545 38252 49602 38261
rect 49545 38215 49576 38252
rect 49852 38215 49877 38261
rect 48905 38200 48943 38215
rect 48995 38200 49154 38215
rect 49206 38200 49365 38215
rect 49417 38200 49576 38215
rect 49628 38200 49787 38215
rect 49839 38200 49877 38215
rect 44605 38128 44812 38174
rect 44858 38128 44925 38174
rect 44971 38128 45038 38174
rect 45084 38128 45151 38174
rect 45197 38128 45264 38174
rect 45310 38128 45323 38174
rect 48905 38160 49877 38200
rect 51035 38177 51343 38217
rect 51035 38174 51073 38177
rect 51125 38174 51253 38177
rect 51305 38174 51343 38177
rect 43362 38091 43524 38098
rect 43362 38045 43373 38091
rect 43513 38045 43524 38091
rect 43362 38034 43524 38045
rect 45584 38114 48546 38150
rect 50454 38128 50467 38174
rect 50513 38128 50571 38174
rect 50617 38128 50674 38174
rect 50720 38128 50777 38174
rect 50823 38128 50880 38174
rect 50926 38128 50983 38174
rect 51029 38128 51073 38174
rect 51132 38128 51189 38174
rect 51235 38128 51253 38174
rect 51338 38128 51395 38174
rect 51441 38128 51454 38174
rect 45584 38068 45619 38114
rect 45665 38068 45777 38114
rect 45823 38068 45935 38114
rect 45981 38068 46093 38114
rect 46139 38068 46251 38114
rect 46297 38068 46409 38114
rect 46455 38068 46568 38114
rect 46614 38068 46726 38114
rect 46772 38068 46884 38114
rect 46930 38068 47042 38114
rect 47088 38068 47200 38114
rect 47246 38068 47358 38114
rect 47404 38068 47516 38114
rect 47562 38068 47675 38114
rect 47721 38068 47833 38114
rect 47879 38068 47991 38114
rect 48037 38068 48149 38114
rect 48195 38068 48307 38114
rect 48353 38068 48465 38114
rect 48511 38068 48546 38114
rect 51035 38125 51073 38128
rect 51125 38125 51253 38128
rect 51305 38125 51343 38128
rect 51035 38084 51343 38125
rect 51589 38100 51600 38522
rect 51646 38100 51657 38522
rect 54085 38523 54540 38641
rect 54085 38477 54440 38523
rect 54486 38477 54540 38523
rect 54085 38449 54540 38477
rect 53585 38398 54540 38449
rect 51789 38352 51802 38398
rect 53776 38360 54540 38398
rect 53776 38352 54440 38360
rect 53585 38330 54440 38352
rect 54085 38314 54440 38330
rect 54486 38314 54540 38360
rect 54085 38238 54540 38314
rect 51797 38184 52105 38224
rect 51797 38174 51835 38184
rect 51887 38174 52015 38184
rect 52067 38174 52105 38184
rect 54085 38192 54223 38238
rect 54269 38197 54540 38238
rect 54269 38192 54440 38197
rect 51789 38128 51802 38174
rect 53776 38128 53789 38174
rect 54085 38151 54440 38192
rect 54486 38151 54540 38197
rect 51589 38089 51657 38100
rect 51797 38091 52105 38128
rect 40215 37987 40523 37994
rect 40788 37987 42986 38001
rect 43753 37987 44514 37994
rect 39492 37964 42986 37987
rect 43704 37964 44514 37987
rect 39492 37953 44514 37964
rect 39492 37950 40253 37953
rect 39492 37904 39740 37950
rect 39786 37904 39862 37950
rect 39908 37904 39985 37950
rect 40031 37904 40108 37950
rect 40154 37904 40253 37950
rect 39492 37901 40253 37904
rect 40305 37901 40433 37953
rect 40485 37950 43790 37953
rect 40485 37904 40836 37950
rect 40882 37904 40994 37950
rect 41040 37904 41152 37950
rect 41198 37904 41310 37950
rect 41356 37904 41469 37950
rect 41515 37904 41627 37950
rect 41673 37904 41785 37950
rect 41831 37904 41943 37950
rect 41989 37904 42101 37950
rect 42147 37904 42259 37950
rect 42305 37904 42418 37950
rect 42464 37904 42576 37950
rect 42622 37904 42734 37950
rect 42780 37904 42892 37950
rect 42938 37904 43739 37950
rect 43785 37904 43790 37950
rect 40485 37901 43790 37904
rect 43842 37950 44001 37953
rect 43842 37904 43906 37950
rect 43952 37904 44001 37950
rect 43842 37901 44001 37904
rect 44053 37950 44213 37953
rect 44265 37950 44424 37953
rect 44053 37904 44071 37950
rect 44117 37904 44213 37950
rect 44282 37904 44424 37950
rect 44053 37901 44213 37904
rect 44265 37901 44424 37904
rect 44476 37901 44514 37953
rect 39492 37890 44514 37901
rect 39492 37867 42986 37890
rect 43704 37867 44514 37890
rect 39492 37415 39608 37867
rect 40215 37860 40523 37867
rect 40788 37853 42986 37867
rect 43753 37860 44514 37867
rect 44796 37987 45346 37994
rect 45584 37987 48546 38068
rect 54085 38074 54540 38151
rect 54085 38028 54223 38074
rect 54269 38034 54540 38074
rect 54269 38028 54440 38034
rect 54085 37994 54440 38028
rect 48800 37987 49982 37994
rect 50308 37987 50859 37994
rect 44796 37953 49982 37987
rect 44796 37950 44834 37953
rect 44886 37950 45045 37953
rect 45097 37950 45256 37953
rect 45308 37950 48838 37953
rect 44796 37904 44812 37950
rect 44886 37904 44925 37950
rect 44971 37904 45038 37950
rect 45097 37904 45151 37950
rect 45197 37904 45256 37950
rect 45310 37904 45619 37950
rect 45665 37904 45777 37950
rect 45823 37904 45935 37950
rect 45981 37904 46093 37950
rect 46139 37904 46251 37950
rect 46297 37904 46409 37950
rect 46455 37904 46568 37950
rect 46614 37904 46726 37950
rect 46772 37904 46884 37950
rect 46930 37904 47042 37950
rect 47088 37904 47200 37950
rect 47246 37904 47358 37950
rect 47404 37904 47516 37950
rect 47562 37904 47675 37950
rect 47721 37904 47833 37950
rect 47879 37904 47991 37950
rect 48037 37904 48149 37950
rect 48195 37904 48307 37950
rect 48353 37904 48465 37950
rect 48511 37904 48838 37950
rect 44796 37901 44834 37904
rect 44886 37901 45045 37904
rect 45097 37901 45256 37904
rect 45308 37901 48838 37904
rect 48890 37901 49048 37953
rect 49100 37901 49259 37953
rect 49311 37901 49471 37953
rect 49523 37901 49682 37953
rect 49734 37901 49892 37953
rect 49944 37901 49982 37953
rect 44796 37867 49982 37901
rect 50307 37953 50859 37987
rect 50307 37901 50346 37953
rect 50398 37950 50557 37953
rect 50609 37950 50768 37953
rect 50820 37950 50859 37953
rect 52278 37988 54440 37994
rect 54486 37988 54540 38034
rect 55927 38687 57736 38801
rect 55927 38644 56267 38687
rect 55927 38598 55961 38644
rect 56007 38641 56267 38644
rect 56313 38641 57736 38687
rect 56007 38598 57736 38641
rect 55927 38523 57736 38598
rect 55927 38481 56267 38523
rect 55927 38435 55961 38481
rect 56007 38477 56267 38481
rect 56313 38477 57736 38523
rect 56007 38435 57736 38477
rect 55927 38360 57736 38435
rect 55927 38317 56267 38360
rect 55927 38271 55961 38317
rect 56007 38314 56267 38317
rect 56313 38314 57736 38360
rect 56007 38271 57736 38314
rect 55927 38197 57736 38271
rect 55927 38154 56267 38197
rect 55927 38108 55961 38154
rect 56007 38151 56267 38154
rect 56313 38151 57736 38197
rect 56007 38108 57736 38151
rect 55927 38034 57736 38108
rect 52278 37953 54540 37988
rect 52278 37950 52316 37953
rect 52368 37950 52527 37953
rect 52579 37950 52738 37953
rect 52790 37950 52948 37953
rect 53000 37950 53159 37953
rect 53211 37950 53371 37953
rect 53423 37950 53582 37953
rect 53634 37950 53792 37953
rect 50398 37904 50467 37950
rect 50513 37904 50557 37950
rect 50617 37904 50674 37950
rect 50720 37904 50768 37950
rect 50823 37904 50880 37950
rect 50926 37904 50983 37950
rect 51029 37904 51086 37950
rect 51132 37904 51189 37950
rect 51235 37904 51292 37950
rect 51338 37904 51395 37950
rect 51441 37904 51454 37950
rect 51789 37904 51802 37950
rect 53776 37904 53792 37950
rect 50398 37901 50557 37904
rect 50609 37901 50768 37904
rect 50820 37901 50859 37904
rect 50307 37867 50859 37901
rect 44796 37860 45346 37867
rect 43362 37809 43524 37820
rect 39737 37726 39866 37755
rect 40246 37737 40362 37774
rect 43362 37763 43373 37809
rect 43513 37763 43524 37809
rect 43362 37756 43524 37763
rect 39727 37680 39740 37726
rect 39786 37715 39862 37726
rect 39827 37680 39862 37715
rect 39908 37680 39985 37726
rect 40031 37680 40108 37726
rect 40154 37680 40167 37726
rect 40246 37691 40281 37737
rect 40327 37691 40362 37737
rect 39737 37663 39775 37680
rect 39827 37663 39866 37680
rect 39737 37636 39866 37663
rect 39737 37623 39865 37636
rect 39923 37500 40085 37540
rect 39923 37448 39994 37500
rect 40046 37448 40085 37500
rect 39008 37369 39021 37415
rect 39067 37369 39144 37415
rect 39190 37369 39267 37415
rect 39313 37369 39326 37415
rect 39492 37369 39641 37415
rect 39687 37369 39730 37415
rect 39014 37337 39323 37369
rect 39492 37337 39608 37369
rect 37853 37225 38161 37230
rect 36438 37191 36953 37225
rect 37439 37191 38161 37225
rect 38658 37205 38726 37327
rect 39923 37317 40085 37448
rect 39809 37314 40085 37317
rect 39809 37306 39994 37314
rect 39809 37260 39844 37306
rect 39890 37262 39994 37306
rect 40046 37293 40085 37314
rect 40246 37293 40362 37691
rect 40718 37715 43524 37756
rect 45584 37786 48546 37867
rect 48800 37860 49982 37867
rect 50308 37860 50859 37867
rect 52278 37901 52316 37904
rect 52368 37901 52527 37904
rect 52579 37901 52738 37904
rect 52790 37901 52948 37904
rect 53000 37901 53159 37904
rect 53211 37901 53371 37904
rect 53423 37901 53582 37904
rect 53634 37901 53792 37904
rect 53844 37901 54003 37953
rect 54055 37901 54214 37953
rect 54266 37901 54540 37953
rect 52278 37866 54540 37901
rect 52278 37860 54440 37866
rect 45584 37740 45619 37786
rect 45665 37740 45777 37786
rect 45823 37740 45935 37786
rect 45981 37740 46093 37786
rect 46139 37740 46251 37786
rect 46297 37740 46409 37786
rect 46455 37740 46568 37786
rect 46614 37740 46726 37786
rect 46772 37740 46884 37786
rect 46930 37740 47042 37786
rect 47088 37740 47200 37786
rect 47246 37740 47358 37786
rect 47404 37740 47516 37786
rect 47562 37740 47675 37786
rect 47721 37740 47833 37786
rect 47879 37740 47991 37786
rect 48037 37740 48149 37786
rect 48195 37740 48307 37786
rect 48353 37740 48465 37786
rect 48511 37740 48546 37786
rect 54085 37826 54440 37860
rect 54085 37780 54223 37826
rect 54269 37820 54440 37826
rect 54486 37820 54540 37866
rect 54758 37953 55840 37994
rect 54758 37950 54855 37953
rect 54758 37904 54793 37950
rect 54839 37904 54855 37950
rect 54758 37901 54855 37904
rect 54907 37950 55066 37953
rect 54907 37904 54956 37950
rect 55002 37904 55066 37950
rect 54907 37901 55066 37904
rect 55118 37950 55278 37953
rect 55330 37950 55489 37953
rect 55164 37904 55278 37950
rect 55330 37904 55439 37950
rect 55485 37904 55489 37950
rect 55118 37901 55278 37904
rect 55330 37901 55489 37904
rect 55541 37950 55840 37953
rect 55541 37904 55599 37950
rect 55645 37904 55760 37950
rect 55806 37904 55840 37950
rect 55541 37901 55840 37904
rect 54758 37861 55840 37901
rect 55927 37988 56267 38034
rect 56313 37988 57736 38034
rect 55927 37866 57736 37988
rect 54817 37860 55579 37861
rect 54269 37780 54540 37820
rect 40718 37663 41935 37715
rect 41987 37663 43524 37715
rect 40718 37622 43524 37663
rect 44605 37680 44812 37726
rect 44858 37680 44925 37726
rect 44971 37680 45038 37726
rect 45084 37680 45151 37726
rect 45197 37680 45264 37726
rect 45310 37680 45323 37726
rect 45584 37704 48546 37740
rect 51035 37729 51343 37770
rect 51035 37726 51073 37729
rect 51125 37726 51253 37729
rect 51305 37726 51343 37729
rect 51589 37754 51657 37765
rect 44341 37614 44509 37625
rect 44341 37568 44358 37614
rect 44498 37568 44509 37614
rect 44341 37524 44509 37568
rect 42229 37484 44509 37524
rect 42229 37432 43445 37484
rect 43497 37432 44509 37484
rect 42229 37391 44509 37432
rect 44605 37293 44721 37680
rect 48905 37654 49877 37694
rect 50454 37680 50467 37726
rect 50513 37680 50571 37726
rect 50617 37680 50674 37726
rect 50720 37680 50777 37726
rect 50823 37680 50880 37726
rect 50926 37680 50983 37726
rect 51029 37680 51073 37726
rect 51132 37680 51189 37726
rect 51235 37680 51253 37726
rect 51338 37680 51395 37726
rect 51441 37680 51454 37726
rect 48905 37639 48943 37654
rect 48995 37639 49154 37654
rect 49206 37639 49365 37654
rect 49417 37639 49576 37654
rect 49628 37639 49787 37654
rect 49839 37639 49877 37654
rect 48765 37593 48778 37639
rect 48824 37593 48881 37639
rect 48927 37602 48943 37639
rect 48927 37593 48984 37602
rect 49030 37593 49087 37639
rect 49133 37602 49154 37639
rect 49133 37593 49190 37602
rect 49236 37593 49293 37639
rect 49339 37602 49365 37639
rect 49339 37593 49396 37602
rect 49442 37593 49499 37639
rect 49545 37602 49576 37639
rect 49545 37593 49602 37602
rect 49852 37593 49877 37639
rect 51035 37677 51073 37680
rect 51125 37677 51253 37680
rect 51305 37677 51343 37680
rect 51035 37637 51343 37677
rect 48557 37547 48687 37588
rect 48905 37562 49877 37593
rect 44901 37502 45241 37531
rect 44799 37456 44812 37502
rect 44858 37456 44925 37502
rect 44971 37491 45038 37502
rect 44991 37456 45038 37491
rect 45084 37456 45151 37502
rect 45197 37491 45264 37502
rect 45203 37456 45264 37491
rect 45310 37456 45323 37502
rect 48557 37495 48596 37547
rect 48648 37495 48687 37547
rect 48557 37492 48687 37495
rect 44901 37439 44939 37456
rect 44991 37439 45151 37456
rect 45203 37439 45241 37456
rect 44901 37398 45241 37439
rect 45400 37383 48379 37416
rect 45400 37337 45464 37383
rect 45604 37375 48379 37383
rect 45604 37337 47864 37375
rect 45400 37323 47864 37337
rect 47916 37323 48379 37375
rect 40046 37278 44918 37293
rect 45400 37282 48379 37323
rect 48557 37352 48622 37492
rect 48668 37352 48687 37492
rect 50262 37502 50812 37531
rect 50262 37491 50467 37502
rect 50513 37491 50571 37502
rect 49820 37415 50160 37456
rect 48765 37369 48778 37415
rect 48824 37369 48881 37415
rect 48927 37369 48984 37415
rect 49030 37369 49087 37415
rect 49133 37369 49190 37415
rect 49236 37369 49293 37415
rect 49339 37369 49396 37415
rect 49442 37369 49499 37415
rect 49545 37369 49602 37415
rect 49852 37369 50160 37415
rect 50262 37439 50300 37491
rect 50352 37456 50467 37491
rect 50563 37456 50571 37491
rect 50617 37456 50674 37502
rect 50720 37491 50777 37502
rect 50720 37456 50722 37491
rect 50352 37439 50511 37456
rect 50563 37439 50722 37456
rect 50774 37456 50777 37491
rect 50823 37456 50880 37502
rect 50926 37456 50983 37502
rect 51029 37456 51086 37502
rect 51132 37456 51189 37502
rect 51235 37456 51292 37502
rect 51338 37456 51395 37502
rect 51441 37456 51454 37502
rect 50774 37439 50812 37456
rect 50262 37398 50812 37439
rect 48557 37329 48687 37352
rect 49820 37337 50160 37369
rect 40046 37262 44812 37278
rect 39890 37260 44812 37262
rect 39809 37257 44812 37260
rect 39809 37211 43739 37257
rect 43785 37211 43906 37257
rect 43952 37211 44071 37257
rect 44117 37211 44236 37257
rect 44282 37232 44812 37257
rect 44858 37232 44925 37278
rect 44971 37232 45038 37278
rect 45084 37232 45151 37278
rect 45197 37232 45264 37278
rect 45310 37232 45323 37278
rect 48557 37277 48596 37329
rect 48648 37277 48687 37329
rect 48557 37237 48687 37277
rect 50044 37280 50160 37337
rect 51589 37332 51600 37754
rect 51646 37332 51657 37754
rect 51797 37726 52105 37763
rect 51789 37680 51802 37726
rect 53776 37680 53789 37726
rect 54085 37703 54540 37780
rect 51797 37670 51835 37680
rect 51887 37670 52015 37680
rect 52067 37670 52105 37680
rect 51797 37630 52105 37670
rect 54085 37662 54440 37703
rect 54085 37616 54223 37662
rect 54269 37657 54440 37662
rect 54486 37657 54540 37703
rect 54269 37616 54540 37657
rect 54085 37540 54540 37616
rect 54085 37524 54440 37540
rect 53585 37502 54440 37524
rect 51789 37456 51802 37502
rect 53776 37494 54440 37502
rect 54486 37494 54540 37540
rect 53776 37456 54540 37494
rect 53585 37405 54540 37456
rect 51589 37280 51657 37332
rect 54085 37377 54540 37405
rect 54085 37331 54440 37377
rect 54486 37331 54540 37377
rect 50044 37243 51657 37280
rect 51797 37278 52105 37300
rect 44282 37211 44918 37232
rect 38658 37191 39723 37205
rect 30683 37167 30855 37173
rect 30583 37127 30855 37167
rect 30901 37127 31040 37173
rect 33484 37160 34643 37189
rect 35260 37145 35273 37191
rect 35523 37145 35543 37191
rect 35626 37145 35683 37191
rect 35729 37145 35754 37191
rect 35832 37145 35889 37191
rect 35935 37145 35965 37191
rect 36038 37145 36095 37191
rect 36141 37145 36176 37191
rect 36244 37145 36301 37191
rect 36347 37145 36360 37191
rect 36438 37145 36854 37191
rect 36900 37145 36971 37191
rect 37017 37145 37088 37191
rect 37134 37145 37206 37191
rect 37252 37145 37324 37191
rect 37370 37145 37442 37191
rect 37488 37189 37909 37191
rect 37488 37145 37891 37189
rect 37955 37145 38026 37191
rect 38072 37189 38143 37191
rect 38123 37145 38143 37189
rect 38189 37145 38261 37191
rect 38307 37145 38379 37191
rect 38425 37145 38497 37191
rect 38543 37145 38556 37191
rect 38658 37145 39021 37191
rect 39067 37145 39144 37191
rect 39190 37145 39267 37191
rect 39313 37145 39641 37191
rect 39687 37145 39730 37191
rect 39809 37173 44918 37211
rect 48905 37191 49877 37231
rect 48765 37145 48778 37191
rect 48824 37145 48881 37191
rect 48927 37145 48943 37191
rect 49030 37145 49087 37191
rect 49133 37145 49154 37191
rect 49236 37145 49293 37191
rect 49339 37145 49365 37191
rect 49442 37145 49499 37191
rect 49545 37145 49576 37191
rect 49852 37145 49877 37191
rect 50044 37197 50516 37243
rect 50562 37197 50703 37243
rect 50749 37197 50890 37243
rect 50936 37197 51076 37243
rect 51122 37197 51263 37243
rect 51309 37197 51657 37243
rect 51789 37232 51802 37278
rect 53776 37232 53789 37278
rect 50044 37187 51657 37197
rect 50481 37160 51657 37187
rect 51797 37207 51835 37232
rect 51887 37207 52015 37232
rect 52067 37207 52105 37232
rect 51797 37167 52105 37207
rect 54085 37213 54540 37331
rect 54085 37173 54440 37213
rect 30583 37094 31040 37127
rect 35294 37139 35332 37145
rect 35384 37139 35543 37145
rect 35595 37139 35754 37145
rect 35806 37139 35965 37145
rect 36017 37139 36176 37145
rect 36228 37139 36266 37145
rect 34870 37094 35025 37101
rect 35294 37099 36266 37139
rect 36438 37105 36953 37145
rect 37439 37137 37891 37145
rect 37943 37137 38071 37145
rect 38123 37137 38161 37145
rect 37439 37105 38161 37137
rect 37853 37097 38161 37105
rect 27387 37001 27790 37053
rect 27842 37001 28001 37053
rect 28053 37001 28212 37053
rect 28264 37001 28423 37053
rect 28475 37001 28634 37053
rect 28686 37050 28845 37053
rect 28686 37004 28810 37050
rect 28686 37001 28845 37004
rect 28897 37001 29056 37053
rect 29108 37001 29196 37053
rect 27387 36887 29196 37001
rect 29283 37053 30365 37094
rect 29283 37050 29582 37053
rect 29283 37004 29317 37050
rect 29363 37004 29478 37050
rect 29524 37004 29582 37050
rect 29283 37001 29582 37004
rect 29634 37050 29793 37053
rect 29845 37050 30005 37053
rect 29634 37004 29638 37050
rect 29684 37004 29793 37050
rect 29845 37004 29959 37050
rect 29634 37001 29793 37004
rect 29845 37001 30005 37004
rect 30057 37050 30216 37053
rect 30057 37004 30121 37050
rect 30167 37004 30216 37050
rect 30057 37001 30216 37004
rect 30268 37050 30365 37053
rect 30268 37004 30284 37050
rect 30330 37004 30365 37050
rect 30268 37001 30365 37004
rect 29283 36961 30365 37001
rect 30583 37053 32842 37094
rect 30583 37050 30854 37053
rect 30583 37004 30637 37050
rect 30683 37004 30854 37050
rect 30583 37001 30854 37004
rect 30906 37001 31065 37053
rect 31117 37001 31276 37053
rect 31328 37001 31486 37053
rect 31538 37001 31697 37053
rect 31749 37001 31909 37053
rect 31961 37001 32120 37053
rect 32172 37001 32330 37053
rect 32382 37001 32541 37053
rect 32593 37001 32752 37053
rect 32804 37001 32842 37053
rect 29544 36960 30306 36961
rect 30583 36960 32842 37001
rect 34717 37053 35025 37094
rect 38658 37085 39723 37145
rect 48905 37139 48943 37145
rect 48995 37139 49154 37145
rect 49206 37139 49365 37145
rect 49417 37139 49576 37145
rect 49628 37139 49787 37145
rect 49839 37139 49877 37145
rect 48905 37099 49877 37139
rect 54085 37127 54223 37173
rect 54269 37167 54440 37173
rect 54486 37167 54540 37213
rect 54269 37127 54540 37167
rect 50099 37094 50255 37101
rect 54085 37094 54540 37127
rect 55927 37820 56267 37866
rect 56313 37820 57736 37866
rect 55927 37744 57736 37820
rect 55927 37698 55961 37744
rect 56007 37703 57736 37744
rect 56007 37698 56267 37703
rect 55927 37657 56267 37698
rect 56313 37657 57736 37703
rect 55927 37581 57736 37657
rect 55927 37535 55961 37581
rect 56007 37540 57736 37581
rect 56007 37535 56267 37540
rect 55927 37494 56267 37535
rect 56313 37494 57736 37540
rect 55927 37417 57736 37494
rect 55927 37371 55961 37417
rect 56007 37377 57736 37417
rect 56007 37371 56267 37377
rect 55927 37331 56267 37371
rect 56313 37331 57736 37377
rect 55927 37254 57736 37331
rect 55927 37208 55961 37254
rect 56007 37213 57736 37254
rect 56007 37208 56267 37213
rect 55927 37167 56267 37208
rect 56313 37167 57736 37213
rect 34717 37001 34755 37053
rect 34807 37050 34935 37053
rect 34807 37004 34916 37050
rect 34807 37001 34935 37004
rect 34987 37001 35025 37053
rect 34717 36960 35025 37001
rect 50099 37053 50408 37094
rect 50099 37001 50138 37053
rect 50190 37050 50318 37053
rect 50206 37004 50318 37050
rect 50190 37001 50318 37004
rect 50370 37001 50408 37053
rect 27387 36841 28810 36887
rect 28856 36844 29196 36887
rect 28856 36841 29116 36844
rect 27387 36798 29116 36841
rect 29162 36798 29196 36844
rect 27387 36723 29196 36798
rect 27387 36677 28810 36723
rect 28856 36681 29196 36723
rect 28856 36677 29116 36681
rect 27387 36635 29116 36677
rect 29162 36635 29196 36681
rect 27387 36560 29196 36635
rect 27387 36514 28810 36560
rect 28856 36517 29196 36560
rect 28856 36514 29116 36517
rect 27387 36471 29116 36514
rect 29162 36471 29196 36517
rect 27387 36397 29196 36471
rect 27387 36351 28810 36397
rect 28856 36354 29196 36397
rect 28856 36351 29116 36354
rect 27387 36308 29116 36351
rect 29162 36308 29196 36354
rect 27387 36234 29196 36308
rect 27387 36188 28810 36234
rect 28856 36188 29196 36234
rect 30583 36927 31040 36960
rect 34870 36953 35025 36960
rect 30583 36887 30855 36927
rect 30583 36841 30637 36887
rect 30683 36881 30855 36887
rect 30901 36881 31040 36927
rect 35294 36915 36266 36955
rect 37853 36949 38161 36957
rect 35294 36909 35332 36915
rect 35384 36909 35543 36915
rect 35595 36909 35754 36915
rect 35806 36909 35965 36915
rect 36017 36909 36176 36915
rect 36228 36909 36266 36915
rect 36438 36909 36953 36949
rect 37439 36917 38161 36949
rect 37439 36909 37891 36917
rect 37943 36909 38071 36917
rect 38123 36909 38161 36917
rect 38658 36909 39723 36969
rect 50099 36960 50408 37001
rect 52278 37053 54540 37094
rect 52278 37001 52316 37053
rect 52368 37001 52527 37053
rect 52579 37001 52738 37053
rect 52790 37001 52948 37053
rect 53000 37001 53159 37053
rect 53211 37001 53371 37053
rect 53423 37001 53582 37053
rect 53634 37001 53792 37053
rect 53844 37001 54003 37053
rect 54055 37001 54214 37053
rect 54266 37050 54540 37053
rect 54266 37004 54440 37050
rect 54486 37004 54540 37050
rect 54266 37001 54540 37004
rect 52278 36960 54540 37001
rect 54758 37053 55840 37094
rect 54758 37050 54855 37053
rect 54758 37004 54793 37050
rect 54839 37004 54855 37050
rect 54758 37001 54855 37004
rect 54907 37050 55066 37053
rect 54907 37004 54956 37050
rect 55002 37004 55066 37050
rect 54907 37001 55066 37004
rect 55118 37050 55278 37053
rect 55330 37050 55489 37053
rect 55164 37004 55278 37050
rect 55330 37004 55439 37050
rect 55485 37004 55489 37050
rect 55118 37001 55278 37004
rect 55330 37001 55489 37004
rect 55541 37050 55840 37053
rect 55541 37004 55599 37050
rect 55645 37004 55760 37050
rect 55806 37004 55840 37050
rect 55541 37001 55840 37004
rect 54758 36961 55840 37001
rect 55927 37053 57736 37167
rect 55927 37001 56015 37053
rect 56067 37001 56226 37053
rect 56278 37050 56437 37053
rect 56313 37004 56437 37050
rect 56278 37001 56437 37004
rect 56489 37001 56648 37053
rect 56700 37001 56859 37053
rect 56911 37001 57070 37053
rect 57122 37001 57281 37053
rect 57333 37001 57736 37053
rect 54817 36960 55579 36961
rect 48905 36915 49877 36955
rect 50099 36953 50255 36960
rect 48905 36909 48943 36915
rect 48995 36909 49154 36915
rect 49206 36909 49365 36915
rect 49417 36909 49576 36915
rect 49628 36909 49787 36915
rect 49839 36909 49877 36915
rect 30683 36841 31040 36881
rect 33484 36865 34643 36894
rect 30583 36764 31040 36841
rect 33019 36825 33327 36865
rect 33019 36822 33057 36825
rect 33109 36822 33237 36825
rect 33289 36822 33327 36825
rect 33484 36857 35082 36865
rect 35260 36863 35273 36909
rect 35523 36863 35543 36909
rect 35626 36863 35683 36909
rect 35729 36863 35754 36909
rect 35832 36863 35889 36909
rect 35935 36863 35965 36909
rect 36038 36863 36095 36909
rect 36141 36863 36176 36909
rect 36244 36863 36301 36909
rect 36347 36863 36360 36909
rect 36438 36863 36854 36909
rect 36900 36863 36971 36909
rect 37017 36863 37088 36909
rect 37134 36863 37206 36909
rect 37252 36863 37324 36909
rect 37370 36863 37442 36909
rect 37488 36865 37891 36909
rect 37488 36863 37909 36865
rect 37955 36863 38026 36909
rect 38123 36865 38143 36909
rect 38072 36863 38143 36865
rect 38189 36863 38261 36909
rect 38307 36863 38379 36909
rect 38425 36863 38497 36909
rect 38543 36863 38556 36909
rect 38658 36863 39021 36909
rect 39067 36863 39144 36909
rect 39190 36863 39267 36909
rect 39313 36863 39641 36909
rect 39687 36863 39730 36909
rect 31336 36776 31349 36822
rect 33323 36776 33336 36822
rect 33484 36811 33816 36857
rect 33862 36811 34002 36857
rect 34048 36811 34189 36857
rect 34235 36811 34376 36857
rect 34422 36811 34562 36857
rect 34608 36811 35082 36857
rect 35294 36823 36266 36863
rect 36438 36829 36953 36863
rect 37439 36829 38161 36863
rect 30583 36723 30855 36764
rect 30583 36677 30637 36723
rect 30683 36718 30855 36723
rect 30901 36718 31040 36764
rect 33019 36773 33057 36776
rect 33109 36773 33237 36776
rect 33289 36773 33327 36776
rect 33019 36732 33327 36773
rect 33484 36774 35082 36811
rect 30683 36677 31040 36718
rect 30583 36649 31040 36677
rect 33484 36692 33552 36774
rect 30583 36601 31493 36649
rect 30583 36560 30855 36601
rect 30583 36514 30637 36560
rect 30683 36555 30855 36560
rect 30901 36598 31493 36601
rect 30901 36555 31349 36598
rect 30683 36552 31349 36555
rect 33323 36552 33336 36598
rect 30683 36530 31493 36552
rect 30683 36514 31040 36530
rect 30583 36438 31040 36514
rect 30583 36397 30855 36438
rect 30583 36351 30637 36397
rect 30683 36392 30855 36397
rect 30901 36392 31040 36438
rect 30683 36351 31040 36392
rect 33019 36377 33327 36417
rect 33019 36374 33057 36377
rect 33109 36374 33237 36377
rect 33289 36374 33327 36377
rect 30583 36274 31040 36351
rect 31336 36328 31349 36374
rect 33323 36328 33336 36374
rect 33019 36325 33057 36328
rect 33109 36325 33237 36328
rect 33289 36325 33327 36328
rect 33019 36284 33327 36325
rect 30583 36234 30855 36274
rect 27387 35985 29196 36188
rect 29283 36153 30365 36194
rect 29283 36150 29582 36153
rect 29283 36104 29317 36150
rect 29363 36104 29478 36150
rect 29524 36104 29582 36150
rect 29283 36101 29582 36104
rect 29634 36150 29793 36153
rect 29845 36150 30005 36153
rect 29634 36104 29638 36150
rect 29684 36104 29793 36150
rect 29845 36104 29959 36150
rect 29634 36101 29793 36104
rect 29845 36101 30005 36104
rect 30057 36150 30216 36153
rect 30057 36104 30121 36150
rect 30167 36104 30216 36150
rect 30057 36101 30216 36104
rect 30268 36150 30365 36153
rect 30268 36104 30284 36150
rect 30330 36104 30365 36150
rect 30268 36101 30365 36104
rect 29283 36061 30365 36101
rect 30583 36188 30637 36234
rect 30683 36228 30855 36234
rect 30901 36228 31040 36274
rect 33484 36270 33495 36692
rect 33541 36270 33552 36692
rect 34964 36717 35082 36774
rect 36438 36729 36554 36829
rect 37853 36824 38161 36829
rect 38658 36849 39723 36863
rect 34964 36685 36360 36717
rect 34228 36615 34718 36656
rect 34228 36598 34267 36615
rect 34319 36598 34447 36615
rect 34499 36598 34627 36615
rect 33671 36552 33684 36598
rect 33730 36552 33787 36598
rect 33833 36552 33890 36598
rect 33936 36552 33993 36598
rect 34039 36552 34096 36598
rect 34142 36552 34199 36598
rect 34245 36563 34267 36598
rect 34245 36552 34302 36563
rect 34348 36552 34405 36598
rect 34499 36563 34508 36598
rect 34451 36552 34508 36563
rect 34554 36552 34612 36598
rect 34679 36563 34718 36615
rect 34964 36639 35273 36685
rect 35523 36639 35580 36685
rect 35626 36639 35683 36685
rect 35729 36639 35786 36685
rect 35832 36639 35889 36685
rect 35935 36639 35992 36685
rect 36038 36639 36095 36685
rect 36141 36639 36198 36685
rect 36244 36639 36301 36685
rect 36347 36639 36360 36685
rect 34964 36595 36360 36639
rect 34658 36552 34718 36563
rect 34228 36523 34718 36552
rect 36438 36589 36475 36729
rect 36521 36589 36554 36729
rect 35294 36461 36266 36495
rect 36438 36486 36554 36589
rect 36640 36729 36773 36749
rect 36640 36690 36697 36729
rect 36640 36638 36678 36690
rect 36640 36589 36697 36638
rect 36743 36589 36773 36729
rect 38658 36727 38726 36849
rect 39809 36843 44918 36881
rect 48765 36863 48778 36909
rect 48824 36863 48881 36909
rect 48927 36863 48943 36909
rect 49030 36863 49087 36909
rect 49133 36863 49154 36909
rect 49236 36863 49293 36909
rect 49339 36863 49365 36909
rect 49442 36863 49499 36909
rect 49545 36863 49576 36909
rect 49852 36863 49877 36909
rect 54085 36927 54540 36960
rect 50481 36867 51657 36894
rect 39809 36797 43739 36843
rect 43785 36797 43906 36843
rect 43952 36797 44071 36843
rect 44117 36797 44236 36843
rect 44282 36822 44918 36843
rect 48905 36823 49877 36863
rect 50044 36857 51657 36867
rect 44282 36797 44812 36822
rect 39809 36794 44812 36797
rect 39809 36748 39844 36794
rect 39890 36792 44812 36794
rect 39890 36748 39994 36792
rect 39809 36740 39994 36748
rect 40046 36776 44812 36792
rect 44858 36776 44925 36822
rect 44971 36776 45038 36822
rect 45084 36776 45151 36822
rect 45197 36776 45264 36822
rect 45310 36776 45323 36822
rect 48557 36777 48687 36817
rect 40046 36761 44918 36776
rect 40046 36740 40085 36761
rect 39809 36737 40085 36740
rect 36924 36717 37685 36724
rect 36923 36685 37931 36717
rect 36841 36639 36854 36685
rect 36900 36683 36971 36685
rect 36900 36639 36961 36683
rect 37017 36639 37088 36685
rect 37134 36683 37206 36685
rect 37134 36639 37172 36683
rect 37252 36639 37324 36685
rect 37370 36683 37442 36685
rect 37370 36639 37384 36683
rect 36923 36631 36961 36639
rect 37013 36631 37172 36639
rect 37224 36631 37384 36639
rect 37436 36639 37442 36683
rect 37488 36683 37909 36685
rect 37488 36639 37595 36683
rect 37436 36631 37595 36639
rect 37647 36639 37909 36683
rect 37955 36639 38026 36685
rect 38072 36639 38143 36685
rect 38189 36639 38261 36685
rect 38307 36639 38379 36685
rect 38425 36639 38497 36685
rect 38543 36639 38556 36685
rect 37647 36631 37931 36639
rect 36923 36598 37931 36631
rect 36923 36597 37685 36598
rect 36924 36591 37685 36597
rect 36640 36566 36773 36589
rect 38658 36587 38669 36727
rect 38715 36587 38726 36727
rect 39014 36685 39323 36717
rect 39492 36685 39608 36717
rect 39008 36639 39021 36685
rect 39067 36639 39144 36685
rect 39190 36639 39267 36685
rect 39313 36639 39326 36685
rect 39492 36639 39641 36685
rect 39687 36639 39730 36685
rect 38658 36576 38726 36587
rect 36438 36461 36953 36486
rect 37439 36483 37931 36486
rect 37439 36461 38161 36483
rect 35260 36415 35273 36461
rect 35523 36455 35580 36461
rect 35523 36415 35543 36455
rect 35626 36415 35683 36461
rect 35729 36455 35786 36461
rect 35729 36415 35754 36455
rect 35832 36415 35889 36461
rect 35935 36455 35992 36461
rect 35935 36415 35965 36455
rect 36038 36415 36095 36461
rect 36141 36455 36198 36461
rect 36141 36415 36176 36455
rect 36244 36415 36301 36461
rect 36347 36415 36360 36461
rect 36438 36415 36854 36461
rect 36900 36415 36971 36461
rect 37017 36415 37088 36461
rect 37134 36415 37206 36461
rect 37252 36415 37324 36461
rect 37370 36415 37442 36461
rect 37488 36443 37909 36461
rect 37488 36415 37891 36443
rect 37955 36415 38026 36461
rect 38072 36443 38143 36461
rect 38123 36415 38143 36443
rect 38189 36415 38261 36461
rect 38307 36415 38379 36461
rect 38425 36415 38497 36461
rect 38543 36415 38556 36461
rect 33781 36374 34089 36409
rect 35294 36403 35332 36415
rect 35384 36403 35543 36415
rect 35595 36403 35754 36415
rect 35806 36403 35965 36415
rect 36017 36403 36176 36415
rect 36228 36403 36266 36415
rect 33671 36328 33684 36374
rect 33730 36328 33787 36374
rect 33833 36369 33890 36374
rect 33871 36328 33890 36369
rect 33936 36328 33993 36374
rect 34039 36369 34096 36374
rect 34051 36328 34096 36369
rect 34142 36328 34199 36374
rect 34245 36328 34302 36374
rect 34348 36328 34405 36374
rect 34451 36328 34508 36374
rect 34554 36328 34612 36374
rect 34658 36328 34671 36374
rect 35294 36363 36266 36403
rect 36438 36366 36953 36415
rect 37439 36391 37891 36415
rect 37943 36391 38071 36415
rect 38123 36391 38161 36415
rect 37439 36366 38161 36391
rect 37853 36350 38161 36366
rect 33781 36317 33819 36328
rect 33871 36317 33999 36328
rect 34051 36317 34089 36328
rect 33781 36276 34089 36317
rect 33484 36259 33552 36270
rect 30683 36194 31040 36228
rect 30683 36188 32842 36194
rect 30583 36153 32842 36188
rect 34247 36187 35008 36194
rect 30583 36101 30854 36153
rect 30906 36101 31065 36153
rect 31117 36101 31276 36153
rect 31328 36150 31486 36153
rect 31538 36150 31697 36153
rect 31749 36150 31909 36153
rect 31961 36150 32120 36153
rect 32172 36150 32330 36153
rect 32382 36150 32541 36153
rect 32593 36150 32752 36153
rect 32804 36150 32842 36153
rect 34246 36153 35008 36187
rect 34246 36150 34284 36153
rect 34336 36150 34495 36153
rect 34547 36150 34707 36153
rect 31328 36104 31349 36150
rect 33323 36104 33336 36150
rect 33671 36104 33684 36150
rect 33730 36104 33787 36150
rect 33833 36104 33890 36150
rect 33936 36104 33993 36150
rect 34039 36104 34096 36150
rect 34142 36104 34199 36150
rect 34245 36104 34284 36150
rect 34348 36104 34405 36150
rect 34451 36104 34495 36150
rect 34554 36104 34612 36150
rect 34658 36104 34707 36150
rect 31328 36101 31486 36104
rect 31538 36101 31697 36104
rect 31749 36101 31909 36104
rect 31961 36101 32120 36104
rect 32172 36101 32330 36104
rect 32382 36101 32541 36104
rect 32593 36101 32752 36104
rect 32804 36101 32842 36104
rect 30583 36061 32842 36101
rect 34246 36101 34284 36104
rect 34336 36101 34495 36104
rect 34547 36101 34707 36104
rect 34759 36101 34918 36153
rect 34970 36101 35008 36153
rect 34246 36067 35008 36101
rect 34247 36061 35008 36067
rect 35182 36187 36364 36194
rect 35182 36153 36958 36187
rect 35182 36101 35220 36153
rect 35272 36101 35430 36153
rect 35482 36101 35641 36153
rect 35693 36101 35853 36153
rect 35905 36101 36064 36153
rect 36116 36101 36274 36153
rect 36326 36150 36958 36153
rect 36326 36104 36489 36150
rect 36723 36104 36958 36150
rect 36326 36101 36958 36104
rect 35182 36067 36958 36101
rect 37946 36153 38842 36194
rect 37946 36150 38330 36153
rect 38382 36150 38541 36153
rect 37946 36104 37957 36150
rect 38473 36104 38541 36150
rect 37946 36101 38330 36104
rect 38382 36101 38541 36104
rect 38593 36101 38752 36153
rect 38804 36101 38842 36153
rect 29544 36060 30306 36061
rect 30748 36060 32842 36061
rect 35182 36060 36364 36067
rect 37946 36061 38842 36101
rect 39014 36153 39323 36639
rect 39014 36101 39052 36153
rect 39104 36150 39232 36153
rect 39108 36104 39220 36150
rect 39104 36101 39232 36104
rect 39284 36101 39323 36153
rect 39014 36067 39323 36101
rect 39492 36187 39608 36639
rect 39923 36606 40085 36737
rect 39923 36554 39994 36606
rect 40046 36554 40085 36606
rect 39923 36514 40085 36554
rect 39737 36418 39865 36431
rect 39737 36391 39866 36418
rect 39737 36374 39775 36391
rect 39827 36374 39866 36391
rect 39727 36328 39740 36374
rect 39827 36339 39862 36374
rect 39786 36328 39862 36339
rect 39908 36328 39985 36374
rect 40031 36328 40108 36374
rect 40154 36328 40167 36374
rect 40246 36363 40362 36761
rect 42229 36622 44509 36663
rect 42229 36570 43445 36622
rect 43497 36570 44509 36622
rect 42229 36530 44509 36570
rect 44341 36486 44509 36530
rect 44341 36440 44358 36486
rect 44498 36440 44509 36486
rect 39737 36299 39866 36328
rect 40246 36317 40281 36363
rect 40327 36317 40362 36363
rect 40246 36280 40362 36317
rect 40718 36391 43524 36432
rect 44341 36429 44509 36440
rect 40718 36339 41935 36391
rect 41987 36339 43524 36391
rect 40718 36298 43524 36339
rect 44605 36374 44721 36761
rect 45400 36731 48379 36772
rect 45400 36717 48241 36731
rect 45400 36671 45464 36717
rect 45604 36679 48241 36717
rect 48293 36679 48379 36731
rect 45604 36671 48379 36679
rect 44901 36615 45241 36656
rect 45400 36638 48379 36671
rect 48557 36725 48596 36777
rect 48648 36725 48687 36777
rect 48557 36702 48687 36725
rect 50044 36811 50516 36857
rect 50562 36811 50703 36857
rect 50749 36811 50890 36857
rect 50936 36811 51076 36857
rect 51122 36811 51263 36857
rect 51309 36811 51657 36857
rect 51797 36847 52105 36887
rect 51797 36822 51835 36847
rect 51887 36822 52015 36847
rect 52067 36822 52105 36847
rect 54085 36881 54223 36927
rect 54269 36887 54540 36927
rect 54269 36881 54440 36887
rect 54085 36841 54440 36881
rect 54486 36841 54540 36887
rect 50044 36774 51657 36811
rect 51789 36776 51802 36822
rect 53776 36776 53789 36822
rect 50044 36717 50160 36774
rect 44901 36598 44939 36615
rect 44991 36598 45151 36615
rect 45203 36598 45241 36615
rect 44799 36552 44812 36598
rect 44858 36552 44925 36598
rect 44991 36563 45038 36598
rect 44971 36552 45038 36563
rect 45084 36552 45151 36598
rect 45203 36563 45264 36598
rect 45197 36552 45264 36563
rect 45310 36552 45323 36598
rect 48557 36562 48622 36702
rect 48668 36562 48687 36702
rect 49820 36685 50160 36717
rect 48765 36639 48778 36685
rect 48824 36639 48881 36685
rect 48927 36639 48984 36685
rect 49030 36639 49087 36685
rect 49133 36639 49190 36685
rect 49236 36639 49293 36685
rect 49339 36639 49396 36685
rect 49442 36639 49499 36685
rect 49545 36639 49602 36685
rect 49852 36639 50160 36685
rect 51589 36722 51657 36774
rect 51797 36754 52105 36776
rect 49820 36598 50160 36639
rect 50262 36615 50812 36656
rect 48557 36559 48687 36562
rect 44901 36523 45241 36552
rect 48557 36507 48596 36559
rect 48648 36507 48687 36559
rect 50262 36563 50300 36615
rect 50352 36598 50511 36615
rect 50563 36598 50722 36615
rect 50352 36563 50467 36598
rect 50563 36563 50571 36598
rect 50262 36552 50467 36563
rect 50513 36552 50571 36563
rect 50617 36552 50674 36598
rect 50720 36563 50722 36598
rect 50774 36598 50812 36615
rect 50774 36563 50777 36598
rect 50720 36552 50777 36563
rect 50823 36552 50880 36598
rect 50926 36552 50983 36598
rect 51029 36552 51086 36598
rect 51132 36552 51189 36598
rect 51235 36552 51292 36598
rect 51338 36552 51395 36598
rect 51441 36552 51454 36598
rect 50262 36523 50812 36552
rect 48557 36466 48687 36507
rect 48905 36461 49877 36492
rect 48765 36415 48778 36461
rect 48824 36415 48881 36461
rect 48927 36452 48984 36461
rect 48927 36415 48943 36452
rect 49030 36415 49087 36461
rect 49133 36452 49190 36461
rect 49133 36415 49154 36452
rect 49236 36415 49293 36461
rect 49339 36452 49396 36461
rect 49339 36415 49365 36452
rect 49442 36415 49499 36461
rect 49545 36452 49602 36461
rect 49545 36415 49576 36452
rect 49852 36415 49877 36461
rect 48905 36400 48943 36415
rect 48995 36400 49154 36415
rect 49206 36400 49365 36415
rect 49417 36400 49576 36415
rect 49628 36400 49787 36415
rect 49839 36400 49877 36415
rect 44605 36328 44812 36374
rect 44858 36328 44925 36374
rect 44971 36328 45038 36374
rect 45084 36328 45151 36374
rect 45197 36328 45264 36374
rect 45310 36328 45323 36374
rect 48905 36360 49877 36400
rect 51035 36377 51343 36417
rect 51035 36374 51073 36377
rect 51125 36374 51253 36377
rect 51305 36374 51343 36377
rect 43362 36291 43524 36298
rect 43362 36245 43373 36291
rect 43513 36245 43524 36291
rect 43362 36234 43524 36245
rect 45584 36314 48546 36350
rect 50454 36328 50467 36374
rect 50513 36328 50571 36374
rect 50617 36328 50674 36374
rect 50720 36328 50777 36374
rect 50823 36328 50880 36374
rect 50926 36328 50983 36374
rect 51029 36328 51073 36374
rect 51132 36328 51189 36374
rect 51235 36328 51253 36374
rect 51338 36328 51395 36374
rect 51441 36328 51454 36374
rect 45584 36268 45619 36314
rect 45665 36268 45777 36314
rect 45823 36268 45935 36314
rect 45981 36268 46093 36314
rect 46139 36268 46251 36314
rect 46297 36268 46409 36314
rect 46455 36268 46568 36314
rect 46614 36268 46726 36314
rect 46772 36268 46884 36314
rect 46930 36268 47042 36314
rect 47088 36268 47200 36314
rect 47246 36268 47358 36314
rect 47404 36268 47516 36314
rect 47562 36268 47675 36314
rect 47721 36268 47833 36314
rect 47879 36268 47991 36314
rect 48037 36268 48149 36314
rect 48195 36268 48307 36314
rect 48353 36268 48465 36314
rect 48511 36268 48546 36314
rect 51035 36325 51073 36328
rect 51125 36325 51253 36328
rect 51305 36325 51343 36328
rect 51035 36284 51343 36325
rect 51589 36300 51600 36722
rect 51646 36300 51657 36722
rect 54085 36723 54540 36841
rect 54085 36677 54440 36723
rect 54486 36677 54540 36723
rect 54085 36649 54540 36677
rect 53585 36598 54540 36649
rect 51789 36552 51802 36598
rect 53776 36560 54540 36598
rect 53776 36552 54440 36560
rect 53585 36530 54440 36552
rect 54085 36514 54440 36530
rect 54486 36514 54540 36560
rect 54085 36438 54540 36514
rect 51797 36384 52105 36424
rect 51797 36374 51835 36384
rect 51887 36374 52015 36384
rect 52067 36374 52105 36384
rect 54085 36392 54223 36438
rect 54269 36397 54540 36438
rect 54269 36392 54440 36397
rect 51789 36328 51802 36374
rect 53776 36328 53789 36374
rect 54085 36351 54440 36392
rect 54486 36351 54540 36397
rect 51589 36289 51657 36300
rect 51797 36291 52105 36328
rect 40215 36187 40523 36193
rect 40788 36187 42986 36201
rect 43753 36187 44514 36194
rect 39492 36164 42986 36187
rect 43704 36164 44514 36187
rect 39492 36153 44514 36164
rect 39492 36150 40253 36153
rect 39492 36104 39740 36150
rect 39786 36104 39862 36150
rect 39908 36104 39985 36150
rect 40031 36104 40108 36150
rect 40154 36104 40253 36150
rect 39492 36101 40253 36104
rect 40305 36101 40433 36153
rect 40485 36150 43790 36153
rect 40485 36104 40836 36150
rect 40882 36104 40994 36150
rect 41040 36104 41152 36150
rect 41198 36104 41310 36150
rect 41356 36104 41469 36150
rect 41515 36104 41627 36150
rect 41673 36104 41785 36150
rect 41831 36104 41943 36150
rect 41989 36104 42101 36150
rect 42147 36104 42259 36150
rect 42305 36104 42418 36150
rect 42464 36104 42576 36150
rect 42622 36104 42734 36150
rect 42780 36104 42892 36150
rect 42938 36104 43739 36150
rect 43785 36104 43790 36150
rect 40485 36101 43790 36104
rect 43842 36150 44001 36153
rect 43842 36104 43906 36150
rect 43952 36104 44001 36150
rect 43842 36101 44001 36104
rect 44053 36150 44213 36153
rect 44265 36150 44424 36153
rect 44053 36104 44071 36150
rect 44117 36104 44213 36150
rect 44282 36104 44424 36150
rect 44053 36101 44213 36104
rect 44265 36101 44424 36104
rect 44476 36101 44514 36153
rect 39492 36090 44514 36101
rect 39492 36067 42986 36090
rect 43704 36067 44514 36090
rect 37946 36060 38324 36061
rect 39014 36060 39322 36067
rect 40215 36060 40523 36067
rect 40788 36053 42986 36067
rect 43753 36061 44514 36067
rect 44796 36187 45346 36194
rect 45584 36187 48546 36268
rect 54085 36274 54540 36351
rect 54085 36228 54223 36274
rect 54269 36234 54540 36274
rect 54269 36228 54440 36234
rect 54085 36194 54440 36228
rect 48800 36187 49982 36194
rect 50308 36187 50859 36194
rect 44796 36153 49982 36187
rect 44796 36150 44834 36153
rect 44886 36150 45045 36153
rect 45097 36150 45256 36153
rect 45308 36150 48838 36153
rect 44796 36104 44812 36150
rect 44886 36104 44925 36150
rect 44971 36104 45038 36150
rect 45097 36104 45151 36150
rect 45197 36104 45256 36150
rect 45310 36104 45619 36150
rect 45665 36104 45777 36150
rect 45823 36104 45935 36150
rect 45981 36104 46093 36150
rect 46139 36104 46251 36150
rect 46297 36104 46409 36150
rect 46455 36104 46568 36150
rect 46614 36104 46726 36150
rect 46772 36104 46884 36150
rect 46930 36104 47042 36150
rect 47088 36104 47200 36150
rect 47246 36104 47358 36150
rect 47404 36104 47516 36150
rect 47562 36104 47675 36150
rect 47721 36104 47833 36150
rect 47879 36104 47991 36150
rect 48037 36104 48149 36150
rect 48195 36104 48307 36150
rect 48353 36104 48465 36150
rect 48511 36104 48838 36150
rect 44796 36101 44834 36104
rect 44886 36101 45045 36104
rect 45097 36101 45256 36104
rect 45308 36101 48838 36104
rect 48890 36101 49048 36153
rect 49100 36101 49259 36153
rect 49311 36101 49471 36153
rect 49523 36101 49682 36153
rect 49734 36101 49892 36153
rect 49944 36101 49982 36153
rect 44796 36067 49982 36101
rect 50307 36153 50859 36187
rect 50307 36101 50346 36153
rect 50398 36150 50557 36153
rect 50609 36150 50768 36153
rect 50820 36150 50859 36153
rect 52278 36188 54440 36194
rect 54486 36188 54540 36234
rect 55927 36887 57736 37001
rect 55927 36844 56267 36887
rect 55927 36798 55961 36844
rect 56007 36841 56267 36844
rect 56313 36841 57736 36887
rect 56007 36798 57736 36841
rect 55927 36723 57736 36798
rect 55927 36681 56267 36723
rect 55927 36635 55961 36681
rect 56007 36677 56267 36681
rect 56313 36677 57736 36723
rect 56007 36635 57736 36677
rect 55927 36560 57736 36635
rect 55927 36517 56267 36560
rect 55927 36471 55961 36517
rect 56007 36514 56267 36517
rect 56313 36514 57736 36560
rect 56007 36471 57736 36514
rect 55927 36397 57736 36471
rect 55927 36354 56267 36397
rect 55927 36308 55961 36354
rect 56007 36351 56267 36354
rect 56313 36351 57736 36397
rect 56007 36308 57736 36351
rect 55927 36234 57736 36308
rect 52278 36153 54540 36188
rect 52278 36150 52316 36153
rect 52368 36150 52527 36153
rect 52579 36150 52738 36153
rect 52790 36150 52948 36153
rect 53000 36150 53159 36153
rect 53211 36150 53371 36153
rect 53423 36150 53582 36153
rect 53634 36150 53792 36153
rect 50398 36104 50467 36150
rect 50513 36104 50557 36150
rect 50617 36104 50674 36150
rect 50720 36104 50768 36150
rect 50823 36104 50880 36150
rect 50926 36104 50983 36150
rect 51029 36104 51086 36150
rect 51132 36104 51189 36150
rect 51235 36104 51292 36150
rect 51338 36104 51395 36150
rect 51441 36104 51454 36150
rect 51789 36104 51802 36150
rect 53776 36104 53792 36150
rect 50398 36101 50557 36104
rect 50609 36101 50768 36104
rect 50820 36101 50859 36104
rect 50307 36067 50859 36101
rect 44796 36061 45346 36067
rect 48800 36060 49982 36067
rect 50308 36060 50859 36067
rect 52278 36101 52316 36104
rect 52368 36101 52527 36104
rect 52579 36101 52738 36104
rect 52790 36101 52948 36104
rect 53000 36101 53159 36104
rect 53211 36101 53371 36104
rect 53423 36101 53582 36104
rect 53634 36101 53792 36104
rect 53844 36101 54003 36153
rect 54055 36101 54214 36153
rect 54266 36101 54540 36153
rect 52278 36061 54540 36101
rect 54758 36153 55840 36194
rect 54758 36150 54855 36153
rect 54758 36104 54793 36150
rect 54839 36104 54855 36150
rect 54758 36101 54855 36104
rect 54907 36150 55066 36153
rect 54907 36104 54956 36150
rect 55002 36104 55066 36150
rect 54907 36101 55066 36104
rect 55118 36150 55278 36153
rect 55330 36150 55489 36153
rect 55164 36104 55278 36150
rect 55330 36104 55439 36150
rect 55485 36104 55489 36150
rect 55118 36101 55278 36104
rect 55330 36101 55489 36104
rect 55541 36150 55840 36153
rect 55541 36104 55599 36150
rect 55645 36104 55760 36150
rect 55806 36104 55840 36150
rect 55541 36101 55840 36104
rect 54758 36061 55840 36101
rect 55927 36188 56267 36234
rect 56313 36188 57736 36234
rect 52278 36060 54377 36061
rect 54817 36060 55579 36061
rect 55927 35985 57736 36188
rect 25334 34959 26030 34971
rect 25334 34909 25346 34959
rect 24362 34907 25346 34909
rect 25398 34907 25470 34959
rect 25522 34907 25594 34959
rect 25646 34907 25718 34959
rect 25770 34907 25842 34959
rect 25894 34907 25966 34959
rect 26018 34909 26030 34959
rect 27387 34960 27828 35985
rect 27387 34909 27469 34960
rect 26018 34907 27469 34909
rect 24362 34835 27469 34907
rect 24362 34783 25346 34835
rect 25398 34783 25470 34835
rect 25522 34783 25594 34835
rect 25646 34783 25718 34835
rect 25770 34783 25842 34835
rect 25894 34783 25966 34835
rect 26018 34783 27469 34835
rect 24362 34739 27469 34783
rect 25334 34711 26030 34739
rect 25334 34659 25346 34711
rect 25398 34659 25470 34711
rect 25522 34659 25594 34711
rect 25646 34659 25718 34711
rect 25770 34659 25842 34711
rect 25894 34659 25966 34711
rect 26018 34659 26030 34711
rect 25334 34647 26030 34659
rect 27387 34596 27469 34739
rect 27729 34655 27828 34960
rect 57295 34909 57736 35985
rect 58812 34979 59508 34991
rect 58812 34927 58824 34979
rect 58876 34927 58948 34979
rect 59000 34927 59072 34979
rect 59124 34927 59196 34979
rect 59248 34927 59320 34979
rect 59372 34927 59444 34979
rect 59496 34927 59508 34979
rect 58812 34909 59508 34927
rect 57295 34855 61058 34909
rect 57295 34803 58824 34855
rect 58876 34803 58948 34855
rect 59000 34803 59072 34855
rect 59124 34803 59196 34855
rect 59248 34803 59320 34855
rect 59372 34803 59444 34855
rect 59496 34803 61058 34855
rect 57295 34739 61058 34803
rect 57295 34655 57736 34739
rect 58812 34731 59508 34739
rect 58812 34679 58824 34731
rect 58876 34679 58948 34731
rect 59000 34679 59072 34731
rect 59124 34679 59196 34731
rect 59248 34679 59320 34731
rect 59372 34679 59444 34731
rect 59496 34679 59508 34731
rect 58812 34667 59508 34679
rect 27729 34596 57736 34655
rect 27387 34199 57736 34596
rect 26772 33432 27214 33519
rect 26772 33380 26861 33432
rect 26913 33380 27073 33432
rect 27125 33380 27214 33432
rect 26772 33215 27214 33380
rect 26772 33163 26861 33215
rect 26913 33163 27073 33215
rect 27125 33163 27214 33215
rect 26772 32997 27214 33163
rect 26772 32945 26861 32997
rect 26913 32945 27073 32997
rect 27125 32945 27214 32997
rect 26772 32779 27214 32945
rect 26772 32727 26861 32779
rect 26913 32727 27073 32779
rect 27125 32727 27214 32779
rect 26772 32562 27214 32727
rect 26772 32510 26861 32562
rect 26913 32510 27073 32562
rect 27125 32510 27214 32562
rect 26772 32344 27214 32510
rect 26772 32292 26861 32344
rect 26913 32292 27073 32344
rect 27125 32292 27214 32344
rect 26772 32127 27214 32292
rect 26772 32075 26861 32127
rect 26913 32075 27073 32127
rect 27125 32075 27214 32127
rect 26772 31909 27214 32075
rect 26772 31857 26861 31909
rect 26913 31857 27073 31909
rect 27125 31857 27214 31909
rect 26772 31691 27214 31857
rect 26772 31639 26861 31691
rect 26913 31639 27073 31691
rect 27125 31639 27214 31691
rect 26772 31474 27214 31639
rect 26772 31422 26861 31474
rect 26913 31422 27073 31474
rect 27125 31422 27214 31474
rect 26772 31256 27214 31422
rect 26772 31204 26861 31256
rect 26913 31204 27073 31256
rect 27125 31204 27214 31256
rect 26772 31038 27214 31204
rect 26772 30986 26861 31038
rect 26913 30986 27073 31038
rect 27125 30986 27214 31038
rect 26772 30821 27214 30986
rect 26772 30769 26861 30821
rect 26913 30769 27073 30821
rect 27125 30769 27214 30821
rect 26772 30603 27214 30769
rect 26772 30551 26861 30603
rect 26913 30551 27073 30603
rect 27125 30551 27214 30603
rect 26772 30386 27214 30551
rect 26772 30334 26861 30386
rect 26913 30334 27073 30386
rect 27125 30334 27214 30386
rect 26772 30168 27214 30334
rect 26772 30116 26861 30168
rect 26913 30116 27073 30168
rect 27125 30116 27214 30168
rect 26772 29950 27214 30116
rect 26772 29898 26861 29950
rect 26913 29898 27073 29950
rect 27125 29898 27214 29950
rect 26772 29733 27214 29898
rect 26772 29681 26861 29733
rect 26913 29681 27073 29733
rect 27125 29681 27214 29733
rect 26772 29515 27214 29681
rect 26772 29463 26861 29515
rect 26913 29463 27073 29515
rect 27125 29463 27214 29515
rect 26772 29297 27214 29463
rect 26772 29245 26861 29297
rect 26913 29245 27073 29297
rect 27125 29245 27214 29297
rect 26772 29080 27214 29245
rect 26772 29028 26861 29080
rect 26913 29028 27073 29080
rect 27125 29028 27214 29080
rect 26772 28862 27214 29028
rect 26772 28810 26861 28862
rect 26913 28810 27073 28862
rect 27125 28810 27214 28862
rect 26772 28644 27214 28810
rect 26772 28592 26861 28644
rect 26913 28592 27073 28644
rect 27125 28592 27214 28644
rect 26772 28427 27214 28592
rect 26772 28375 26861 28427
rect 26913 28375 27073 28427
rect 27125 28375 27214 28427
rect 26772 28209 27214 28375
rect 26772 28157 26861 28209
rect 26913 28157 27073 28209
rect 27125 28157 27214 28209
rect 26772 27992 27214 28157
rect 26772 27940 26861 27992
rect 26913 27940 27073 27992
rect 27125 27940 27214 27992
rect 26772 27774 27214 27940
rect 26772 27722 26861 27774
rect 26913 27722 27073 27774
rect 27125 27722 27214 27774
rect 26772 27556 27214 27722
rect 26772 27504 26861 27556
rect 26913 27504 27073 27556
rect 27125 27504 27214 27556
rect 26772 27339 27214 27504
rect 26772 27287 26861 27339
rect 26913 27287 27073 27339
rect 27125 27287 27214 27339
rect 26772 27121 27214 27287
rect 26772 27069 26861 27121
rect 26913 27069 27073 27121
rect 27125 27069 27214 27121
rect 26772 26903 27214 27069
rect 26772 26851 26861 26903
rect 26913 26851 27073 26903
rect 27125 26851 27214 26903
rect 26772 26686 27214 26851
rect 26772 26634 26861 26686
rect 26913 26634 27073 26686
rect 27125 26634 27214 26686
rect 26772 26468 27214 26634
rect 26772 26416 26861 26468
rect 26913 26416 27073 26468
rect 27125 26416 27214 26468
rect 26772 26250 27214 26416
rect 26772 26198 26861 26250
rect 26913 26198 27073 26250
rect 27125 26198 27214 26250
rect 26772 26033 27214 26198
rect 26772 25981 26861 26033
rect 26913 25981 27073 26033
rect 27125 25981 27214 26033
rect 26772 25815 27214 25981
rect 26772 25763 26861 25815
rect 26913 25763 27073 25815
rect 27125 25763 27214 25815
rect 26772 25598 27214 25763
rect 26772 25546 26861 25598
rect 26913 25546 27073 25598
rect 27125 25546 27214 25598
rect 26772 25380 27214 25546
rect 26772 25328 26861 25380
rect 26913 25328 27073 25380
rect 27125 25328 27214 25380
rect 26772 25162 27214 25328
rect 26772 25110 26861 25162
rect 26913 25110 27073 25162
rect 27125 25110 27214 25162
rect 26772 24945 27214 25110
rect 26772 24893 26861 24945
rect 26913 24893 27073 24945
rect 27125 24893 27214 24945
rect 26772 24727 27214 24893
rect 26772 24675 26861 24727
rect 26913 24675 27073 24727
rect 27125 24675 27214 24727
rect 26772 24509 27214 24675
rect 26772 24457 26861 24509
rect 26913 24457 27073 24509
rect 27125 24457 27214 24509
rect 26772 24292 27214 24457
rect 26772 24240 26861 24292
rect 26913 24240 27073 24292
rect 27125 24240 27214 24292
rect 26772 24074 27214 24240
rect 26772 24022 26861 24074
rect 26913 24022 27073 24074
rect 27125 24022 27214 24074
rect 26772 23857 27214 24022
rect 26772 23805 26861 23857
rect 26913 23805 27073 23857
rect 27125 23805 27214 23857
rect 26772 23639 27214 23805
rect 26772 23587 26861 23639
rect 26913 23587 27073 23639
rect 27125 23587 27214 23639
rect 26772 23421 27214 23587
rect 26772 23369 26861 23421
rect 26913 23369 27073 23421
rect 27125 23369 27214 23421
rect 26772 23204 27214 23369
rect 26772 23152 26861 23204
rect 26913 23152 27073 23204
rect 27125 23152 27214 23204
rect 26772 22986 27214 23152
rect 26772 22934 26861 22986
rect 26913 22934 27073 22986
rect 27125 22934 27214 22986
rect 26772 22768 27214 22934
rect 26772 22716 26861 22768
rect 26913 22716 27073 22768
rect 27125 22716 27214 22768
rect 26772 22551 27214 22716
rect 26772 22499 26861 22551
rect 26913 22499 27073 22551
rect 27125 22499 27214 22551
rect 26772 22333 27214 22499
rect 26772 22281 26861 22333
rect 26913 22281 27073 22333
rect 27125 22281 27214 22333
rect 26772 22115 27214 22281
rect 26772 22063 26861 22115
rect 26913 22063 27073 22115
rect 27125 22063 27214 22115
rect 26772 21898 27214 22063
rect 26772 21846 26861 21898
rect 26913 21846 27073 21898
rect 27125 21846 27214 21898
rect 26772 21680 27214 21846
rect 26772 21628 26861 21680
rect 26913 21628 27073 21680
rect 27125 21628 27214 21680
rect 26772 21463 27214 21628
rect 26772 21411 26861 21463
rect 26913 21411 27073 21463
rect 27125 21411 27214 21463
rect 26772 21245 27214 21411
rect 26772 21193 26861 21245
rect 26913 21193 27073 21245
rect 27125 21193 27214 21245
rect 26772 21027 27214 21193
rect 26772 20975 26861 21027
rect 26913 20975 27073 21027
rect 27125 20975 27214 21027
rect 26772 20810 27214 20975
rect 26772 20758 26861 20810
rect 26913 20758 27073 20810
rect 27125 20758 27214 20810
rect 26772 20592 27214 20758
rect 26772 20540 26861 20592
rect 26913 20540 27073 20592
rect 27125 20540 27214 20592
rect 26772 20374 27214 20540
rect 26772 20322 26861 20374
rect 26913 20322 27073 20374
rect 27125 20322 27214 20374
rect 26772 20157 27214 20322
rect 26772 20105 26861 20157
rect 26913 20105 27073 20157
rect 27125 20105 27214 20157
rect 26772 19939 27214 20105
rect 26772 19887 26861 19939
rect 26913 19887 27073 19939
rect 27125 19887 27214 19939
rect 26772 19722 27214 19887
rect 26772 19670 26861 19722
rect 26913 19670 27073 19722
rect 27125 19670 27214 19722
rect 26772 19504 27214 19670
rect 26772 19452 26861 19504
rect 26913 19452 27073 19504
rect 27125 19452 27214 19504
rect 26772 19286 27214 19452
rect 26772 19234 26861 19286
rect 26913 19234 27073 19286
rect 27125 19234 27214 19286
rect 26772 19068 27214 19234
rect 26772 19016 26861 19068
rect 26913 19016 27073 19068
rect 27125 19016 27214 19068
rect 26772 18851 27214 19016
rect 26772 18799 26861 18851
rect 26913 18799 27073 18851
rect 27125 18799 27214 18851
rect 26772 18633 27214 18799
rect 26772 18581 26861 18633
rect 26913 18581 27073 18633
rect 27125 18581 27214 18633
rect 26772 18416 27214 18581
rect 26772 18364 26861 18416
rect 26913 18364 27073 18416
rect 27125 18364 27214 18416
rect 26772 18198 27214 18364
rect 26772 18146 26861 18198
rect 26913 18146 27073 18198
rect 27125 18146 27214 18198
rect 26772 17980 27214 18146
rect 26772 17928 26861 17980
rect 26913 17928 27073 17980
rect 27125 17928 27214 17980
rect 26772 17763 27214 17928
rect 26772 17711 26861 17763
rect 26913 17711 27073 17763
rect 27125 17711 27214 17763
rect 26772 17545 27214 17711
rect 26772 17493 26861 17545
rect 26913 17493 27073 17545
rect 27125 17493 27214 17545
rect 26772 17327 27214 17493
rect 26772 17275 26861 17327
rect 26913 17275 27073 17327
rect 27125 17275 27214 17327
rect 26772 17110 27214 17275
rect 26772 17058 26861 17110
rect 26913 17058 27073 17110
rect 27125 17058 27214 17110
rect 26772 16892 27214 17058
rect 26772 16840 26861 16892
rect 26913 16840 27073 16892
rect 27125 16840 27214 16892
rect 26772 16675 27214 16840
rect 26772 16623 26861 16675
rect 26913 16623 27073 16675
rect 27125 16623 27214 16675
rect 26772 16457 27214 16623
rect 26772 16405 26861 16457
rect 26913 16405 27073 16457
rect 27125 16405 27214 16457
rect 26772 16239 27214 16405
rect 26772 16187 26861 16239
rect 26913 16187 27073 16239
rect 27125 16187 27214 16239
rect 26772 16022 27214 16187
rect 26772 15970 26861 16022
rect 26913 15970 27073 16022
rect 27125 15970 27214 16022
rect 26772 15804 27214 15970
rect 26772 15752 26861 15804
rect 26913 15752 27073 15804
rect 27125 15752 27214 15804
rect 26772 15586 27214 15752
rect 26772 15534 26861 15586
rect 26913 15534 27073 15586
rect 27125 15534 27214 15586
rect 26772 15369 27214 15534
rect 26772 15317 26861 15369
rect 26913 15317 27073 15369
rect 27125 15317 27214 15369
rect 26772 15151 27214 15317
rect 26772 15099 26861 15151
rect 26913 15099 27073 15151
rect 27125 15099 27214 15151
rect 26772 14933 27214 15099
rect 26772 14881 26861 14933
rect 26913 14881 27073 14933
rect 27125 14881 27214 14933
rect 26772 14716 27214 14881
rect 26772 14664 26861 14716
rect 26913 14664 27073 14716
rect 27125 14664 27214 14716
rect 26772 14498 27214 14664
rect 26772 14446 26861 14498
rect 26913 14446 27073 14498
rect 27125 14446 27214 14498
rect 26772 14281 27214 14446
rect 26772 14229 26861 14281
rect 26913 14229 27073 14281
rect 27125 14229 27214 14281
rect 26772 14063 27214 14229
rect 26772 14011 26861 14063
rect 26913 14011 27073 14063
rect 27125 14011 27214 14063
rect 26772 13845 27214 14011
rect 26772 13793 26861 13845
rect 26913 13793 27073 13845
rect 27125 13793 27214 13845
rect 26772 13628 27214 13793
rect 26772 13576 26861 13628
rect 26913 13576 27073 13628
rect 27125 13576 27214 13628
rect 26772 13410 27214 13576
rect 26772 13358 26861 13410
rect 26913 13358 27073 13410
rect 27125 13358 27214 13410
rect 26772 13192 27214 13358
rect 26772 13140 26861 13192
rect 26913 13140 27073 13192
rect 27125 13140 27214 13192
rect 26772 12975 27214 13140
rect 26772 12923 26861 12975
rect 26913 12923 27073 12975
rect 27125 12923 27214 12975
rect 26772 12757 27214 12923
rect 26772 12705 26861 12757
rect 26913 12705 27073 12757
rect 27125 12705 27214 12757
rect 26772 12540 27214 12705
rect 26772 12488 26861 12540
rect 26913 12488 27073 12540
rect 27125 12488 27214 12540
rect 26772 12322 27214 12488
rect 26772 12270 26861 12322
rect 26913 12270 27073 12322
rect 27125 12270 27214 12322
rect 26772 12104 27214 12270
rect 26772 12052 26861 12104
rect 26913 12052 27073 12104
rect 27125 12052 27214 12104
rect 26772 11887 27214 12052
rect 26772 11835 26861 11887
rect 26913 11835 27073 11887
rect 27125 11835 27214 11887
rect 26772 11669 27214 11835
rect 26772 11617 26861 11669
rect 26913 11617 27073 11669
rect 27125 11617 27214 11669
rect 26772 11451 27214 11617
rect 26772 11399 26861 11451
rect 26913 11399 27073 11451
rect 27125 11399 27214 11451
rect 26772 11234 27214 11399
rect 26772 11182 26861 11234
rect 26913 11182 27073 11234
rect 27125 11182 27214 11234
rect 26772 11016 27214 11182
rect 26772 10964 26861 11016
rect 26913 10964 27073 11016
rect 27125 10964 27214 11016
rect 26772 10798 27214 10964
rect 26772 10746 26861 10798
rect 26913 10746 27073 10798
rect 27125 10746 27214 10798
rect 26772 10581 27214 10746
rect 26772 10529 26861 10581
rect 26913 10529 27073 10581
rect 27125 10529 27214 10581
rect 26772 10363 27214 10529
rect 26772 10311 26861 10363
rect 26913 10311 27073 10363
rect 27125 10311 27214 10363
rect 26772 10146 27214 10311
rect 26772 10094 26861 10146
rect 26913 10094 27073 10146
rect 27125 10094 27214 10146
rect 26772 9928 27214 10094
rect 26772 9876 26861 9928
rect 26913 9876 27073 9928
rect 27125 9876 27214 9928
rect 26772 9710 27214 9876
rect 26772 9658 26861 9710
rect 26913 9658 27073 9710
rect 27125 9658 27214 9710
rect 26772 9493 27214 9658
rect 26772 9441 26861 9493
rect 26913 9441 27073 9493
rect 27125 9441 27214 9493
rect 26772 9275 27214 9441
rect 26772 9223 26861 9275
rect 26913 9223 27073 9275
rect 27125 9223 27214 9275
rect 26772 9057 27214 9223
rect 26772 9005 26861 9057
rect 26913 9005 27073 9057
rect 27125 9005 27214 9057
rect 26772 8840 27214 9005
rect 26772 8788 26861 8840
rect 26913 8788 27073 8840
rect 27125 8788 27214 8840
rect 26772 8622 27214 8788
rect 26772 8570 26861 8622
rect 26913 8570 27073 8622
rect 27125 8570 27214 8622
rect 26772 8404 27214 8570
rect 26772 8352 26861 8404
rect 26913 8352 27073 8404
rect 27125 8352 27214 8404
rect 26772 8187 27214 8352
rect 26772 8135 26861 8187
rect 26913 8135 27073 8187
rect 27125 8135 27214 8187
rect 26772 7969 27214 8135
rect 26772 7917 26861 7969
rect 26913 7917 27073 7969
rect 27125 7917 27214 7969
rect 26772 7752 27214 7917
rect 26772 7700 26861 7752
rect 26913 7700 27073 7752
rect 27125 7700 27214 7752
rect 26772 7534 27214 7700
rect 26772 7482 26861 7534
rect 26913 7482 27073 7534
rect 27125 7482 27214 7534
rect 26772 7316 27214 7482
rect 26772 7264 26861 7316
rect 26913 7264 27073 7316
rect 27125 7264 27214 7316
rect 26772 7099 27214 7264
rect 26772 7047 26861 7099
rect 26913 7047 27073 7099
rect 27125 7047 27214 7099
rect 26772 6881 27214 7047
rect 26772 6829 26861 6881
rect 26913 6829 27073 6881
rect 27125 6829 27214 6881
rect 26772 6663 27214 6829
rect 26772 6611 26861 6663
rect 26913 6611 27073 6663
rect 27125 6611 27214 6663
rect 26772 6446 27214 6611
rect 26772 6394 26861 6446
rect 26913 6394 27073 6446
rect 27125 6394 27214 6446
rect 26772 6228 27214 6394
rect 26772 6176 26861 6228
rect 26913 6176 27073 6228
rect 27125 6176 27214 6228
rect 26772 6011 27214 6176
rect 26772 5959 26861 6011
rect 26913 5959 27073 6011
rect 27125 5959 27214 6011
rect 26772 5793 27214 5959
rect 26772 5741 26861 5793
rect 26913 5741 27073 5793
rect 27125 5741 27214 5793
rect 26772 5575 27214 5741
rect 26772 5523 26861 5575
rect 26913 5523 27073 5575
rect 27125 5523 27214 5575
rect 26772 5358 27214 5523
rect 26772 5306 26861 5358
rect 26913 5306 27073 5358
rect 27125 5306 27214 5358
rect 26772 4587 27214 5306
rect 26772 4535 26861 4587
rect 26913 4535 27073 4587
rect 27125 4535 27214 4587
rect 26772 4370 27214 4535
rect 26772 4318 26861 4370
rect 26913 4318 27073 4370
rect 27125 4318 27214 4370
rect 26772 4152 27214 4318
rect 26772 4100 26861 4152
rect 26913 4100 27073 4152
rect 27125 4100 27214 4152
rect 26772 3934 27214 4100
rect 26772 3882 26861 3934
rect 26913 3882 27073 3934
rect 27125 3882 27214 3934
rect 26772 3717 27214 3882
rect 26772 3665 26861 3717
rect 26913 3665 27073 3717
rect 27125 3665 27214 3717
rect 26772 1777 27214 3665
rect 27387 33432 27828 34199
rect 27387 33380 27476 33432
rect 27528 33380 27688 33432
rect 27740 33380 27828 33432
rect 27387 33215 27828 33380
rect 27387 33163 27476 33215
rect 27528 33163 27688 33215
rect 27740 33163 27828 33215
rect 27387 32997 27828 33163
rect 27387 32945 27476 32997
rect 27528 32945 27688 32997
rect 27740 32945 27828 32997
rect 27387 32779 27828 32945
rect 27387 32727 27476 32779
rect 27528 32727 27688 32779
rect 27740 32727 27828 32779
rect 27387 32562 27828 32727
rect 27387 32510 27476 32562
rect 27528 32510 27688 32562
rect 27740 32510 27828 32562
rect 27387 32344 27828 32510
rect 27387 32292 27476 32344
rect 27528 32292 27688 32344
rect 27740 32292 27828 32344
rect 27387 32127 27828 32292
rect 27387 32075 27476 32127
rect 27528 32075 27688 32127
rect 27740 32075 27828 32127
rect 27387 31909 27828 32075
rect 27387 31857 27476 31909
rect 27528 31857 27688 31909
rect 27740 31857 27828 31909
rect 27387 31691 27828 31857
rect 27387 31639 27476 31691
rect 27528 31639 27688 31691
rect 27740 31639 27828 31691
rect 27387 31474 27828 31639
rect 27387 31422 27476 31474
rect 27528 31422 27688 31474
rect 27740 31422 27828 31474
rect 27387 31256 27828 31422
rect 27387 31204 27476 31256
rect 27528 31204 27688 31256
rect 27740 31204 27828 31256
rect 27387 31038 27828 31204
rect 27387 30986 27476 31038
rect 27528 30986 27688 31038
rect 27740 30986 27828 31038
rect 27387 30821 27828 30986
rect 27387 30769 27476 30821
rect 27528 30769 27688 30821
rect 27740 30769 27828 30821
rect 27387 30603 27828 30769
rect 27387 30551 27476 30603
rect 27528 30551 27688 30603
rect 27740 30551 27828 30603
rect 27387 30386 27828 30551
rect 27387 30334 27476 30386
rect 27528 30334 27688 30386
rect 27740 30334 27828 30386
rect 27387 30168 27828 30334
rect 27387 30116 27476 30168
rect 27528 30116 27688 30168
rect 27740 30116 27828 30168
rect 27387 29950 27828 30116
rect 27387 29898 27476 29950
rect 27528 29898 27688 29950
rect 27740 29898 27828 29950
rect 27387 29733 27828 29898
rect 27387 29681 27476 29733
rect 27528 29681 27688 29733
rect 27740 29681 27828 29733
rect 27387 29515 27828 29681
rect 27387 29463 27476 29515
rect 27528 29463 27688 29515
rect 27740 29463 27828 29515
rect 27387 29297 27828 29463
rect 27387 29245 27476 29297
rect 27528 29245 27688 29297
rect 27740 29245 27828 29297
rect 27387 29080 27828 29245
rect 27387 29028 27476 29080
rect 27528 29028 27688 29080
rect 27740 29028 27828 29080
rect 27387 28862 27828 29028
rect 27387 28810 27476 28862
rect 27528 28810 27688 28862
rect 27740 28810 27828 28862
rect 27387 28644 27828 28810
rect 27387 28592 27476 28644
rect 27528 28592 27688 28644
rect 27740 28592 27828 28644
rect 27387 28427 27828 28592
rect 27387 28375 27476 28427
rect 27528 28375 27688 28427
rect 27740 28375 27828 28427
rect 27387 28209 27828 28375
rect 27387 28157 27476 28209
rect 27528 28157 27688 28209
rect 27740 28157 27828 28209
rect 27387 27992 27828 28157
rect 27387 27940 27476 27992
rect 27528 27940 27688 27992
rect 27740 27940 27828 27992
rect 27387 27774 27828 27940
rect 27387 27722 27476 27774
rect 27528 27722 27688 27774
rect 27740 27722 27828 27774
rect 27387 27556 27828 27722
rect 27387 27504 27476 27556
rect 27528 27504 27688 27556
rect 27740 27504 27828 27556
rect 27387 27339 27828 27504
rect 27387 27287 27476 27339
rect 27528 27287 27688 27339
rect 27740 27287 27828 27339
rect 27387 27121 27828 27287
rect 27387 27069 27476 27121
rect 27528 27069 27688 27121
rect 27740 27069 27828 27121
rect 27387 26903 27828 27069
rect 27387 26851 27476 26903
rect 27528 26851 27688 26903
rect 27740 26851 27828 26903
rect 27387 26686 27828 26851
rect 27387 26634 27476 26686
rect 27528 26634 27688 26686
rect 27740 26634 27828 26686
rect 27387 26468 27828 26634
rect 27387 26416 27476 26468
rect 27528 26416 27688 26468
rect 27740 26416 27828 26468
rect 27387 26250 27828 26416
rect 27387 26198 27476 26250
rect 27528 26198 27688 26250
rect 27740 26198 27828 26250
rect 27387 26033 27828 26198
rect 27387 25981 27476 26033
rect 27528 25981 27688 26033
rect 27740 25981 27828 26033
rect 27387 25815 27828 25981
rect 27387 25763 27476 25815
rect 27528 25763 27688 25815
rect 27740 25763 27828 25815
rect 27387 25598 27828 25763
rect 27387 25546 27476 25598
rect 27528 25546 27688 25598
rect 27740 25546 27828 25598
rect 27387 25380 27828 25546
rect 27387 25328 27476 25380
rect 27528 25328 27688 25380
rect 27740 25328 27828 25380
rect 27387 25162 27828 25328
rect 27387 25110 27476 25162
rect 27528 25110 27688 25162
rect 27740 25110 27828 25162
rect 27387 24945 27828 25110
rect 27387 24893 27476 24945
rect 27528 24893 27688 24945
rect 27740 24893 27828 24945
rect 27387 24727 27828 24893
rect 27387 24675 27476 24727
rect 27528 24675 27688 24727
rect 27740 24675 27828 24727
rect 27387 24509 27828 24675
rect 27387 24457 27476 24509
rect 27528 24457 27688 24509
rect 27740 24457 27828 24509
rect 27387 24292 27828 24457
rect 27387 24240 27476 24292
rect 27528 24240 27688 24292
rect 27740 24240 27828 24292
rect 27387 24074 27828 24240
rect 27387 24022 27476 24074
rect 27528 24022 27688 24074
rect 27740 24022 27828 24074
rect 27387 23857 27828 24022
rect 27387 23805 27476 23857
rect 27528 23805 27688 23857
rect 27740 23805 27828 23857
rect 27387 23639 27828 23805
rect 27387 23587 27476 23639
rect 27528 23587 27688 23639
rect 27740 23587 27828 23639
rect 27387 23421 27828 23587
rect 27387 23369 27476 23421
rect 27528 23369 27688 23421
rect 27740 23369 27828 23421
rect 27387 23204 27828 23369
rect 27387 23152 27476 23204
rect 27528 23152 27688 23204
rect 27740 23152 27828 23204
rect 27387 22986 27828 23152
rect 27387 22934 27476 22986
rect 27528 22934 27688 22986
rect 27740 22934 27828 22986
rect 27387 22768 27828 22934
rect 27387 22716 27476 22768
rect 27528 22716 27688 22768
rect 27740 22716 27828 22768
rect 27387 22551 27828 22716
rect 27387 22499 27476 22551
rect 27528 22499 27688 22551
rect 27740 22499 27828 22551
rect 27387 22333 27828 22499
rect 27387 22281 27476 22333
rect 27528 22281 27688 22333
rect 27740 22281 27828 22333
rect 27387 22115 27828 22281
rect 27387 22063 27476 22115
rect 27528 22063 27688 22115
rect 27740 22063 27828 22115
rect 27387 21898 27828 22063
rect 27387 21846 27476 21898
rect 27528 21846 27688 21898
rect 27740 21846 27828 21898
rect 27387 21680 27828 21846
rect 27387 21628 27476 21680
rect 27528 21628 27688 21680
rect 27740 21628 27828 21680
rect 27387 21463 27828 21628
rect 27387 21411 27476 21463
rect 27528 21411 27688 21463
rect 27740 21411 27828 21463
rect 27387 21245 27828 21411
rect 27387 21193 27476 21245
rect 27528 21193 27688 21245
rect 27740 21193 27828 21245
rect 27387 21027 27828 21193
rect 27387 20975 27476 21027
rect 27528 20975 27688 21027
rect 27740 20975 27828 21027
rect 27387 20810 27828 20975
rect 27387 20758 27476 20810
rect 27528 20758 27688 20810
rect 27740 20758 27828 20810
rect 27387 20592 27828 20758
rect 27387 20540 27476 20592
rect 27528 20540 27688 20592
rect 27740 20540 27828 20592
rect 27387 20374 27828 20540
rect 27387 20322 27476 20374
rect 27528 20322 27688 20374
rect 27740 20322 27828 20374
rect 27387 20157 27828 20322
rect 27387 20105 27476 20157
rect 27528 20105 27688 20157
rect 27740 20105 27828 20157
rect 27387 19939 27828 20105
rect 27387 19887 27476 19939
rect 27528 19887 27688 19939
rect 27740 19887 27828 19939
rect 27387 19722 27828 19887
rect 27387 19670 27476 19722
rect 27528 19670 27688 19722
rect 27740 19670 27828 19722
rect 27387 19504 27828 19670
rect 27387 19452 27476 19504
rect 27528 19452 27688 19504
rect 27740 19452 27828 19504
rect 27387 19286 27828 19452
rect 27387 19234 27476 19286
rect 27528 19234 27688 19286
rect 27740 19234 27828 19286
rect 27387 19068 27828 19234
rect 27387 19016 27476 19068
rect 27528 19016 27688 19068
rect 27740 19016 27828 19068
rect 27387 18851 27828 19016
rect 27387 18799 27476 18851
rect 27528 18799 27688 18851
rect 27740 18799 27828 18851
rect 27387 18633 27828 18799
rect 27387 18581 27476 18633
rect 27528 18581 27688 18633
rect 27740 18581 27828 18633
rect 27387 18416 27828 18581
rect 27387 18364 27476 18416
rect 27528 18364 27688 18416
rect 27740 18364 27828 18416
rect 27387 18198 27828 18364
rect 27387 18146 27476 18198
rect 27528 18146 27688 18198
rect 27740 18146 27828 18198
rect 27387 17980 27828 18146
rect 27387 17928 27476 17980
rect 27528 17928 27688 17980
rect 27740 17928 27828 17980
rect 27387 17763 27828 17928
rect 27387 17711 27476 17763
rect 27528 17711 27688 17763
rect 27740 17711 27828 17763
rect 27387 17545 27828 17711
rect 27387 17493 27476 17545
rect 27528 17493 27688 17545
rect 27740 17493 27828 17545
rect 27387 17327 27828 17493
rect 27387 17275 27476 17327
rect 27528 17275 27688 17327
rect 27740 17275 27828 17327
rect 27387 17110 27828 17275
rect 27387 17058 27476 17110
rect 27528 17058 27688 17110
rect 27740 17058 27828 17110
rect 27387 16892 27828 17058
rect 27387 16840 27476 16892
rect 27528 16840 27688 16892
rect 27740 16840 27828 16892
rect 27387 16675 27828 16840
rect 27387 16623 27476 16675
rect 27528 16623 27688 16675
rect 27740 16623 27828 16675
rect 27387 16457 27828 16623
rect 27387 16405 27476 16457
rect 27528 16405 27688 16457
rect 27740 16405 27828 16457
rect 27387 16239 27828 16405
rect 27387 16187 27476 16239
rect 27528 16187 27688 16239
rect 27740 16187 27828 16239
rect 27387 16022 27828 16187
rect 27387 15970 27476 16022
rect 27528 15970 27688 16022
rect 27740 15970 27828 16022
rect 27387 15804 27828 15970
rect 27387 15752 27476 15804
rect 27528 15752 27688 15804
rect 27740 15752 27828 15804
rect 27387 15586 27828 15752
rect 27387 15534 27476 15586
rect 27528 15534 27688 15586
rect 27740 15534 27828 15586
rect 27387 15369 27828 15534
rect 27387 15317 27476 15369
rect 27528 15317 27688 15369
rect 27740 15317 27828 15369
rect 27387 15151 27828 15317
rect 27387 15099 27476 15151
rect 27528 15099 27688 15151
rect 27740 15099 27828 15151
rect 27387 14933 27828 15099
rect 27387 14881 27476 14933
rect 27528 14881 27688 14933
rect 27740 14881 27828 14933
rect 27387 14716 27828 14881
rect 27387 14664 27476 14716
rect 27528 14664 27688 14716
rect 27740 14664 27828 14716
rect 27387 14498 27828 14664
rect 27387 14446 27476 14498
rect 27528 14446 27688 14498
rect 27740 14446 27828 14498
rect 27387 14281 27828 14446
rect 27387 14229 27476 14281
rect 27528 14229 27688 14281
rect 27740 14229 27828 14281
rect 27387 14063 27828 14229
rect 27387 14011 27476 14063
rect 27528 14011 27688 14063
rect 27740 14011 27828 14063
rect 27387 13845 27828 14011
rect 27387 13793 27476 13845
rect 27528 13793 27688 13845
rect 27740 13793 27828 13845
rect 27387 13628 27828 13793
rect 27387 13576 27476 13628
rect 27528 13576 27688 13628
rect 27740 13576 27828 13628
rect 27387 13410 27828 13576
rect 27387 13358 27476 13410
rect 27528 13358 27688 13410
rect 27740 13358 27828 13410
rect 27387 13192 27828 13358
rect 27387 13140 27476 13192
rect 27528 13140 27688 13192
rect 27740 13140 27828 13192
rect 27387 12975 27828 13140
rect 27387 12923 27476 12975
rect 27528 12923 27688 12975
rect 27740 12923 27828 12975
rect 27387 12757 27828 12923
rect 27387 12705 27476 12757
rect 27528 12705 27688 12757
rect 27740 12705 27828 12757
rect 27387 12540 27828 12705
rect 27387 12488 27476 12540
rect 27528 12488 27688 12540
rect 27740 12488 27828 12540
rect 27387 12322 27828 12488
rect 27387 12270 27476 12322
rect 27528 12270 27688 12322
rect 27740 12270 27828 12322
rect 27387 12104 27828 12270
rect 27387 12052 27476 12104
rect 27528 12052 27688 12104
rect 27740 12052 27828 12104
rect 27387 11887 27828 12052
rect 27387 11835 27476 11887
rect 27528 11835 27688 11887
rect 27740 11835 27828 11887
rect 27387 11669 27828 11835
rect 27387 11617 27476 11669
rect 27528 11617 27688 11669
rect 27740 11617 27828 11669
rect 27387 11451 27828 11617
rect 27387 11399 27476 11451
rect 27528 11399 27688 11451
rect 27740 11399 27828 11451
rect 27387 11234 27828 11399
rect 27387 11182 27476 11234
rect 27528 11182 27688 11234
rect 27740 11182 27828 11234
rect 27387 11016 27828 11182
rect 27387 10964 27476 11016
rect 27528 10964 27688 11016
rect 27740 10964 27828 11016
rect 27387 10798 27828 10964
rect 27387 10746 27476 10798
rect 27528 10746 27688 10798
rect 27740 10746 27828 10798
rect 27387 10581 27828 10746
rect 27387 10529 27476 10581
rect 27528 10529 27688 10581
rect 27740 10529 27828 10581
rect 27387 10363 27828 10529
rect 27387 10311 27476 10363
rect 27528 10311 27688 10363
rect 27740 10311 27828 10363
rect 27387 10146 27828 10311
rect 27387 10094 27476 10146
rect 27528 10094 27688 10146
rect 27740 10094 27828 10146
rect 27387 9928 27828 10094
rect 27387 9876 27476 9928
rect 27528 9876 27688 9928
rect 27740 9876 27828 9928
rect 27387 9710 27828 9876
rect 27387 9658 27476 9710
rect 27528 9658 27688 9710
rect 27740 9658 27828 9710
rect 27387 9493 27828 9658
rect 27387 9441 27476 9493
rect 27528 9441 27688 9493
rect 27740 9441 27828 9493
rect 27387 9275 27828 9441
rect 27387 9223 27476 9275
rect 27528 9223 27688 9275
rect 27740 9223 27828 9275
rect 27387 9057 27828 9223
rect 27387 9005 27476 9057
rect 27528 9005 27688 9057
rect 27740 9005 27828 9057
rect 27387 8840 27828 9005
rect 27387 8788 27476 8840
rect 27528 8788 27688 8840
rect 27740 8788 27828 8840
rect 27387 8622 27828 8788
rect 27387 8570 27476 8622
rect 27528 8570 27688 8622
rect 27740 8570 27828 8622
rect 27387 8404 27828 8570
rect 27387 8352 27476 8404
rect 27528 8352 27688 8404
rect 27740 8352 27828 8404
rect 27387 8187 27828 8352
rect 27387 8135 27476 8187
rect 27528 8135 27688 8187
rect 27740 8135 27828 8187
rect 27387 7969 27828 8135
rect 27387 7917 27476 7969
rect 27528 7917 27688 7969
rect 27740 7917 27828 7969
rect 27387 7752 27828 7917
rect 27387 7700 27476 7752
rect 27528 7700 27688 7752
rect 27740 7700 27828 7752
rect 27387 7534 27828 7700
rect 27387 7482 27476 7534
rect 27528 7482 27688 7534
rect 27740 7482 27828 7534
rect 27387 7316 27828 7482
rect 27387 7264 27476 7316
rect 27528 7264 27688 7316
rect 27740 7264 27828 7316
rect 27387 7099 27828 7264
rect 27387 7047 27476 7099
rect 27528 7047 27688 7099
rect 27740 7047 27828 7099
rect 27387 6881 27828 7047
rect 27387 6829 27476 6881
rect 27528 6829 27688 6881
rect 27740 6829 27828 6881
rect 27387 6663 27828 6829
rect 27387 6611 27476 6663
rect 27528 6611 27688 6663
rect 27740 6611 27828 6663
rect 27387 6446 27828 6611
rect 27387 6394 27476 6446
rect 27528 6394 27688 6446
rect 27740 6394 27828 6446
rect 27387 6228 27828 6394
rect 57295 33432 57736 34199
rect 57295 33380 57383 33432
rect 57435 33380 57595 33432
rect 57647 33380 57736 33432
rect 57295 33215 57736 33380
rect 57295 33163 57383 33215
rect 57435 33163 57595 33215
rect 57647 33163 57736 33215
rect 57295 32997 57736 33163
rect 57295 32945 57383 32997
rect 57435 32945 57595 32997
rect 57647 32945 57736 32997
rect 57295 32779 57736 32945
rect 57295 32727 57383 32779
rect 57435 32727 57595 32779
rect 57647 32727 57736 32779
rect 57295 32562 57736 32727
rect 57295 32510 57383 32562
rect 57435 32510 57595 32562
rect 57647 32510 57736 32562
rect 57295 32344 57736 32510
rect 57295 32292 57383 32344
rect 57435 32292 57595 32344
rect 57647 32292 57736 32344
rect 57295 32127 57736 32292
rect 57295 32075 57383 32127
rect 57435 32075 57595 32127
rect 57647 32075 57736 32127
rect 57295 31909 57736 32075
rect 57295 31857 57383 31909
rect 57435 31857 57595 31909
rect 57647 31857 57736 31909
rect 57295 31691 57736 31857
rect 57295 31639 57383 31691
rect 57435 31639 57595 31691
rect 57647 31639 57736 31691
rect 57295 31474 57736 31639
rect 57295 31422 57383 31474
rect 57435 31422 57595 31474
rect 57647 31422 57736 31474
rect 57295 31256 57736 31422
rect 57295 31204 57383 31256
rect 57435 31204 57595 31256
rect 57647 31204 57736 31256
rect 57295 31038 57736 31204
rect 57295 30986 57383 31038
rect 57435 30986 57595 31038
rect 57647 30986 57736 31038
rect 57295 30821 57736 30986
rect 57295 30769 57383 30821
rect 57435 30769 57595 30821
rect 57647 30769 57736 30821
rect 57295 30603 57736 30769
rect 57295 30551 57383 30603
rect 57435 30551 57595 30603
rect 57647 30551 57736 30603
rect 57295 30386 57736 30551
rect 57295 30334 57383 30386
rect 57435 30334 57595 30386
rect 57647 30334 57736 30386
rect 57295 30168 57736 30334
rect 57295 30116 57383 30168
rect 57435 30116 57595 30168
rect 57647 30116 57736 30168
rect 57295 29950 57736 30116
rect 57295 29898 57383 29950
rect 57435 29898 57595 29950
rect 57647 29898 57736 29950
rect 57295 29733 57736 29898
rect 57295 29681 57383 29733
rect 57435 29681 57595 29733
rect 57647 29681 57736 29733
rect 57295 29515 57736 29681
rect 57295 29463 57383 29515
rect 57435 29463 57595 29515
rect 57647 29463 57736 29515
rect 57295 29297 57736 29463
rect 57295 29245 57383 29297
rect 57435 29245 57595 29297
rect 57647 29245 57736 29297
rect 57295 29080 57736 29245
rect 57295 29028 57383 29080
rect 57435 29028 57595 29080
rect 57647 29028 57736 29080
rect 57295 28862 57736 29028
rect 57295 28810 57383 28862
rect 57435 28810 57595 28862
rect 57647 28810 57736 28862
rect 57295 28644 57736 28810
rect 57295 28592 57383 28644
rect 57435 28592 57595 28644
rect 57647 28592 57736 28644
rect 57295 28427 57736 28592
rect 57295 28375 57383 28427
rect 57435 28375 57595 28427
rect 57647 28375 57736 28427
rect 57295 28209 57736 28375
rect 57295 28157 57383 28209
rect 57435 28157 57595 28209
rect 57647 28157 57736 28209
rect 57295 27992 57736 28157
rect 57295 27940 57383 27992
rect 57435 27940 57595 27992
rect 57647 27940 57736 27992
rect 57295 27774 57736 27940
rect 57295 27722 57383 27774
rect 57435 27722 57595 27774
rect 57647 27722 57736 27774
rect 57295 27556 57736 27722
rect 57295 27504 57383 27556
rect 57435 27504 57595 27556
rect 57647 27504 57736 27556
rect 57295 27339 57736 27504
rect 57295 27287 57383 27339
rect 57435 27287 57595 27339
rect 57647 27287 57736 27339
rect 57295 27121 57736 27287
rect 57295 27069 57383 27121
rect 57435 27069 57595 27121
rect 57647 27069 57736 27121
rect 57295 26903 57736 27069
rect 57295 26851 57383 26903
rect 57435 26851 57595 26903
rect 57647 26851 57736 26903
rect 57295 26686 57736 26851
rect 57295 26634 57383 26686
rect 57435 26634 57595 26686
rect 57647 26634 57736 26686
rect 57295 26468 57736 26634
rect 57295 26416 57383 26468
rect 57435 26416 57595 26468
rect 57647 26416 57736 26468
rect 57295 26250 57736 26416
rect 57295 26198 57383 26250
rect 57435 26198 57595 26250
rect 57647 26198 57736 26250
rect 57295 26033 57736 26198
rect 57295 25981 57383 26033
rect 57435 25981 57595 26033
rect 57647 25981 57736 26033
rect 57295 25815 57736 25981
rect 57295 25763 57383 25815
rect 57435 25763 57595 25815
rect 57647 25763 57736 25815
rect 57295 25598 57736 25763
rect 57295 25546 57383 25598
rect 57435 25546 57595 25598
rect 57647 25546 57736 25598
rect 57295 25380 57736 25546
rect 57295 25328 57383 25380
rect 57435 25328 57595 25380
rect 57647 25328 57736 25380
rect 57295 25162 57736 25328
rect 57295 25110 57383 25162
rect 57435 25110 57595 25162
rect 57647 25110 57736 25162
rect 57295 24945 57736 25110
rect 57295 24893 57383 24945
rect 57435 24893 57595 24945
rect 57647 24893 57736 24945
rect 57295 24727 57736 24893
rect 57295 24675 57383 24727
rect 57435 24675 57595 24727
rect 57647 24675 57736 24727
rect 57295 24509 57736 24675
rect 57295 24457 57383 24509
rect 57435 24457 57595 24509
rect 57647 24457 57736 24509
rect 57295 24292 57736 24457
rect 57295 24240 57383 24292
rect 57435 24240 57595 24292
rect 57647 24240 57736 24292
rect 57295 24074 57736 24240
rect 57295 24022 57383 24074
rect 57435 24022 57595 24074
rect 57647 24022 57736 24074
rect 57295 23857 57736 24022
rect 57295 23805 57383 23857
rect 57435 23805 57595 23857
rect 57647 23805 57736 23857
rect 57295 23639 57736 23805
rect 57295 23587 57383 23639
rect 57435 23587 57595 23639
rect 57647 23587 57736 23639
rect 57295 23421 57736 23587
rect 57295 23369 57383 23421
rect 57435 23369 57595 23421
rect 57647 23369 57736 23421
rect 57295 23204 57736 23369
rect 57295 23152 57383 23204
rect 57435 23152 57595 23204
rect 57647 23152 57736 23204
rect 57295 22986 57736 23152
rect 57295 22934 57383 22986
rect 57435 22934 57595 22986
rect 57647 22934 57736 22986
rect 57295 22768 57736 22934
rect 57295 22716 57383 22768
rect 57435 22716 57595 22768
rect 57647 22716 57736 22768
rect 57295 22551 57736 22716
rect 57295 22499 57383 22551
rect 57435 22499 57595 22551
rect 57647 22499 57736 22551
rect 57295 22333 57736 22499
rect 57295 22281 57383 22333
rect 57435 22281 57595 22333
rect 57647 22281 57736 22333
rect 57295 22115 57736 22281
rect 57295 22063 57383 22115
rect 57435 22063 57595 22115
rect 57647 22063 57736 22115
rect 57295 21898 57736 22063
rect 57295 21846 57383 21898
rect 57435 21846 57595 21898
rect 57647 21846 57736 21898
rect 57295 21680 57736 21846
rect 57295 21628 57383 21680
rect 57435 21628 57595 21680
rect 57647 21628 57736 21680
rect 57295 21463 57736 21628
rect 57295 21411 57383 21463
rect 57435 21411 57595 21463
rect 57647 21411 57736 21463
rect 57295 21245 57736 21411
rect 57295 21193 57383 21245
rect 57435 21193 57595 21245
rect 57647 21193 57736 21245
rect 57295 21027 57736 21193
rect 57295 20975 57383 21027
rect 57435 20975 57595 21027
rect 57647 20975 57736 21027
rect 57295 20810 57736 20975
rect 57295 20758 57383 20810
rect 57435 20758 57595 20810
rect 57647 20758 57736 20810
rect 57295 20592 57736 20758
rect 57295 20540 57383 20592
rect 57435 20540 57595 20592
rect 57647 20540 57736 20592
rect 57295 20374 57736 20540
rect 57295 20322 57383 20374
rect 57435 20322 57595 20374
rect 57647 20322 57736 20374
rect 57295 20157 57736 20322
rect 57295 20105 57383 20157
rect 57435 20105 57595 20157
rect 57647 20105 57736 20157
rect 57295 19939 57736 20105
rect 57295 19887 57383 19939
rect 57435 19887 57595 19939
rect 57647 19887 57736 19939
rect 57295 19722 57736 19887
rect 57295 19670 57383 19722
rect 57435 19670 57595 19722
rect 57647 19670 57736 19722
rect 57295 19504 57736 19670
rect 57295 19452 57383 19504
rect 57435 19452 57595 19504
rect 57647 19452 57736 19504
rect 57295 19286 57736 19452
rect 57295 19234 57383 19286
rect 57435 19234 57595 19286
rect 57647 19234 57736 19286
rect 57295 19068 57736 19234
rect 57295 19016 57383 19068
rect 57435 19016 57595 19068
rect 57647 19016 57736 19068
rect 57295 18851 57736 19016
rect 57295 18799 57383 18851
rect 57435 18799 57595 18851
rect 57647 18799 57736 18851
rect 57295 18633 57736 18799
rect 57295 18581 57383 18633
rect 57435 18581 57595 18633
rect 57647 18581 57736 18633
rect 57295 18416 57736 18581
rect 57295 18364 57383 18416
rect 57435 18364 57595 18416
rect 57647 18364 57736 18416
rect 57295 18198 57736 18364
rect 57295 18146 57383 18198
rect 57435 18146 57595 18198
rect 57647 18146 57736 18198
rect 57295 17980 57736 18146
rect 57295 17928 57383 17980
rect 57435 17928 57595 17980
rect 57647 17928 57736 17980
rect 57295 17763 57736 17928
rect 57295 17711 57383 17763
rect 57435 17711 57595 17763
rect 57647 17711 57736 17763
rect 57295 17545 57736 17711
rect 57295 17493 57383 17545
rect 57435 17493 57595 17545
rect 57647 17493 57736 17545
rect 57295 17327 57736 17493
rect 57295 17275 57383 17327
rect 57435 17275 57595 17327
rect 57647 17275 57736 17327
rect 57295 17110 57736 17275
rect 57295 17058 57383 17110
rect 57435 17058 57595 17110
rect 57647 17058 57736 17110
rect 57295 16892 57736 17058
rect 57295 16840 57383 16892
rect 57435 16840 57595 16892
rect 57647 16840 57736 16892
rect 57295 16675 57736 16840
rect 57295 16623 57383 16675
rect 57435 16623 57595 16675
rect 57647 16623 57736 16675
rect 57295 16457 57736 16623
rect 57295 16405 57383 16457
rect 57435 16405 57595 16457
rect 57647 16405 57736 16457
rect 57295 16239 57736 16405
rect 57295 16187 57383 16239
rect 57435 16187 57595 16239
rect 57647 16187 57736 16239
rect 57295 16022 57736 16187
rect 57295 15970 57383 16022
rect 57435 15970 57595 16022
rect 57647 15970 57736 16022
rect 57295 15804 57736 15970
rect 57295 15752 57383 15804
rect 57435 15752 57595 15804
rect 57647 15752 57736 15804
rect 57295 15586 57736 15752
rect 57295 15534 57383 15586
rect 57435 15534 57595 15586
rect 57647 15534 57736 15586
rect 57295 15369 57736 15534
rect 57295 15317 57383 15369
rect 57435 15317 57595 15369
rect 57647 15317 57736 15369
rect 57295 15151 57736 15317
rect 57295 15099 57383 15151
rect 57435 15099 57595 15151
rect 57647 15099 57736 15151
rect 57295 14933 57736 15099
rect 57295 14881 57383 14933
rect 57435 14881 57595 14933
rect 57647 14881 57736 14933
rect 57295 14716 57736 14881
rect 57295 14664 57383 14716
rect 57435 14664 57595 14716
rect 57647 14664 57736 14716
rect 57295 14498 57736 14664
rect 57295 14446 57383 14498
rect 57435 14446 57595 14498
rect 57647 14446 57736 14498
rect 57295 14281 57736 14446
rect 57295 14229 57383 14281
rect 57435 14229 57595 14281
rect 57647 14229 57736 14281
rect 57295 14063 57736 14229
rect 57295 14011 57383 14063
rect 57435 14011 57595 14063
rect 57647 14011 57736 14063
rect 57295 13845 57736 14011
rect 57295 13793 57383 13845
rect 57435 13793 57595 13845
rect 57647 13793 57736 13845
rect 57295 13628 57736 13793
rect 57295 13576 57383 13628
rect 57435 13576 57595 13628
rect 57647 13576 57736 13628
rect 57295 13410 57736 13576
rect 57295 13358 57383 13410
rect 57435 13358 57595 13410
rect 57647 13358 57736 13410
rect 57295 13192 57736 13358
rect 57295 13140 57383 13192
rect 57435 13140 57595 13192
rect 57647 13140 57736 13192
rect 57295 12975 57736 13140
rect 57295 12923 57383 12975
rect 57435 12923 57595 12975
rect 57647 12923 57736 12975
rect 57295 12757 57736 12923
rect 57295 12705 57383 12757
rect 57435 12705 57595 12757
rect 57647 12705 57736 12757
rect 57295 12540 57736 12705
rect 57295 12488 57383 12540
rect 57435 12488 57595 12540
rect 57647 12488 57736 12540
rect 57295 12322 57736 12488
rect 57295 12270 57383 12322
rect 57435 12270 57595 12322
rect 57647 12270 57736 12322
rect 57295 12104 57736 12270
rect 57295 12052 57383 12104
rect 57435 12052 57595 12104
rect 57647 12052 57736 12104
rect 57295 11887 57736 12052
rect 57295 11835 57383 11887
rect 57435 11835 57595 11887
rect 57647 11835 57736 11887
rect 57295 11669 57736 11835
rect 57295 11617 57383 11669
rect 57435 11617 57595 11669
rect 57647 11617 57736 11669
rect 57295 11451 57736 11617
rect 57295 11399 57383 11451
rect 57435 11399 57595 11451
rect 57647 11399 57736 11451
rect 57295 11234 57736 11399
rect 57295 11182 57383 11234
rect 57435 11182 57595 11234
rect 57647 11182 57736 11234
rect 57295 11016 57736 11182
rect 57295 10964 57383 11016
rect 57435 10964 57595 11016
rect 57647 10964 57736 11016
rect 57295 10798 57736 10964
rect 57295 10746 57383 10798
rect 57435 10746 57595 10798
rect 57647 10746 57736 10798
rect 57295 10581 57736 10746
rect 57295 10529 57383 10581
rect 57435 10529 57595 10581
rect 57647 10529 57736 10581
rect 57295 10363 57736 10529
rect 57295 10311 57383 10363
rect 57435 10311 57595 10363
rect 57647 10311 57736 10363
rect 57295 10146 57736 10311
rect 57295 10094 57383 10146
rect 57435 10094 57595 10146
rect 57647 10094 57736 10146
rect 57295 9928 57736 10094
rect 57295 9876 57383 9928
rect 57435 9876 57595 9928
rect 57647 9876 57736 9928
rect 57295 9710 57736 9876
rect 57295 9658 57383 9710
rect 57435 9658 57595 9710
rect 57647 9658 57736 9710
rect 57295 9493 57736 9658
rect 57295 9441 57383 9493
rect 57435 9441 57595 9493
rect 57647 9441 57736 9493
rect 57295 9275 57736 9441
rect 57295 9223 57383 9275
rect 57435 9223 57595 9275
rect 57647 9223 57736 9275
rect 57295 9057 57736 9223
rect 57295 9005 57383 9057
rect 57435 9005 57595 9057
rect 57647 9005 57736 9057
rect 57295 8840 57736 9005
rect 57295 8788 57383 8840
rect 57435 8788 57595 8840
rect 57647 8788 57736 8840
rect 57295 8622 57736 8788
rect 57295 8570 57383 8622
rect 57435 8570 57595 8622
rect 57647 8570 57736 8622
rect 57295 8404 57736 8570
rect 57295 8352 57383 8404
rect 57435 8352 57595 8404
rect 57647 8352 57736 8404
rect 57295 8187 57736 8352
rect 57295 8135 57383 8187
rect 57435 8135 57595 8187
rect 57647 8135 57736 8187
rect 57295 7969 57736 8135
rect 57295 7917 57383 7969
rect 57435 7917 57595 7969
rect 57647 7917 57736 7969
rect 57295 7752 57736 7917
rect 57295 7700 57383 7752
rect 57435 7700 57595 7752
rect 57647 7700 57736 7752
rect 57295 7534 57736 7700
rect 57295 7482 57383 7534
rect 57435 7482 57595 7534
rect 57647 7482 57736 7534
rect 57295 7316 57736 7482
rect 57295 7264 57383 7316
rect 57435 7264 57595 7316
rect 57647 7264 57736 7316
rect 57295 7099 57736 7264
rect 57295 7047 57383 7099
rect 57435 7047 57595 7099
rect 57647 7047 57736 7099
rect 57295 6881 57736 7047
rect 57295 6829 57383 6881
rect 57435 6829 57595 6881
rect 57647 6829 57736 6881
rect 57295 6663 57736 6829
rect 57295 6611 57383 6663
rect 57435 6611 57595 6663
rect 57647 6611 57736 6663
rect 57295 6446 57736 6611
rect 57295 6394 57383 6446
rect 57435 6394 57595 6446
rect 57647 6394 57736 6446
rect 49896 6349 50076 6361
rect 49896 6347 49908 6349
rect 49728 6301 49908 6347
rect 49896 6297 49908 6301
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 27387 6176 27476 6228
rect 27528 6176 27688 6228
rect 27740 6176 27828 6228
rect 27387 6011 27828 6176
rect 27387 5959 27476 6011
rect 27528 5959 27688 6011
rect 27740 5959 27828 6011
rect 27387 5793 27828 5959
rect 27387 5741 27476 5793
rect 27528 5741 27688 5793
rect 27740 5741 27828 5793
rect 27387 5575 27828 5741
rect 27387 5523 27476 5575
rect 27528 5523 27688 5575
rect 27740 5523 27828 5575
rect 27387 5358 27828 5523
rect 27387 5306 27476 5358
rect 27528 5306 27688 5358
rect 27740 5306 27828 5358
rect 27387 4587 27828 5306
rect 57295 6228 57736 6394
rect 57295 6176 57383 6228
rect 57435 6176 57595 6228
rect 57647 6176 57736 6228
rect 57295 6011 57736 6176
rect 57295 5959 57383 6011
rect 57435 5959 57595 6011
rect 57647 5959 57736 6011
rect 57295 5793 57736 5959
rect 57295 5741 57383 5793
rect 57435 5741 57595 5793
rect 57647 5741 57736 5793
rect 57295 5575 57736 5741
rect 57295 5523 57383 5575
rect 57435 5523 57595 5575
rect 57647 5523 57736 5575
rect 57295 5358 57736 5523
rect 57295 5306 57383 5358
rect 57435 5306 57595 5358
rect 57647 5306 57736 5358
rect 51642 5199 51822 5211
rect 51642 5196 51654 5199
rect 49963 5150 51654 5196
rect 51642 5147 51654 5150
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 27387 4535 27476 4587
rect 27528 4535 27688 4587
rect 27740 4535 27828 4587
rect 27387 4370 27828 4535
rect 27387 4318 27476 4370
rect 27528 4318 27688 4370
rect 27740 4318 27828 4370
rect 27387 4152 27828 4318
rect 27387 4100 27476 4152
rect 27528 4100 27688 4152
rect 27740 4100 27828 4152
rect 27387 3934 27828 4100
rect 27387 3882 27476 3934
rect 27528 3882 27688 3934
rect 27740 3882 27828 3934
rect 57295 4587 57736 5306
rect 57295 4535 57383 4587
rect 57435 4535 57595 4587
rect 57647 4535 57736 4587
rect 57295 4370 57736 4535
rect 57295 4318 57383 4370
rect 57435 4318 57595 4370
rect 57647 4318 57736 4370
rect 57295 4152 57736 4318
rect 57295 4100 57383 4152
rect 57435 4100 57595 4152
rect 57647 4100 57736 4152
rect 57295 3934 57736 4100
rect 27387 3717 27828 3882
rect 27387 3665 27476 3717
rect 27528 3665 27688 3717
rect 27740 3665 27828 3717
rect 27387 1925 27828 3665
rect 28628 3906 40180 3917
rect 28628 3860 28639 3906
rect 28685 3860 28755 3906
rect 28801 3860 28871 3906
rect 28917 3860 28987 3906
rect 29033 3860 29103 3906
rect 29149 3860 29219 3906
rect 29265 3860 29335 3906
rect 29381 3860 29451 3906
rect 29497 3860 29567 3906
rect 29613 3860 29683 3906
rect 29729 3860 29799 3906
rect 29845 3860 29915 3906
rect 29961 3860 30031 3906
rect 30077 3860 30147 3906
rect 30193 3860 30263 3906
rect 30309 3860 30379 3906
rect 30425 3860 30495 3906
rect 30541 3860 30611 3906
rect 30657 3860 30727 3906
rect 30773 3860 30843 3906
rect 30889 3860 30959 3906
rect 31005 3860 31075 3906
rect 31121 3860 31191 3906
rect 31237 3860 31307 3906
rect 31353 3860 31423 3906
rect 31469 3860 31539 3906
rect 31585 3860 31655 3906
rect 31701 3860 31771 3906
rect 31817 3860 31887 3906
rect 31933 3860 32003 3906
rect 32049 3860 32119 3906
rect 32165 3860 32235 3906
rect 32281 3860 32351 3906
rect 32397 3860 32467 3906
rect 32513 3860 32583 3906
rect 32629 3860 32699 3906
rect 32745 3860 32815 3906
rect 32861 3860 32931 3906
rect 32977 3860 33047 3906
rect 33093 3860 33163 3906
rect 33209 3860 33279 3906
rect 33325 3860 33395 3906
rect 33441 3860 33511 3906
rect 33557 3860 33627 3906
rect 33673 3860 33743 3906
rect 33789 3860 33859 3906
rect 33905 3860 33975 3906
rect 34021 3860 34091 3906
rect 34137 3860 34207 3906
rect 34253 3860 34323 3906
rect 34369 3860 34439 3906
rect 34485 3860 34555 3906
rect 34601 3860 34671 3906
rect 34717 3860 34787 3906
rect 34833 3860 34903 3906
rect 34949 3860 35019 3906
rect 35065 3860 35135 3906
rect 35181 3860 35251 3906
rect 35297 3860 35367 3906
rect 35413 3860 35483 3906
rect 35529 3860 35599 3906
rect 35645 3860 35715 3906
rect 35761 3860 35831 3906
rect 35877 3860 35947 3906
rect 35993 3860 36063 3906
rect 36109 3860 36179 3906
rect 36225 3860 36295 3906
rect 36341 3860 36411 3906
rect 36457 3860 36527 3906
rect 36573 3860 36643 3906
rect 36689 3860 36759 3906
rect 36805 3860 36875 3906
rect 36921 3860 36991 3906
rect 37037 3860 37107 3906
rect 37153 3860 37223 3906
rect 37269 3860 37339 3906
rect 37385 3860 37455 3906
rect 37501 3860 37571 3906
rect 37617 3860 37687 3906
rect 37733 3860 37803 3906
rect 37849 3860 37919 3906
rect 37965 3860 38035 3906
rect 38081 3860 38151 3906
rect 38197 3860 38267 3906
rect 38313 3860 38383 3906
rect 38429 3860 38499 3906
rect 38545 3860 38615 3906
rect 38661 3860 38731 3906
rect 38777 3860 38847 3906
rect 38893 3860 38963 3906
rect 39009 3860 39079 3906
rect 39125 3860 39195 3906
rect 39241 3860 39311 3906
rect 39357 3860 39427 3906
rect 39473 3860 39543 3906
rect 39589 3860 39659 3906
rect 39705 3860 39775 3906
rect 39821 3860 39891 3906
rect 39937 3860 40007 3906
rect 40053 3860 40123 3906
rect 40169 3860 40180 3906
rect 28628 3790 40180 3860
rect 28628 3744 28639 3790
rect 28685 3744 28755 3790
rect 28801 3744 28871 3790
rect 28917 3744 28987 3790
rect 29033 3744 29103 3790
rect 29149 3744 29219 3790
rect 29265 3744 29335 3790
rect 29381 3744 29451 3790
rect 29497 3744 29567 3790
rect 29613 3744 29683 3790
rect 29729 3744 29799 3790
rect 29845 3744 29915 3790
rect 29961 3744 30031 3790
rect 30077 3744 30147 3790
rect 30193 3744 30263 3790
rect 30309 3744 30379 3790
rect 30425 3744 30495 3790
rect 30541 3744 30611 3790
rect 30657 3744 30727 3790
rect 30773 3744 30843 3790
rect 30889 3744 30959 3790
rect 31005 3744 31075 3790
rect 31121 3744 31191 3790
rect 31237 3744 31307 3790
rect 31353 3744 31423 3790
rect 31469 3744 31539 3790
rect 31585 3744 31655 3790
rect 31701 3744 31771 3790
rect 31817 3744 31887 3790
rect 31933 3744 32003 3790
rect 32049 3744 32119 3790
rect 32165 3744 32235 3790
rect 32281 3744 32351 3790
rect 32397 3744 32467 3790
rect 32513 3744 32583 3790
rect 32629 3744 32699 3790
rect 32745 3744 32815 3790
rect 32861 3744 32931 3790
rect 32977 3744 33047 3790
rect 33093 3744 33163 3790
rect 33209 3744 33279 3790
rect 33325 3744 33395 3790
rect 33441 3744 33511 3790
rect 33557 3744 33627 3790
rect 33673 3744 33743 3790
rect 33789 3744 33859 3790
rect 33905 3744 33975 3790
rect 34021 3744 34091 3790
rect 34137 3744 34207 3790
rect 34253 3744 34323 3790
rect 34369 3744 34439 3790
rect 34485 3744 34555 3790
rect 34601 3744 34671 3790
rect 34717 3744 34787 3790
rect 34833 3744 34903 3790
rect 34949 3744 35019 3790
rect 35065 3744 35135 3790
rect 35181 3744 35251 3790
rect 35297 3744 35367 3790
rect 35413 3744 35483 3790
rect 35529 3744 35599 3790
rect 35645 3744 35715 3790
rect 35761 3744 35831 3790
rect 35877 3744 35947 3790
rect 35993 3744 36063 3790
rect 36109 3744 36179 3790
rect 36225 3744 36295 3790
rect 36341 3744 36411 3790
rect 36457 3744 36527 3790
rect 36573 3744 36643 3790
rect 36689 3744 36759 3790
rect 36805 3744 36875 3790
rect 36921 3744 36991 3790
rect 37037 3744 37107 3790
rect 37153 3744 37223 3790
rect 37269 3744 37339 3790
rect 37385 3744 37455 3790
rect 37501 3744 37571 3790
rect 37617 3744 37687 3790
rect 37733 3744 37803 3790
rect 37849 3744 37919 3790
rect 37965 3744 38035 3790
rect 38081 3744 38151 3790
rect 38197 3744 38267 3790
rect 38313 3744 38383 3790
rect 38429 3744 38499 3790
rect 38545 3744 38615 3790
rect 38661 3744 38731 3790
rect 38777 3744 38847 3790
rect 38893 3744 38963 3790
rect 39009 3744 39079 3790
rect 39125 3744 39195 3790
rect 39241 3744 39311 3790
rect 39357 3744 39427 3790
rect 39473 3744 39543 3790
rect 39589 3744 39659 3790
rect 39705 3744 39775 3790
rect 39821 3744 39891 3790
rect 39937 3744 40007 3790
rect 40053 3744 40123 3790
rect 40169 3744 40180 3790
rect 28628 3674 40180 3744
rect 28628 3628 28639 3674
rect 28685 3628 28755 3674
rect 28801 3628 28871 3674
rect 28917 3628 28987 3674
rect 29033 3628 29103 3674
rect 29149 3628 29219 3674
rect 29265 3628 29335 3674
rect 29381 3628 29451 3674
rect 29497 3628 29567 3674
rect 29613 3628 29683 3674
rect 29729 3628 29799 3674
rect 29845 3628 29915 3674
rect 29961 3628 30031 3674
rect 30077 3628 30147 3674
rect 30193 3628 30263 3674
rect 30309 3628 30379 3674
rect 30425 3628 30495 3674
rect 30541 3628 30611 3674
rect 30657 3628 30727 3674
rect 30773 3628 30843 3674
rect 30889 3628 30959 3674
rect 31005 3628 31075 3674
rect 31121 3628 31191 3674
rect 31237 3628 31307 3674
rect 31353 3628 31423 3674
rect 31469 3628 31539 3674
rect 31585 3628 31655 3674
rect 31701 3628 31771 3674
rect 31817 3628 31887 3674
rect 31933 3628 32003 3674
rect 32049 3628 32119 3674
rect 32165 3628 32235 3674
rect 32281 3628 32351 3674
rect 32397 3628 32467 3674
rect 32513 3628 32583 3674
rect 32629 3628 32699 3674
rect 32745 3628 32815 3674
rect 32861 3628 32931 3674
rect 32977 3628 33047 3674
rect 33093 3628 33163 3674
rect 33209 3628 33279 3674
rect 33325 3628 33395 3674
rect 33441 3628 33511 3674
rect 33557 3628 33627 3674
rect 33673 3628 33743 3674
rect 33789 3628 33859 3674
rect 33905 3628 33975 3674
rect 34021 3628 34091 3674
rect 34137 3628 34207 3674
rect 34253 3628 34323 3674
rect 34369 3628 34439 3674
rect 34485 3628 34555 3674
rect 34601 3628 34671 3674
rect 34717 3628 34787 3674
rect 34833 3628 34903 3674
rect 34949 3628 35019 3674
rect 35065 3628 35135 3674
rect 35181 3628 35251 3674
rect 35297 3628 35367 3674
rect 35413 3628 35483 3674
rect 35529 3628 35599 3674
rect 35645 3628 35715 3674
rect 35761 3628 35831 3674
rect 35877 3628 35947 3674
rect 35993 3628 36063 3674
rect 36109 3628 36179 3674
rect 36225 3628 36295 3674
rect 36341 3628 36411 3674
rect 36457 3628 36527 3674
rect 36573 3628 36643 3674
rect 36689 3628 36759 3674
rect 36805 3628 36875 3674
rect 36921 3628 36991 3674
rect 37037 3628 37107 3674
rect 37153 3628 37223 3674
rect 37269 3628 37339 3674
rect 37385 3628 37455 3674
rect 37501 3628 37571 3674
rect 37617 3628 37687 3674
rect 37733 3628 37803 3674
rect 37849 3628 37919 3674
rect 37965 3628 38035 3674
rect 38081 3628 38151 3674
rect 38197 3628 38267 3674
rect 38313 3628 38383 3674
rect 38429 3628 38499 3674
rect 38545 3628 38615 3674
rect 38661 3628 38731 3674
rect 38777 3628 38847 3674
rect 38893 3628 38963 3674
rect 39009 3628 39079 3674
rect 39125 3628 39195 3674
rect 39241 3628 39311 3674
rect 39357 3628 39427 3674
rect 39473 3628 39543 3674
rect 39589 3628 39659 3674
rect 39705 3628 39775 3674
rect 39821 3628 39891 3674
rect 39937 3628 40007 3674
rect 40053 3628 40123 3674
rect 40169 3628 40180 3674
rect 28628 3558 40180 3628
rect 28628 3512 28639 3558
rect 28685 3512 28755 3558
rect 28801 3512 28871 3558
rect 28917 3512 28987 3558
rect 29033 3512 29103 3558
rect 29149 3512 29219 3558
rect 29265 3512 29335 3558
rect 29381 3512 29451 3558
rect 29497 3512 29567 3558
rect 29613 3512 29683 3558
rect 29729 3512 29799 3558
rect 29845 3512 29915 3558
rect 29961 3512 30031 3558
rect 30077 3512 30147 3558
rect 30193 3512 30263 3558
rect 30309 3512 30379 3558
rect 30425 3512 30495 3558
rect 30541 3512 30611 3558
rect 30657 3512 30727 3558
rect 30773 3512 30843 3558
rect 30889 3512 30959 3558
rect 31005 3512 31075 3558
rect 31121 3512 31191 3558
rect 31237 3512 31307 3558
rect 31353 3512 31423 3558
rect 31469 3512 31539 3558
rect 31585 3512 31655 3558
rect 31701 3512 31771 3558
rect 31817 3512 31887 3558
rect 31933 3512 32003 3558
rect 32049 3512 32119 3558
rect 32165 3512 32235 3558
rect 32281 3512 32351 3558
rect 32397 3512 32467 3558
rect 32513 3512 32583 3558
rect 32629 3512 32699 3558
rect 32745 3512 32815 3558
rect 32861 3512 32931 3558
rect 32977 3512 33047 3558
rect 33093 3512 33163 3558
rect 33209 3512 33279 3558
rect 33325 3512 33395 3558
rect 33441 3512 33511 3558
rect 33557 3512 33627 3558
rect 33673 3512 33743 3558
rect 33789 3512 33859 3558
rect 33905 3512 33975 3558
rect 34021 3512 34091 3558
rect 34137 3512 34207 3558
rect 34253 3512 34323 3558
rect 34369 3512 34439 3558
rect 34485 3512 34555 3558
rect 34601 3512 34671 3558
rect 34717 3512 34787 3558
rect 34833 3512 34903 3558
rect 34949 3512 35019 3558
rect 35065 3512 35135 3558
rect 35181 3512 35251 3558
rect 35297 3512 35367 3558
rect 35413 3512 35483 3558
rect 35529 3512 35599 3558
rect 35645 3512 35715 3558
rect 35761 3512 35831 3558
rect 35877 3512 35947 3558
rect 35993 3512 36063 3558
rect 36109 3512 36179 3558
rect 36225 3512 36295 3558
rect 36341 3512 36411 3558
rect 36457 3512 36527 3558
rect 36573 3512 36643 3558
rect 36689 3512 36759 3558
rect 36805 3512 36875 3558
rect 36921 3512 36991 3558
rect 37037 3512 37107 3558
rect 37153 3512 37223 3558
rect 37269 3512 37339 3558
rect 37385 3512 37455 3558
rect 37501 3512 37571 3558
rect 37617 3512 37687 3558
rect 37733 3512 37803 3558
rect 37849 3512 37919 3558
rect 37965 3512 38035 3558
rect 38081 3512 38151 3558
rect 38197 3512 38267 3558
rect 38313 3512 38383 3558
rect 38429 3512 38499 3558
rect 38545 3512 38615 3558
rect 38661 3512 38731 3558
rect 38777 3512 38847 3558
rect 38893 3512 38963 3558
rect 39009 3512 39079 3558
rect 39125 3512 39195 3558
rect 39241 3512 39311 3558
rect 39357 3512 39427 3558
rect 39473 3512 39543 3558
rect 39589 3512 39659 3558
rect 39705 3512 39775 3558
rect 39821 3512 39891 3558
rect 39937 3512 40007 3558
rect 40053 3512 40123 3558
rect 40169 3512 40180 3558
rect 28628 3442 40180 3512
rect 28628 3396 28639 3442
rect 28685 3396 28755 3442
rect 28801 3396 28871 3442
rect 28917 3396 28987 3442
rect 29033 3396 29103 3442
rect 29149 3396 29219 3442
rect 29265 3396 29335 3442
rect 29381 3396 29451 3442
rect 29497 3396 29567 3442
rect 29613 3396 29683 3442
rect 29729 3396 29799 3442
rect 29845 3396 29915 3442
rect 29961 3396 30031 3442
rect 30077 3396 30147 3442
rect 30193 3396 30263 3442
rect 30309 3396 30379 3442
rect 30425 3396 30495 3442
rect 30541 3396 30611 3442
rect 30657 3396 30727 3442
rect 30773 3396 30843 3442
rect 30889 3396 30959 3442
rect 31005 3396 31075 3442
rect 31121 3396 31191 3442
rect 31237 3396 31307 3442
rect 31353 3396 31423 3442
rect 31469 3396 31539 3442
rect 31585 3396 31655 3442
rect 31701 3396 31771 3442
rect 31817 3396 31887 3442
rect 31933 3396 32003 3442
rect 32049 3396 32119 3442
rect 32165 3396 32235 3442
rect 32281 3396 32351 3442
rect 32397 3396 32467 3442
rect 32513 3396 32583 3442
rect 32629 3396 32699 3442
rect 32745 3396 32815 3442
rect 32861 3396 32931 3442
rect 32977 3396 33047 3442
rect 33093 3396 33163 3442
rect 33209 3396 33279 3442
rect 33325 3396 33395 3442
rect 33441 3396 33511 3442
rect 33557 3396 33627 3442
rect 33673 3396 33743 3442
rect 33789 3396 33859 3442
rect 33905 3396 33975 3442
rect 34021 3396 34091 3442
rect 34137 3396 34207 3442
rect 34253 3396 34323 3442
rect 34369 3396 34439 3442
rect 34485 3396 34555 3442
rect 34601 3396 34671 3442
rect 34717 3396 34787 3442
rect 34833 3396 34903 3442
rect 34949 3396 35019 3442
rect 35065 3396 35135 3442
rect 35181 3396 35251 3442
rect 35297 3396 35367 3442
rect 35413 3396 35483 3442
rect 35529 3396 35599 3442
rect 35645 3396 35715 3442
rect 35761 3396 35831 3442
rect 35877 3396 35947 3442
rect 35993 3396 36063 3442
rect 36109 3396 36179 3442
rect 36225 3396 36295 3442
rect 36341 3396 36411 3442
rect 36457 3396 36527 3442
rect 36573 3396 36643 3442
rect 36689 3396 36759 3442
rect 36805 3396 36875 3442
rect 36921 3396 36991 3442
rect 37037 3396 37107 3442
rect 37153 3396 37223 3442
rect 37269 3396 37339 3442
rect 37385 3396 37455 3442
rect 37501 3396 37571 3442
rect 37617 3396 37687 3442
rect 37733 3396 37803 3442
rect 37849 3396 37919 3442
rect 37965 3396 38035 3442
rect 38081 3396 38151 3442
rect 38197 3396 38267 3442
rect 38313 3396 38383 3442
rect 38429 3396 38499 3442
rect 38545 3396 38615 3442
rect 38661 3396 38731 3442
rect 38777 3396 38847 3442
rect 38893 3396 38963 3442
rect 39009 3396 39079 3442
rect 39125 3396 39195 3442
rect 39241 3396 39311 3442
rect 39357 3396 39427 3442
rect 39473 3396 39543 3442
rect 39589 3396 39659 3442
rect 39705 3396 39775 3442
rect 39821 3396 39891 3442
rect 39937 3396 40007 3442
rect 40053 3396 40123 3442
rect 40169 3396 40180 3442
rect 28628 3326 40180 3396
rect 28628 3280 28639 3326
rect 28685 3280 28755 3326
rect 28801 3280 28871 3326
rect 28917 3280 28987 3326
rect 29033 3280 29103 3326
rect 29149 3280 29219 3326
rect 29265 3280 29335 3326
rect 29381 3280 29451 3326
rect 29497 3280 29567 3326
rect 29613 3280 29683 3326
rect 29729 3280 29799 3326
rect 29845 3280 29915 3326
rect 29961 3280 30031 3326
rect 30077 3280 30147 3326
rect 30193 3280 30263 3326
rect 30309 3280 30379 3326
rect 30425 3280 30495 3326
rect 30541 3280 30611 3326
rect 30657 3280 30727 3326
rect 30773 3280 30843 3326
rect 30889 3280 30959 3326
rect 31005 3280 31075 3326
rect 31121 3280 31191 3326
rect 31237 3280 31307 3326
rect 31353 3280 31423 3326
rect 31469 3280 31539 3326
rect 31585 3280 31655 3326
rect 31701 3280 31771 3326
rect 31817 3280 31887 3326
rect 31933 3280 32003 3326
rect 32049 3280 32119 3326
rect 32165 3280 32235 3326
rect 32281 3280 32351 3326
rect 32397 3280 32467 3326
rect 32513 3280 32583 3326
rect 32629 3280 32699 3326
rect 32745 3280 32815 3326
rect 32861 3280 32931 3326
rect 32977 3280 33047 3326
rect 33093 3280 33163 3326
rect 33209 3280 33279 3326
rect 33325 3280 33395 3326
rect 33441 3280 33511 3326
rect 33557 3280 33627 3326
rect 33673 3280 33743 3326
rect 33789 3280 33859 3326
rect 33905 3280 33975 3326
rect 34021 3280 34091 3326
rect 34137 3280 34207 3326
rect 34253 3280 34323 3326
rect 34369 3280 34439 3326
rect 34485 3280 34555 3326
rect 34601 3280 34671 3326
rect 34717 3280 34787 3326
rect 34833 3280 34903 3326
rect 34949 3280 35019 3326
rect 35065 3280 35135 3326
rect 35181 3280 35251 3326
rect 35297 3280 35367 3326
rect 35413 3280 35483 3326
rect 35529 3280 35599 3326
rect 35645 3280 35715 3326
rect 35761 3280 35831 3326
rect 35877 3280 35947 3326
rect 35993 3280 36063 3326
rect 36109 3280 36179 3326
rect 36225 3280 36295 3326
rect 36341 3280 36411 3326
rect 36457 3280 36527 3326
rect 36573 3280 36643 3326
rect 36689 3280 36759 3326
rect 36805 3280 36875 3326
rect 36921 3280 36991 3326
rect 37037 3280 37107 3326
rect 37153 3280 37223 3326
rect 37269 3280 37339 3326
rect 37385 3280 37455 3326
rect 37501 3280 37571 3326
rect 37617 3280 37687 3326
rect 37733 3280 37803 3326
rect 37849 3280 37919 3326
rect 37965 3280 38035 3326
rect 38081 3280 38151 3326
rect 38197 3280 38267 3326
rect 38313 3280 38383 3326
rect 38429 3280 38499 3326
rect 38545 3280 38615 3326
rect 38661 3280 38731 3326
rect 38777 3280 38847 3326
rect 38893 3280 38963 3326
rect 39009 3280 39079 3326
rect 39125 3280 39195 3326
rect 39241 3280 39311 3326
rect 39357 3280 39427 3326
rect 39473 3280 39543 3326
rect 39589 3280 39659 3326
rect 39705 3280 39775 3326
rect 39821 3280 39891 3326
rect 39937 3280 40007 3326
rect 40053 3280 40123 3326
rect 40169 3280 40180 3326
rect 50834 3906 56586 3917
rect 50834 3860 50845 3906
rect 50891 3860 50961 3906
rect 51007 3860 51077 3906
rect 51123 3860 51193 3906
rect 51239 3860 51309 3906
rect 51355 3860 51425 3906
rect 51471 3860 51541 3906
rect 51587 3860 51657 3906
rect 51703 3860 51773 3906
rect 51819 3860 51889 3906
rect 51935 3860 52005 3906
rect 52051 3860 52121 3906
rect 52167 3860 52237 3906
rect 52283 3860 52353 3906
rect 52399 3860 52469 3906
rect 52515 3860 52585 3906
rect 52631 3860 52701 3906
rect 52747 3860 52817 3906
rect 52863 3860 52933 3906
rect 52979 3860 53049 3906
rect 53095 3860 53165 3906
rect 53211 3860 53281 3906
rect 53327 3860 53397 3906
rect 53443 3860 53513 3906
rect 53559 3860 53629 3906
rect 53675 3860 53745 3906
rect 53791 3860 53861 3906
rect 53907 3860 53977 3906
rect 54023 3860 54093 3906
rect 54139 3860 54209 3906
rect 54255 3860 54325 3906
rect 54371 3860 54441 3906
rect 54487 3860 54557 3906
rect 54603 3860 54673 3906
rect 54719 3860 54789 3906
rect 54835 3860 54905 3906
rect 54951 3860 55021 3906
rect 55067 3860 55137 3906
rect 55183 3860 55253 3906
rect 55299 3860 55369 3906
rect 55415 3860 55485 3906
rect 55531 3860 55601 3906
rect 55647 3860 55717 3906
rect 55763 3860 55833 3906
rect 55879 3860 55949 3906
rect 55995 3860 56065 3906
rect 56111 3860 56181 3906
rect 56227 3860 56297 3906
rect 56343 3860 56413 3906
rect 56459 3860 56529 3906
rect 56575 3860 56586 3906
rect 50834 3790 56586 3860
rect 50834 3744 50845 3790
rect 50891 3744 50961 3790
rect 51007 3744 51077 3790
rect 51123 3744 51193 3790
rect 51239 3744 51309 3790
rect 51355 3744 51425 3790
rect 51471 3744 51541 3790
rect 51587 3744 51657 3790
rect 51703 3744 51773 3790
rect 51819 3744 51889 3790
rect 51935 3744 52005 3790
rect 52051 3744 52121 3790
rect 52167 3744 52237 3790
rect 52283 3744 52353 3790
rect 52399 3744 52469 3790
rect 52515 3744 52585 3790
rect 52631 3744 52701 3790
rect 52747 3744 52817 3790
rect 52863 3744 52933 3790
rect 52979 3744 53049 3790
rect 53095 3744 53165 3790
rect 53211 3744 53281 3790
rect 53327 3744 53397 3790
rect 53443 3744 53513 3790
rect 53559 3744 53629 3790
rect 53675 3744 53745 3790
rect 53791 3744 53861 3790
rect 53907 3744 53977 3790
rect 54023 3744 54093 3790
rect 54139 3744 54209 3790
rect 54255 3744 54325 3790
rect 54371 3744 54441 3790
rect 54487 3744 54557 3790
rect 54603 3744 54673 3790
rect 54719 3744 54789 3790
rect 54835 3744 54905 3790
rect 54951 3744 55021 3790
rect 55067 3744 55137 3790
rect 55183 3744 55253 3790
rect 55299 3744 55369 3790
rect 55415 3744 55485 3790
rect 55531 3744 55601 3790
rect 55647 3744 55717 3790
rect 55763 3744 55833 3790
rect 55879 3744 55949 3790
rect 55995 3744 56065 3790
rect 56111 3744 56181 3790
rect 56227 3744 56297 3790
rect 56343 3744 56413 3790
rect 56459 3744 56529 3790
rect 56575 3744 56586 3790
rect 50834 3674 56586 3744
rect 50834 3628 50845 3674
rect 50891 3628 50961 3674
rect 51007 3628 51077 3674
rect 51123 3628 51193 3674
rect 51239 3628 51309 3674
rect 51355 3628 51425 3674
rect 51471 3628 51541 3674
rect 51587 3628 51657 3674
rect 51703 3628 51773 3674
rect 51819 3628 51889 3674
rect 51935 3628 52005 3674
rect 52051 3628 52121 3674
rect 52167 3628 52237 3674
rect 52283 3628 52353 3674
rect 52399 3628 52469 3674
rect 52515 3628 52585 3674
rect 52631 3628 52701 3674
rect 52747 3628 52817 3674
rect 52863 3628 52933 3674
rect 52979 3628 53049 3674
rect 53095 3628 53165 3674
rect 53211 3628 53281 3674
rect 53327 3628 53397 3674
rect 53443 3628 53513 3674
rect 53559 3628 53629 3674
rect 53675 3628 53745 3674
rect 53791 3628 53861 3674
rect 53907 3628 53977 3674
rect 54023 3628 54093 3674
rect 54139 3628 54209 3674
rect 54255 3628 54325 3674
rect 54371 3628 54441 3674
rect 54487 3628 54557 3674
rect 54603 3628 54673 3674
rect 54719 3628 54789 3674
rect 54835 3628 54905 3674
rect 54951 3628 55021 3674
rect 55067 3628 55137 3674
rect 55183 3628 55253 3674
rect 55299 3628 55369 3674
rect 55415 3628 55485 3674
rect 55531 3628 55601 3674
rect 55647 3628 55717 3674
rect 55763 3628 55833 3674
rect 55879 3628 55949 3674
rect 55995 3628 56065 3674
rect 56111 3628 56181 3674
rect 56227 3628 56297 3674
rect 56343 3628 56413 3674
rect 56459 3628 56529 3674
rect 56575 3628 56586 3674
rect 50834 3558 56586 3628
rect 50834 3512 50845 3558
rect 50891 3512 50961 3558
rect 51007 3512 51077 3558
rect 51123 3512 51193 3558
rect 51239 3512 51309 3558
rect 51355 3512 51425 3558
rect 51471 3512 51541 3558
rect 51587 3512 51657 3558
rect 51703 3512 51773 3558
rect 51819 3512 51889 3558
rect 51935 3512 52005 3558
rect 52051 3512 52121 3558
rect 52167 3512 52237 3558
rect 52283 3512 52353 3558
rect 52399 3512 52469 3558
rect 52515 3512 52585 3558
rect 52631 3512 52701 3558
rect 52747 3512 52817 3558
rect 52863 3512 52933 3558
rect 52979 3512 53049 3558
rect 53095 3512 53165 3558
rect 53211 3512 53281 3558
rect 53327 3512 53397 3558
rect 53443 3512 53513 3558
rect 53559 3512 53629 3558
rect 53675 3512 53745 3558
rect 53791 3512 53861 3558
rect 53907 3512 53977 3558
rect 54023 3512 54093 3558
rect 54139 3512 54209 3558
rect 54255 3512 54325 3558
rect 54371 3512 54441 3558
rect 54487 3512 54557 3558
rect 54603 3512 54673 3558
rect 54719 3512 54789 3558
rect 54835 3512 54905 3558
rect 54951 3512 55021 3558
rect 55067 3512 55137 3558
rect 55183 3512 55253 3558
rect 55299 3512 55369 3558
rect 55415 3512 55485 3558
rect 55531 3512 55601 3558
rect 55647 3512 55717 3558
rect 55763 3512 55833 3558
rect 55879 3512 55949 3558
rect 55995 3512 56065 3558
rect 56111 3512 56181 3558
rect 56227 3512 56297 3558
rect 56343 3512 56413 3558
rect 56459 3512 56529 3558
rect 56575 3512 56586 3558
rect 50834 3442 56586 3512
rect 50834 3396 50845 3442
rect 50891 3396 50961 3442
rect 51007 3396 51077 3442
rect 51123 3396 51193 3442
rect 51239 3396 51309 3442
rect 51355 3396 51425 3442
rect 51471 3396 51541 3442
rect 51587 3396 51657 3442
rect 51703 3396 51773 3442
rect 51819 3396 51889 3442
rect 51935 3396 52005 3442
rect 52051 3396 52121 3442
rect 52167 3396 52237 3442
rect 52283 3396 52353 3442
rect 52399 3396 52469 3442
rect 52515 3396 52585 3442
rect 52631 3396 52701 3442
rect 52747 3396 52817 3442
rect 52863 3396 52933 3442
rect 52979 3396 53049 3442
rect 53095 3396 53165 3442
rect 53211 3396 53281 3442
rect 53327 3396 53397 3442
rect 53443 3396 53513 3442
rect 53559 3396 53629 3442
rect 53675 3396 53745 3442
rect 53791 3396 53861 3442
rect 53907 3396 53977 3442
rect 54023 3396 54093 3442
rect 54139 3396 54209 3442
rect 54255 3396 54325 3442
rect 54371 3396 54441 3442
rect 54487 3396 54557 3442
rect 54603 3396 54673 3442
rect 54719 3396 54789 3442
rect 54835 3396 54905 3442
rect 54951 3396 55021 3442
rect 55067 3396 55137 3442
rect 55183 3396 55253 3442
rect 55299 3396 55369 3442
rect 55415 3396 55485 3442
rect 55531 3396 55601 3442
rect 55647 3396 55717 3442
rect 55763 3396 55833 3442
rect 55879 3396 55949 3442
rect 55995 3396 56065 3442
rect 56111 3396 56181 3442
rect 56227 3396 56297 3442
rect 56343 3396 56413 3442
rect 56459 3396 56529 3442
rect 56575 3396 56586 3442
rect 50834 3326 56586 3396
rect 28628 3210 40180 3280
rect 40611 3282 40791 3294
rect 40611 3230 40623 3282
rect 40779 3230 40791 3282
rect 40611 3218 40791 3230
rect 50834 3280 50845 3326
rect 50891 3280 50961 3326
rect 51007 3280 51077 3326
rect 51123 3280 51193 3326
rect 51239 3280 51309 3326
rect 51355 3280 51425 3326
rect 51471 3280 51541 3326
rect 51587 3280 51657 3326
rect 51703 3280 51773 3326
rect 51819 3280 51889 3326
rect 51935 3280 52005 3326
rect 52051 3280 52121 3326
rect 52167 3280 52237 3326
rect 52283 3280 52353 3326
rect 52399 3280 52469 3326
rect 52515 3280 52585 3326
rect 52631 3280 52701 3326
rect 52747 3280 52817 3326
rect 52863 3280 52933 3326
rect 52979 3280 53049 3326
rect 53095 3280 53165 3326
rect 53211 3280 53281 3326
rect 53327 3280 53397 3326
rect 53443 3280 53513 3326
rect 53559 3280 53629 3326
rect 53675 3280 53745 3326
rect 53791 3280 53861 3326
rect 53907 3280 53977 3326
rect 54023 3280 54093 3326
rect 54139 3280 54209 3326
rect 54255 3280 54325 3326
rect 54371 3280 54441 3326
rect 54487 3280 54557 3326
rect 54603 3280 54673 3326
rect 54719 3280 54789 3326
rect 54835 3280 54905 3326
rect 54951 3280 55021 3326
rect 55067 3280 55137 3326
rect 55183 3280 55253 3326
rect 55299 3280 55369 3326
rect 55415 3280 55485 3326
rect 55531 3280 55601 3326
rect 55647 3280 55717 3326
rect 55763 3280 55833 3326
rect 55879 3280 55949 3326
rect 55995 3280 56065 3326
rect 56111 3280 56181 3326
rect 56227 3280 56297 3326
rect 56343 3280 56413 3326
rect 56459 3280 56529 3326
rect 56575 3280 56586 3326
rect 28628 3164 28639 3210
rect 28685 3164 28755 3210
rect 28801 3164 28871 3210
rect 28917 3164 28987 3210
rect 29033 3164 29103 3210
rect 29149 3164 29219 3210
rect 29265 3164 29335 3210
rect 29381 3164 29451 3210
rect 29497 3164 29567 3210
rect 29613 3164 29683 3210
rect 29729 3164 29799 3210
rect 29845 3164 29915 3210
rect 29961 3164 30031 3210
rect 30077 3164 30147 3210
rect 30193 3164 30263 3210
rect 30309 3164 30379 3210
rect 30425 3164 30495 3210
rect 30541 3164 30611 3210
rect 30657 3164 30727 3210
rect 30773 3164 30843 3210
rect 30889 3164 30959 3210
rect 31005 3164 31075 3210
rect 31121 3164 31191 3210
rect 31237 3164 31307 3210
rect 31353 3164 31423 3210
rect 31469 3164 31539 3210
rect 31585 3164 31655 3210
rect 31701 3164 31771 3210
rect 31817 3164 31887 3210
rect 31933 3164 32003 3210
rect 32049 3164 32119 3210
rect 32165 3164 32235 3210
rect 32281 3164 32351 3210
rect 32397 3164 32467 3210
rect 32513 3164 32583 3210
rect 32629 3164 32699 3210
rect 32745 3164 32815 3210
rect 32861 3164 32931 3210
rect 32977 3164 33047 3210
rect 33093 3164 33163 3210
rect 33209 3164 33279 3210
rect 33325 3164 33395 3210
rect 33441 3164 33511 3210
rect 33557 3164 33627 3210
rect 33673 3164 33743 3210
rect 33789 3164 33859 3210
rect 33905 3164 33975 3210
rect 34021 3164 34091 3210
rect 34137 3164 34207 3210
rect 34253 3164 34323 3210
rect 34369 3164 34439 3210
rect 34485 3164 34555 3210
rect 34601 3164 34671 3210
rect 34717 3164 34787 3210
rect 34833 3164 34903 3210
rect 34949 3164 35019 3210
rect 35065 3164 35135 3210
rect 35181 3164 35251 3210
rect 35297 3164 35367 3210
rect 35413 3164 35483 3210
rect 35529 3164 35599 3210
rect 35645 3164 35715 3210
rect 35761 3164 35831 3210
rect 35877 3164 35947 3210
rect 35993 3164 36063 3210
rect 36109 3164 36179 3210
rect 36225 3164 36295 3210
rect 36341 3164 36411 3210
rect 36457 3164 36527 3210
rect 36573 3164 36643 3210
rect 36689 3164 36759 3210
rect 36805 3164 36875 3210
rect 36921 3164 36991 3210
rect 37037 3164 37107 3210
rect 37153 3164 37223 3210
rect 37269 3164 37339 3210
rect 37385 3164 37455 3210
rect 37501 3164 37571 3210
rect 37617 3164 37687 3210
rect 37733 3164 37803 3210
rect 37849 3164 37919 3210
rect 37965 3164 38035 3210
rect 38081 3164 38151 3210
rect 38197 3164 38267 3210
rect 38313 3164 38383 3210
rect 38429 3164 38499 3210
rect 38545 3164 38615 3210
rect 38661 3164 38731 3210
rect 38777 3164 38847 3210
rect 38893 3164 38963 3210
rect 39009 3164 39079 3210
rect 39125 3164 39195 3210
rect 39241 3164 39311 3210
rect 39357 3164 39427 3210
rect 39473 3164 39543 3210
rect 39589 3164 39659 3210
rect 39705 3164 39775 3210
rect 39821 3164 39891 3210
rect 39937 3164 40007 3210
rect 40053 3164 40123 3210
rect 40169 3164 40180 3210
rect 28628 3094 40180 3164
rect 28628 3048 28639 3094
rect 28685 3048 28755 3094
rect 28801 3048 28871 3094
rect 28917 3048 28987 3094
rect 29033 3048 29103 3094
rect 29149 3048 29219 3094
rect 29265 3048 29335 3094
rect 29381 3048 29451 3094
rect 29497 3048 29567 3094
rect 29613 3048 29683 3094
rect 29729 3048 29799 3094
rect 29845 3048 29915 3094
rect 29961 3048 30031 3094
rect 30077 3048 30147 3094
rect 30193 3048 30263 3094
rect 30309 3048 30379 3094
rect 30425 3048 30495 3094
rect 30541 3048 30611 3094
rect 30657 3048 30727 3094
rect 30773 3048 30843 3094
rect 30889 3048 30959 3094
rect 31005 3048 31075 3094
rect 31121 3048 31191 3094
rect 31237 3048 31307 3094
rect 31353 3048 31423 3094
rect 31469 3048 31539 3094
rect 31585 3048 31655 3094
rect 31701 3048 31771 3094
rect 31817 3048 31887 3094
rect 31933 3048 32003 3094
rect 32049 3048 32119 3094
rect 32165 3048 32235 3094
rect 32281 3048 32351 3094
rect 32397 3048 32467 3094
rect 32513 3048 32583 3094
rect 32629 3048 32699 3094
rect 32745 3048 32815 3094
rect 32861 3048 32931 3094
rect 32977 3048 33047 3094
rect 33093 3048 33163 3094
rect 33209 3048 33279 3094
rect 33325 3048 33395 3094
rect 33441 3048 33511 3094
rect 33557 3048 33627 3094
rect 33673 3048 33743 3094
rect 33789 3048 33859 3094
rect 33905 3048 33975 3094
rect 34021 3048 34091 3094
rect 34137 3048 34207 3094
rect 34253 3048 34323 3094
rect 34369 3048 34439 3094
rect 34485 3048 34555 3094
rect 34601 3048 34671 3094
rect 34717 3048 34787 3094
rect 34833 3048 34903 3094
rect 34949 3048 35019 3094
rect 35065 3048 35135 3094
rect 35181 3048 35251 3094
rect 35297 3048 35367 3094
rect 35413 3048 35483 3094
rect 35529 3048 35599 3094
rect 35645 3048 35715 3094
rect 35761 3048 35831 3094
rect 35877 3048 35947 3094
rect 35993 3048 36063 3094
rect 36109 3048 36179 3094
rect 36225 3048 36295 3094
rect 36341 3048 36411 3094
rect 36457 3048 36527 3094
rect 36573 3048 36643 3094
rect 36689 3048 36759 3094
rect 36805 3048 36875 3094
rect 36921 3048 36991 3094
rect 37037 3048 37107 3094
rect 37153 3048 37223 3094
rect 37269 3048 37339 3094
rect 37385 3048 37455 3094
rect 37501 3048 37571 3094
rect 37617 3048 37687 3094
rect 37733 3048 37803 3094
rect 37849 3048 37919 3094
rect 37965 3048 38035 3094
rect 38081 3048 38151 3094
rect 38197 3048 38267 3094
rect 38313 3048 38383 3094
rect 38429 3048 38499 3094
rect 38545 3048 38615 3094
rect 38661 3048 38731 3094
rect 38777 3048 38847 3094
rect 38893 3048 38963 3094
rect 39009 3048 39079 3094
rect 39125 3048 39195 3094
rect 39241 3048 39311 3094
rect 39357 3048 39427 3094
rect 39473 3048 39543 3094
rect 39589 3048 39659 3094
rect 39705 3048 39775 3094
rect 39821 3048 39891 3094
rect 39937 3048 40007 3094
rect 40053 3048 40123 3094
rect 40169 3048 40180 3094
rect 28628 2978 40180 3048
rect 28628 2932 28639 2978
rect 28685 2932 28755 2978
rect 28801 2932 28871 2978
rect 28917 2932 28987 2978
rect 29033 2932 29103 2978
rect 29149 2932 29219 2978
rect 29265 2932 29335 2978
rect 29381 2932 29451 2978
rect 29497 2932 29567 2978
rect 29613 2932 29683 2978
rect 29729 2932 29799 2978
rect 29845 2932 29915 2978
rect 29961 2932 30031 2978
rect 30077 2932 30147 2978
rect 30193 2932 30263 2978
rect 30309 2932 30379 2978
rect 30425 2932 30495 2978
rect 30541 2932 30611 2978
rect 30657 2932 30727 2978
rect 30773 2932 30843 2978
rect 30889 2932 30959 2978
rect 31005 2932 31075 2978
rect 31121 2932 31191 2978
rect 31237 2932 31307 2978
rect 31353 2932 31423 2978
rect 31469 2932 31539 2978
rect 31585 2932 31655 2978
rect 31701 2932 31771 2978
rect 31817 2932 31887 2978
rect 31933 2932 32003 2978
rect 32049 2932 32119 2978
rect 32165 2932 32235 2978
rect 32281 2932 32351 2978
rect 32397 2932 32467 2978
rect 32513 2932 32583 2978
rect 32629 2932 32699 2978
rect 32745 2932 32815 2978
rect 32861 2932 32931 2978
rect 32977 2932 33047 2978
rect 33093 2932 33163 2978
rect 33209 2932 33279 2978
rect 33325 2932 33395 2978
rect 33441 2932 33511 2978
rect 33557 2932 33627 2978
rect 33673 2932 33743 2978
rect 33789 2932 33859 2978
rect 33905 2932 33975 2978
rect 34021 2932 34091 2978
rect 34137 2932 34207 2978
rect 34253 2932 34323 2978
rect 34369 2932 34439 2978
rect 34485 2932 34555 2978
rect 34601 2932 34671 2978
rect 34717 2932 34787 2978
rect 34833 2932 34903 2978
rect 34949 2932 35019 2978
rect 35065 2932 35135 2978
rect 35181 2932 35251 2978
rect 35297 2932 35367 2978
rect 35413 2932 35483 2978
rect 35529 2932 35599 2978
rect 35645 2932 35715 2978
rect 35761 2932 35831 2978
rect 35877 2932 35947 2978
rect 35993 2932 36063 2978
rect 36109 2932 36179 2978
rect 36225 2932 36295 2978
rect 36341 2932 36411 2978
rect 36457 2932 36527 2978
rect 36573 2932 36643 2978
rect 36689 2932 36759 2978
rect 36805 2932 36875 2978
rect 36921 2932 36991 2978
rect 37037 2932 37107 2978
rect 37153 2932 37223 2978
rect 37269 2932 37339 2978
rect 37385 2932 37455 2978
rect 37501 2932 37571 2978
rect 37617 2932 37687 2978
rect 37733 2932 37803 2978
rect 37849 2932 37919 2978
rect 37965 2932 38035 2978
rect 38081 2932 38151 2978
rect 38197 2932 38267 2978
rect 38313 2932 38383 2978
rect 38429 2932 38499 2978
rect 38545 2932 38615 2978
rect 38661 2932 38731 2978
rect 38777 2932 38847 2978
rect 38893 2932 38963 2978
rect 39009 2932 39079 2978
rect 39125 2932 39195 2978
rect 39241 2932 39311 2978
rect 39357 2932 39427 2978
rect 39473 2932 39543 2978
rect 39589 2932 39659 2978
rect 39705 2932 39775 2978
rect 39821 2932 39891 2978
rect 39937 2932 40007 2978
rect 40053 2932 40123 2978
rect 40169 2932 40180 2978
rect 28628 2862 40180 2932
rect 28628 2816 28639 2862
rect 28685 2816 28755 2862
rect 28801 2816 28871 2862
rect 28917 2816 28987 2862
rect 29033 2816 29103 2862
rect 29149 2816 29219 2862
rect 29265 2816 29335 2862
rect 29381 2816 29451 2862
rect 29497 2816 29567 2862
rect 29613 2816 29683 2862
rect 29729 2816 29799 2862
rect 29845 2816 29915 2862
rect 29961 2816 30031 2862
rect 30077 2816 30147 2862
rect 30193 2816 30263 2862
rect 30309 2816 30379 2862
rect 30425 2816 30495 2862
rect 30541 2816 30611 2862
rect 30657 2816 30727 2862
rect 30773 2816 30843 2862
rect 30889 2816 30959 2862
rect 31005 2816 31075 2862
rect 31121 2816 31191 2862
rect 31237 2816 31307 2862
rect 31353 2816 31423 2862
rect 31469 2816 31539 2862
rect 31585 2816 31655 2862
rect 31701 2816 31771 2862
rect 31817 2816 31887 2862
rect 31933 2816 32003 2862
rect 32049 2816 32119 2862
rect 32165 2816 32235 2862
rect 32281 2816 32351 2862
rect 32397 2816 32467 2862
rect 32513 2816 32583 2862
rect 32629 2816 32699 2862
rect 32745 2816 32815 2862
rect 32861 2816 32931 2862
rect 32977 2816 33047 2862
rect 33093 2816 33163 2862
rect 33209 2816 33279 2862
rect 33325 2816 33395 2862
rect 33441 2816 33511 2862
rect 33557 2816 33627 2862
rect 33673 2816 33743 2862
rect 33789 2816 33859 2862
rect 33905 2816 33975 2862
rect 34021 2816 34091 2862
rect 34137 2816 34207 2862
rect 34253 2816 34323 2862
rect 34369 2816 34439 2862
rect 34485 2816 34555 2862
rect 34601 2816 34671 2862
rect 34717 2816 34787 2862
rect 34833 2816 34903 2862
rect 34949 2816 35019 2862
rect 35065 2816 35135 2862
rect 35181 2816 35251 2862
rect 35297 2816 35367 2862
rect 35413 2816 35483 2862
rect 35529 2816 35599 2862
rect 35645 2816 35715 2862
rect 35761 2816 35831 2862
rect 35877 2816 35947 2862
rect 35993 2816 36063 2862
rect 36109 2816 36179 2862
rect 36225 2816 36295 2862
rect 36341 2816 36411 2862
rect 36457 2816 36527 2862
rect 36573 2816 36643 2862
rect 36689 2816 36759 2862
rect 36805 2816 36875 2862
rect 36921 2816 36991 2862
rect 37037 2816 37107 2862
rect 37153 2816 37223 2862
rect 37269 2816 37339 2862
rect 37385 2816 37455 2862
rect 37501 2816 37571 2862
rect 37617 2816 37687 2862
rect 37733 2816 37803 2862
rect 37849 2816 37919 2862
rect 37965 2816 38035 2862
rect 38081 2816 38151 2862
rect 38197 2816 38267 2862
rect 38313 2816 38383 2862
rect 38429 2816 38499 2862
rect 38545 2816 38615 2862
rect 38661 2816 38731 2862
rect 38777 2816 38847 2862
rect 38893 2816 38963 2862
rect 39009 2816 39079 2862
rect 39125 2816 39195 2862
rect 39241 2816 39311 2862
rect 39357 2816 39427 2862
rect 39473 2816 39543 2862
rect 39589 2816 39659 2862
rect 39705 2816 39775 2862
rect 39821 2816 39891 2862
rect 39937 2816 40007 2862
rect 40053 2816 40123 2862
rect 40169 2816 40180 2862
rect 28628 2746 40180 2816
rect 28628 2700 28639 2746
rect 28685 2700 28755 2746
rect 28801 2700 28871 2746
rect 28917 2700 28987 2746
rect 29033 2700 29103 2746
rect 29149 2700 29219 2746
rect 29265 2700 29335 2746
rect 29381 2700 29451 2746
rect 29497 2700 29567 2746
rect 29613 2700 29683 2746
rect 29729 2700 29799 2746
rect 29845 2700 29915 2746
rect 29961 2700 30031 2746
rect 30077 2700 30147 2746
rect 30193 2700 30263 2746
rect 30309 2700 30379 2746
rect 30425 2700 30495 2746
rect 30541 2700 30611 2746
rect 30657 2700 30727 2746
rect 30773 2700 30843 2746
rect 30889 2700 30959 2746
rect 31005 2700 31075 2746
rect 31121 2700 31191 2746
rect 31237 2700 31307 2746
rect 31353 2700 31423 2746
rect 31469 2700 31539 2746
rect 31585 2700 31655 2746
rect 31701 2700 31771 2746
rect 31817 2700 31887 2746
rect 31933 2700 32003 2746
rect 32049 2700 32119 2746
rect 32165 2700 32235 2746
rect 32281 2700 32351 2746
rect 32397 2700 32467 2746
rect 32513 2700 32583 2746
rect 32629 2700 32699 2746
rect 32745 2700 32815 2746
rect 32861 2700 32931 2746
rect 32977 2700 33047 2746
rect 33093 2700 33163 2746
rect 33209 2700 33279 2746
rect 33325 2700 33395 2746
rect 33441 2700 33511 2746
rect 33557 2700 33627 2746
rect 33673 2700 33743 2746
rect 33789 2700 33859 2746
rect 33905 2700 33975 2746
rect 34021 2700 34091 2746
rect 34137 2700 34207 2746
rect 34253 2700 34323 2746
rect 34369 2700 34439 2746
rect 34485 2700 34555 2746
rect 34601 2700 34671 2746
rect 34717 2700 34787 2746
rect 34833 2700 34903 2746
rect 34949 2700 35019 2746
rect 35065 2700 35135 2746
rect 35181 2700 35251 2746
rect 35297 2700 35367 2746
rect 35413 2700 35483 2746
rect 35529 2700 35599 2746
rect 35645 2700 35715 2746
rect 35761 2700 35831 2746
rect 35877 2700 35947 2746
rect 35993 2700 36063 2746
rect 36109 2700 36179 2746
rect 36225 2700 36295 2746
rect 36341 2700 36411 2746
rect 36457 2700 36527 2746
rect 36573 2700 36643 2746
rect 36689 2700 36759 2746
rect 36805 2700 36875 2746
rect 36921 2700 36991 2746
rect 37037 2700 37107 2746
rect 37153 2700 37223 2746
rect 37269 2700 37339 2746
rect 37385 2700 37455 2746
rect 37501 2700 37571 2746
rect 37617 2700 37687 2746
rect 37733 2700 37803 2746
rect 37849 2700 37919 2746
rect 37965 2700 38035 2746
rect 38081 2700 38151 2746
rect 38197 2700 38267 2746
rect 38313 2700 38383 2746
rect 38429 2700 38499 2746
rect 38545 2700 38615 2746
rect 38661 2700 38731 2746
rect 38777 2700 38847 2746
rect 38893 2700 38963 2746
rect 39009 2700 39079 2746
rect 39125 2700 39195 2746
rect 39241 2700 39311 2746
rect 39357 2700 39427 2746
rect 39473 2700 39543 2746
rect 39589 2700 39659 2746
rect 39705 2700 39775 2746
rect 39821 2700 39891 2746
rect 39937 2700 40007 2746
rect 40053 2700 40123 2746
rect 40169 2700 40180 2746
rect 28628 2630 40180 2700
rect 28628 2584 28639 2630
rect 28685 2584 28755 2630
rect 28801 2584 28871 2630
rect 28917 2584 28987 2630
rect 29033 2584 29103 2630
rect 29149 2584 29219 2630
rect 29265 2584 29335 2630
rect 29381 2584 29451 2630
rect 29497 2584 29567 2630
rect 29613 2584 29683 2630
rect 29729 2584 29799 2630
rect 29845 2584 29915 2630
rect 29961 2584 30031 2630
rect 30077 2584 30147 2630
rect 30193 2584 30263 2630
rect 30309 2584 30379 2630
rect 30425 2584 30495 2630
rect 30541 2584 30611 2630
rect 30657 2584 30727 2630
rect 30773 2584 30843 2630
rect 30889 2584 30959 2630
rect 31005 2584 31075 2630
rect 31121 2584 31191 2630
rect 31237 2584 31307 2630
rect 31353 2584 31423 2630
rect 31469 2584 31539 2630
rect 31585 2584 31655 2630
rect 31701 2584 31771 2630
rect 31817 2584 31887 2630
rect 31933 2584 32003 2630
rect 32049 2584 32119 2630
rect 32165 2584 32235 2630
rect 32281 2584 32351 2630
rect 32397 2584 32467 2630
rect 32513 2584 32583 2630
rect 32629 2584 32699 2630
rect 32745 2584 32815 2630
rect 32861 2584 32931 2630
rect 32977 2584 33047 2630
rect 33093 2584 33163 2630
rect 33209 2584 33279 2630
rect 33325 2584 33395 2630
rect 33441 2584 33511 2630
rect 33557 2584 33627 2630
rect 33673 2584 33743 2630
rect 33789 2584 33859 2630
rect 33905 2584 33975 2630
rect 34021 2584 34091 2630
rect 34137 2584 34207 2630
rect 34253 2584 34323 2630
rect 34369 2584 34439 2630
rect 34485 2584 34555 2630
rect 34601 2584 34671 2630
rect 34717 2584 34787 2630
rect 34833 2584 34903 2630
rect 34949 2584 35019 2630
rect 35065 2584 35135 2630
rect 35181 2584 35251 2630
rect 35297 2584 35367 2630
rect 35413 2584 35483 2630
rect 35529 2584 35599 2630
rect 35645 2584 35715 2630
rect 35761 2584 35831 2630
rect 35877 2584 35947 2630
rect 35993 2584 36063 2630
rect 36109 2584 36179 2630
rect 36225 2584 36295 2630
rect 36341 2584 36411 2630
rect 36457 2584 36527 2630
rect 36573 2584 36643 2630
rect 36689 2584 36759 2630
rect 36805 2584 36875 2630
rect 36921 2584 36991 2630
rect 37037 2584 37107 2630
rect 37153 2584 37223 2630
rect 37269 2584 37339 2630
rect 37385 2584 37455 2630
rect 37501 2584 37571 2630
rect 37617 2584 37687 2630
rect 37733 2584 37803 2630
rect 37849 2584 37919 2630
rect 37965 2584 38035 2630
rect 38081 2584 38151 2630
rect 38197 2584 38267 2630
rect 38313 2584 38383 2630
rect 38429 2584 38499 2630
rect 38545 2584 38615 2630
rect 38661 2584 38731 2630
rect 38777 2584 38847 2630
rect 38893 2584 38963 2630
rect 39009 2584 39079 2630
rect 39125 2584 39195 2630
rect 39241 2584 39311 2630
rect 39357 2584 39427 2630
rect 39473 2584 39543 2630
rect 39589 2584 39659 2630
rect 39705 2584 39775 2630
rect 39821 2584 39891 2630
rect 39937 2584 40007 2630
rect 40053 2584 40123 2630
rect 40169 2584 40180 2630
rect 28628 2514 40180 2584
rect 28628 2468 28639 2514
rect 28685 2468 28755 2514
rect 28801 2468 28871 2514
rect 28917 2468 28987 2514
rect 29033 2468 29103 2514
rect 29149 2468 29219 2514
rect 29265 2468 29335 2514
rect 29381 2468 29451 2514
rect 29497 2468 29567 2514
rect 29613 2468 29683 2514
rect 29729 2468 29799 2514
rect 29845 2468 29915 2514
rect 29961 2468 30031 2514
rect 30077 2468 30147 2514
rect 30193 2468 30263 2514
rect 30309 2468 30379 2514
rect 30425 2468 30495 2514
rect 30541 2468 30611 2514
rect 30657 2468 30727 2514
rect 30773 2468 30843 2514
rect 30889 2468 30959 2514
rect 31005 2468 31075 2514
rect 31121 2468 31191 2514
rect 31237 2468 31307 2514
rect 31353 2468 31423 2514
rect 31469 2468 31539 2514
rect 31585 2468 31655 2514
rect 31701 2468 31771 2514
rect 31817 2468 31887 2514
rect 31933 2468 32003 2514
rect 32049 2468 32119 2514
rect 32165 2468 32235 2514
rect 32281 2468 32351 2514
rect 32397 2468 32467 2514
rect 32513 2468 32583 2514
rect 32629 2468 32699 2514
rect 32745 2468 32815 2514
rect 32861 2468 32931 2514
rect 32977 2468 33047 2514
rect 33093 2468 33163 2514
rect 33209 2468 33279 2514
rect 33325 2468 33395 2514
rect 33441 2468 33511 2514
rect 33557 2468 33627 2514
rect 33673 2468 33743 2514
rect 33789 2468 33859 2514
rect 33905 2468 33975 2514
rect 34021 2468 34091 2514
rect 34137 2468 34207 2514
rect 34253 2468 34323 2514
rect 34369 2468 34439 2514
rect 34485 2468 34555 2514
rect 34601 2468 34671 2514
rect 34717 2468 34787 2514
rect 34833 2468 34903 2514
rect 34949 2468 35019 2514
rect 35065 2468 35135 2514
rect 35181 2468 35251 2514
rect 35297 2468 35367 2514
rect 35413 2468 35483 2514
rect 35529 2468 35599 2514
rect 35645 2468 35715 2514
rect 35761 2468 35831 2514
rect 35877 2468 35947 2514
rect 35993 2468 36063 2514
rect 36109 2468 36179 2514
rect 36225 2468 36295 2514
rect 36341 2468 36411 2514
rect 36457 2468 36527 2514
rect 36573 2468 36643 2514
rect 36689 2468 36759 2514
rect 36805 2468 36875 2514
rect 36921 2468 36991 2514
rect 37037 2468 37107 2514
rect 37153 2468 37223 2514
rect 37269 2468 37339 2514
rect 37385 2468 37455 2514
rect 37501 2468 37571 2514
rect 37617 2468 37687 2514
rect 37733 2468 37803 2514
rect 37849 2468 37919 2514
rect 37965 2468 38035 2514
rect 38081 2468 38151 2514
rect 38197 2468 38267 2514
rect 38313 2468 38383 2514
rect 38429 2468 38499 2514
rect 38545 2468 38615 2514
rect 38661 2468 38731 2514
rect 38777 2468 38847 2514
rect 38893 2468 38963 2514
rect 39009 2468 39079 2514
rect 39125 2468 39195 2514
rect 39241 2468 39311 2514
rect 39357 2468 39427 2514
rect 39473 2468 39543 2514
rect 39589 2468 39659 2514
rect 39705 2468 39775 2514
rect 39821 2468 39891 2514
rect 39937 2468 40007 2514
rect 40053 2468 40123 2514
rect 40169 2468 40180 2514
rect 28628 2398 40180 2468
rect 28628 2352 28639 2398
rect 28685 2352 28755 2398
rect 28801 2352 28871 2398
rect 28917 2352 28987 2398
rect 29033 2352 29103 2398
rect 29149 2352 29219 2398
rect 29265 2352 29335 2398
rect 29381 2352 29451 2398
rect 29497 2352 29567 2398
rect 29613 2352 29683 2398
rect 29729 2352 29799 2398
rect 29845 2352 29915 2398
rect 29961 2352 30031 2398
rect 30077 2352 30147 2398
rect 30193 2352 30263 2398
rect 30309 2352 30379 2398
rect 30425 2352 30495 2398
rect 30541 2352 30611 2398
rect 30657 2352 30727 2398
rect 30773 2352 30843 2398
rect 30889 2352 30959 2398
rect 31005 2352 31075 2398
rect 31121 2352 31191 2398
rect 31237 2352 31307 2398
rect 31353 2352 31423 2398
rect 31469 2352 31539 2398
rect 31585 2352 31655 2398
rect 31701 2352 31771 2398
rect 31817 2352 31887 2398
rect 31933 2352 32003 2398
rect 32049 2352 32119 2398
rect 32165 2352 32235 2398
rect 32281 2352 32351 2398
rect 32397 2352 32467 2398
rect 32513 2352 32583 2398
rect 32629 2352 32699 2398
rect 32745 2352 32815 2398
rect 32861 2352 32931 2398
rect 32977 2352 33047 2398
rect 33093 2352 33163 2398
rect 33209 2352 33279 2398
rect 33325 2352 33395 2398
rect 33441 2352 33511 2398
rect 33557 2352 33627 2398
rect 33673 2352 33743 2398
rect 33789 2352 33859 2398
rect 33905 2352 33975 2398
rect 34021 2352 34091 2398
rect 34137 2352 34207 2398
rect 34253 2352 34323 2398
rect 34369 2352 34439 2398
rect 34485 2352 34555 2398
rect 34601 2352 34671 2398
rect 34717 2352 34787 2398
rect 34833 2352 34903 2398
rect 34949 2352 35019 2398
rect 35065 2352 35135 2398
rect 35181 2352 35251 2398
rect 35297 2352 35367 2398
rect 35413 2352 35483 2398
rect 35529 2352 35599 2398
rect 35645 2352 35715 2398
rect 35761 2352 35831 2398
rect 35877 2352 35947 2398
rect 35993 2352 36063 2398
rect 36109 2352 36179 2398
rect 36225 2352 36295 2398
rect 36341 2352 36411 2398
rect 36457 2352 36527 2398
rect 36573 2352 36643 2398
rect 36689 2352 36759 2398
rect 36805 2352 36875 2398
rect 36921 2352 36991 2398
rect 37037 2352 37107 2398
rect 37153 2352 37223 2398
rect 37269 2352 37339 2398
rect 37385 2352 37455 2398
rect 37501 2352 37571 2398
rect 37617 2352 37687 2398
rect 37733 2352 37803 2398
rect 37849 2352 37919 2398
rect 37965 2352 38035 2398
rect 38081 2352 38151 2398
rect 38197 2352 38267 2398
rect 38313 2352 38383 2398
rect 38429 2352 38499 2398
rect 38545 2352 38615 2398
rect 38661 2352 38731 2398
rect 38777 2352 38847 2398
rect 38893 2352 38963 2398
rect 39009 2352 39079 2398
rect 39125 2352 39195 2398
rect 39241 2352 39311 2398
rect 39357 2352 39427 2398
rect 39473 2352 39543 2398
rect 39589 2352 39659 2398
rect 39705 2352 39775 2398
rect 39821 2352 39891 2398
rect 39937 2352 40007 2398
rect 40053 2352 40123 2398
rect 40169 2352 40180 2398
rect 28628 2282 40180 2352
rect 28628 2236 28639 2282
rect 28685 2236 28755 2282
rect 28801 2236 28871 2282
rect 28917 2236 28987 2282
rect 29033 2236 29103 2282
rect 29149 2236 29219 2282
rect 29265 2236 29335 2282
rect 29381 2236 29451 2282
rect 29497 2236 29567 2282
rect 29613 2236 29683 2282
rect 29729 2236 29799 2282
rect 29845 2236 29915 2282
rect 29961 2236 30031 2282
rect 30077 2236 30147 2282
rect 30193 2236 30263 2282
rect 30309 2236 30379 2282
rect 30425 2236 30495 2282
rect 30541 2236 30611 2282
rect 30657 2236 30727 2282
rect 30773 2236 30843 2282
rect 30889 2236 30959 2282
rect 31005 2236 31075 2282
rect 31121 2236 31191 2282
rect 31237 2236 31307 2282
rect 31353 2236 31423 2282
rect 31469 2236 31539 2282
rect 31585 2236 31655 2282
rect 31701 2236 31771 2282
rect 31817 2236 31887 2282
rect 31933 2236 32003 2282
rect 32049 2236 32119 2282
rect 32165 2236 32235 2282
rect 32281 2236 32351 2282
rect 32397 2236 32467 2282
rect 32513 2236 32583 2282
rect 32629 2236 32699 2282
rect 32745 2236 32815 2282
rect 32861 2236 32931 2282
rect 32977 2236 33047 2282
rect 33093 2236 33163 2282
rect 33209 2236 33279 2282
rect 33325 2236 33395 2282
rect 33441 2236 33511 2282
rect 33557 2236 33627 2282
rect 33673 2236 33743 2282
rect 33789 2236 33859 2282
rect 33905 2236 33975 2282
rect 34021 2236 34091 2282
rect 34137 2236 34207 2282
rect 34253 2236 34323 2282
rect 34369 2236 34439 2282
rect 34485 2236 34555 2282
rect 34601 2236 34671 2282
rect 34717 2236 34787 2282
rect 34833 2236 34903 2282
rect 34949 2236 35019 2282
rect 35065 2236 35135 2282
rect 35181 2236 35251 2282
rect 35297 2236 35367 2282
rect 35413 2236 35483 2282
rect 35529 2236 35599 2282
rect 35645 2236 35715 2282
rect 35761 2236 35831 2282
rect 35877 2236 35947 2282
rect 35993 2236 36063 2282
rect 36109 2236 36179 2282
rect 36225 2236 36295 2282
rect 36341 2236 36411 2282
rect 36457 2236 36527 2282
rect 36573 2236 36643 2282
rect 36689 2236 36759 2282
rect 36805 2236 36875 2282
rect 36921 2236 36991 2282
rect 37037 2236 37107 2282
rect 37153 2236 37223 2282
rect 37269 2236 37339 2282
rect 37385 2236 37455 2282
rect 37501 2236 37571 2282
rect 37617 2236 37687 2282
rect 37733 2236 37803 2282
rect 37849 2236 37919 2282
rect 37965 2236 38035 2282
rect 38081 2236 38151 2282
rect 38197 2236 38267 2282
rect 38313 2236 38383 2282
rect 38429 2236 38499 2282
rect 38545 2236 38615 2282
rect 38661 2236 38731 2282
rect 38777 2236 38847 2282
rect 38893 2236 38963 2282
rect 39009 2236 39079 2282
rect 39125 2236 39195 2282
rect 39241 2236 39311 2282
rect 39357 2236 39427 2282
rect 39473 2236 39543 2282
rect 39589 2236 39659 2282
rect 39705 2236 39775 2282
rect 39821 2236 39891 2282
rect 39937 2236 40007 2282
rect 40053 2236 40123 2282
rect 40169 2236 40180 2282
rect 28628 2166 40180 2236
rect 28628 2120 28639 2166
rect 28685 2120 28755 2166
rect 28801 2120 28871 2166
rect 28917 2120 28987 2166
rect 29033 2120 29103 2166
rect 29149 2120 29219 2166
rect 29265 2120 29335 2166
rect 29381 2120 29451 2166
rect 29497 2120 29567 2166
rect 29613 2120 29683 2166
rect 29729 2120 29799 2166
rect 29845 2120 29915 2166
rect 29961 2120 30031 2166
rect 30077 2120 30147 2166
rect 30193 2120 30263 2166
rect 30309 2120 30379 2166
rect 30425 2120 30495 2166
rect 30541 2120 30611 2166
rect 30657 2120 30727 2166
rect 30773 2120 30843 2166
rect 30889 2120 30959 2166
rect 31005 2120 31075 2166
rect 31121 2120 31191 2166
rect 31237 2120 31307 2166
rect 31353 2120 31423 2166
rect 31469 2120 31539 2166
rect 31585 2120 31655 2166
rect 31701 2120 31771 2166
rect 31817 2120 31887 2166
rect 31933 2120 32003 2166
rect 32049 2120 32119 2166
rect 32165 2120 32235 2166
rect 32281 2120 32351 2166
rect 32397 2120 32467 2166
rect 32513 2120 32583 2166
rect 32629 2120 32699 2166
rect 32745 2120 32815 2166
rect 32861 2120 32931 2166
rect 32977 2120 33047 2166
rect 33093 2120 33163 2166
rect 33209 2120 33279 2166
rect 33325 2120 33395 2166
rect 33441 2120 33511 2166
rect 33557 2120 33627 2166
rect 33673 2120 33743 2166
rect 33789 2120 33859 2166
rect 33905 2120 33975 2166
rect 34021 2120 34091 2166
rect 34137 2120 34207 2166
rect 34253 2120 34323 2166
rect 34369 2120 34439 2166
rect 34485 2120 34555 2166
rect 34601 2120 34671 2166
rect 34717 2120 34787 2166
rect 34833 2120 34903 2166
rect 34949 2120 35019 2166
rect 35065 2120 35135 2166
rect 35181 2120 35251 2166
rect 35297 2120 35367 2166
rect 35413 2120 35483 2166
rect 35529 2120 35599 2166
rect 35645 2120 35715 2166
rect 35761 2120 35831 2166
rect 35877 2120 35947 2166
rect 35993 2120 36063 2166
rect 36109 2120 36179 2166
rect 36225 2120 36295 2166
rect 36341 2120 36411 2166
rect 36457 2120 36527 2166
rect 36573 2120 36643 2166
rect 36689 2120 36759 2166
rect 36805 2120 36875 2166
rect 36921 2120 36991 2166
rect 37037 2120 37107 2166
rect 37153 2120 37223 2166
rect 37269 2120 37339 2166
rect 37385 2120 37455 2166
rect 37501 2120 37571 2166
rect 37617 2120 37687 2166
rect 37733 2120 37803 2166
rect 37849 2120 37919 2166
rect 37965 2120 38035 2166
rect 38081 2120 38151 2166
rect 38197 2120 38267 2166
rect 38313 2120 38383 2166
rect 38429 2120 38499 2166
rect 38545 2120 38615 2166
rect 38661 2120 38731 2166
rect 38777 2120 38847 2166
rect 38893 2120 38963 2166
rect 39009 2120 39079 2166
rect 39125 2120 39195 2166
rect 39241 2120 39311 2166
rect 39357 2120 39427 2166
rect 39473 2120 39543 2166
rect 39589 2120 39659 2166
rect 39705 2120 39775 2166
rect 39821 2120 39891 2166
rect 39937 2120 40007 2166
rect 40053 2120 40123 2166
rect 40169 2120 40180 2166
rect 28628 2050 40180 2120
rect 28628 2004 28639 2050
rect 28685 2004 28755 2050
rect 28801 2004 28871 2050
rect 28917 2004 28987 2050
rect 29033 2004 29103 2050
rect 29149 2004 29219 2050
rect 29265 2004 29335 2050
rect 29381 2004 29451 2050
rect 29497 2004 29567 2050
rect 29613 2004 29683 2050
rect 29729 2004 29799 2050
rect 29845 2004 29915 2050
rect 29961 2004 30031 2050
rect 30077 2004 30147 2050
rect 30193 2004 30263 2050
rect 30309 2004 30379 2050
rect 30425 2004 30495 2050
rect 30541 2004 30611 2050
rect 30657 2004 30727 2050
rect 30773 2004 30843 2050
rect 30889 2004 30959 2050
rect 31005 2004 31075 2050
rect 31121 2004 31191 2050
rect 31237 2004 31307 2050
rect 31353 2004 31423 2050
rect 31469 2004 31539 2050
rect 31585 2004 31655 2050
rect 31701 2004 31771 2050
rect 31817 2004 31887 2050
rect 31933 2004 32003 2050
rect 32049 2004 32119 2050
rect 32165 2004 32235 2050
rect 32281 2004 32351 2050
rect 32397 2004 32467 2050
rect 32513 2004 32583 2050
rect 32629 2004 32699 2050
rect 32745 2004 32815 2050
rect 32861 2004 32931 2050
rect 32977 2004 33047 2050
rect 33093 2004 33163 2050
rect 33209 2004 33279 2050
rect 33325 2004 33395 2050
rect 33441 2004 33511 2050
rect 33557 2004 33627 2050
rect 33673 2004 33743 2050
rect 33789 2004 33859 2050
rect 33905 2004 33975 2050
rect 34021 2004 34091 2050
rect 34137 2004 34207 2050
rect 34253 2004 34323 2050
rect 34369 2004 34439 2050
rect 34485 2004 34555 2050
rect 34601 2004 34671 2050
rect 34717 2004 34787 2050
rect 34833 2004 34903 2050
rect 34949 2004 35019 2050
rect 35065 2004 35135 2050
rect 35181 2004 35251 2050
rect 35297 2004 35367 2050
rect 35413 2004 35483 2050
rect 35529 2004 35599 2050
rect 35645 2004 35715 2050
rect 35761 2004 35831 2050
rect 35877 2004 35947 2050
rect 35993 2004 36063 2050
rect 36109 2004 36179 2050
rect 36225 2004 36295 2050
rect 36341 2004 36411 2050
rect 36457 2004 36527 2050
rect 36573 2004 36643 2050
rect 36689 2004 36759 2050
rect 36805 2004 36875 2050
rect 36921 2004 36991 2050
rect 37037 2004 37107 2050
rect 37153 2004 37223 2050
rect 37269 2004 37339 2050
rect 37385 2004 37455 2050
rect 37501 2004 37571 2050
rect 37617 2004 37687 2050
rect 37733 2004 37803 2050
rect 37849 2004 37919 2050
rect 37965 2004 38035 2050
rect 38081 2004 38151 2050
rect 38197 2004 38267 2050
rect 38313 2004 38383 2050
rect 38429 2004 38499 2050
rect 38545 2004 38615 2050
rect 38661 2004 38731 2050
rect 38777 2004 38847 2050
rect 38893 2004 38963 2050
rect 39009 2004 39079 2050
rect 39125 2004 39195 2050
rect 39241 2004 39311 2050
rect 39357 2004 39427 2050
rect 39473 2004 39543 2050
rect 39589 2004 39659 2050
rect 39705 2004 39775 2050
rect 39821 2004 39891 2050
rect 39937 2004 40007 2050
rect 40053 2004 40123 2050
rect 40169 2004 40180 2050
rect 28628 1934 40180 2004
rect 28628 1925 28639 1934
rect 27387 1888 28639 1925
rect 28685 1888 28755 1934
rect 28801 1888 28871 1934
rect 28917 1888 28987 1934
rect 29033 1888 29103 1934
rect 29149 1888 29219 1934
rect 29265 1888 29335 1934
rect 29381 1888 29451 1934
rect 29497 1888 29567 1934
rect 29613 1888 29683 1934
rect 29729 1888 29799 1934
rect 29845 1888 29915 1934
rect 29961 1888 30031 1934
rect 30077 1888 30147 1934
rect 30193 1888 30263 1934
rect 30309 1888 30379 1934
rect 30425 1888 30495 1934
rect 30541 1888 30611 1934
rect 30657 1888 30727 1934
rect 30773 1888 30843 1934
rect 30889 1888 30959 1934
rect 31005 1888 31075 1934
rect 31121 1888 31191 1934
rect 31237 1888 31307 1934
rect 31353 1888 31423 1934
rect 31469 1888 31539 1934
rect 31585 1888 31655 1934
rect 31701 1888 31771 1934
rect 31817 1888 31887 1934
rect 31933 1888 32003 1934
rect 32049 1888 32119 1934
rect 32165 1888 32235 1934
rect 32281 1888 32351 1934
rect 32397 1888 32467 1934
rect 32513 1888 32583 1934
rect 32629 1888 32699 1934
rect 32745 1888 32815 1934
rect 32861 1888 32931 1934
rect 32977 1888 33047 1934
rect 33093 1888 33163 1934
rect 33209 1888 33279 1934
rect 33325 1888 33395 1934
rect 33441 1888 33511 1934
rect 33557 1888 33627 1934
rect 33673 1888 33743 1934
rect 33789 1888 33859 1934
rect 33905 1888 33975 1934
rect 34021 1888 34091 1934
rect 34137 1888 34207 1934
rect 34253 1888 34323 1934
rect 34369 1888 34439 1934
rect 34485 1888 34555 1934
rect 34601 1888 34671 1934
rect 34717 1888 34787 1934
rect 34833 1888 34903 1934
rect 34949 1888 35019 1934
rect 35065 1888 35135 1934
rect 35181 1888 35251 1934
rect 35297 1888 35367 1934
rect 35413 1888 35483 1934
rect 35529 1888 35599 1934
rect 35645 1888 35715 1934
rect 35761 1888 35831 1934
rect 35877 1888 35947 1934
rect 35993 1888 36063 1934
rect 36109 1888 36179 1934
rect 36225 1888 36295 1934
rect 36341 1888 36411 1934
rect 36457 1888 36527 1934
rect 36573 1888 36643 1934
rect 36689 1888 36759 1934
rect 36805 1888 36875 1934
rect 36921 1888 36991 1934
rect 37037 1888 37107 1934
rect 37153 1888 37223 1934
rect 37269 1888 37339 1934
rect 37385 1888 37455 1934
rect 37501 1888 37571 1934
rect 37617 1888 37687 1934
rect 37733 1888 37803 1934
rect 37849 1888 37919 1934
rect 37965 1888 38035 1934
rect 38081 1888 38151 1934
rect 38197 1888 38267 1934
rect 38313 1888 38383 1934
rect 38429 1888 38499 1934
rect 38545 1888 38615 1934
rect 38661 1888 38731 1934
rect 38777 1888 38847 1934
rect 38893 1888 38963 1934
rect 39009 1888 39079 1934
rect 39125 1888 39195 1934
rect 39241 1888 39311 1934
rect 39357 1888 39427 1934
rect 39473 1888 39543 1934
rect 39589 1888 39659 1934
rect 39705 1888 39775 1934
rect 39821 1888 39891 1934
rect 39937 1888 40007 1934
rect 40053 1888 40123 1934
rect 40169 1925 40180 1934
rect 50834 3210 56586 3280
rect 50834 3164 50845 3210
rect 50891 3164 50961 3210
rect 51007 3164 51077 3210
rect 51123 3164 51193 3210
rect 51239 3164 51309 3210
rect 51355 3164 51425 3210
rect 51471 3164 51541 3210
rect 51587 3164 51657 3210
rect 51703 3164 51773 3210
rect 51819 3164 51889 3210
rect 51935 3164 52005 3210
rect 52051 3164 52121 3210
rect 52167 3164 52237 3210
rect 52283 3164 52353 3210
rect 52399 3164 52469 3210
rect 52515 3164 52585 3210
rect 52631 3164 52701 3210
rect 52747 3164 52817 3210
rect 52863 3164 52933 3210
rect 52979 3164 53049 3210
rect 53095 3164 53165 3210
rect 53211 3164 53281 3210
rect 53327 3164 53397 3210
rect 53443 3164 53513 3210
rect 53559 3164 53629 3210
rect 53675 3164 53745 3210
rect 53791 3164 53861 3210
rect 53907 3164 53977 3210
rect 54023 3164 54093 3210
rect 54139 3164 54209 3210
rect 54255 3164 54325 3210
rect 54371 3164 54441 3210
rect 54487 3164 54557 3210
rect 54603 3164 54673 3210
rect 54719 3164 54789 3210
rect 54835 3164 54905 3210
rect 54951 3164 55021 3210
rect 55067 3164 55137 3210
rect 55183 3164 55253 3210
rect 55299 3164 55369 3210
rect 55415 3164 55485 3210
rect 55531 3164 55601 3210
rect 55647 3164 55717 3210
rect 55763 3164 55833 3210
rect 55879 3164 55949 3210
rect 55995 3164 56065 3210
rect 56111 3164 56181 3210
rect 56227 3164 56297 3210
rect 56343 3164 56413 3210
rect 56459 3164 56529 3210
rect 56575 3164 56586 3210
rect 50834 3094 56586 3164
rect 50834 3048 50845 3094
rect 50891 3048 50961 3094
rect 51007 3048 51077 3094
rect 51123 3048 51193 3094
rect 51239 3048 51309 3094
rect 51355 3048 51425 3094
rect 51471 3048 51541 3094
rect 51587 3048 51657 3094
rect 51703 3048 51773 3094
rect 51819 3048 51889 3094
rect 51935 3048 52005 3094
rect 52051 3048 52121 3094
rect 52167 3048 52237 3094
rect 52283 3048 52353 3094
rect 52399 3048 52469 3094
rect 52515 3048 52585 3094
rect 52631 3048 52701 3094
rect 52747 3048 52817 3094
rect 52863 3048 52933 3094
rect 52979 3048 53049 3094
rect 53095 3048 53165 3094
rect 53211 3048 53281 3094
rect 53327 3048 53397 3094
rect 53443 3048 53513 3094
rect 53559 3048 53629 3094
rect 53675 3048 53745 3094
rect 53791 3048 53861 3094
rect 53907 3048 53977 3094
rect 54023 3048 54093 3094
rect 54139 3048 54209 3094
rect 54255 3048 54325 3094
rect 54371 3048 54441 3094
rect 54487 3048 54557 3094
rect 54603 3048 54673 3094
rect 54719 3048 54789 3094
rect 54835 3048 54905 3094
rect 54951 3048 55021 3094
rect 55067 3048 55137 3094
rect 55183 3048 55253 3094
rect 55299 3048 55369 3094
rect 55415 3048 55485 3094
rect 55531 3048 55601 3094
rect 55647 3048 55717 3094
rect 55763 3048 55833 3094
rect 55879 3048 55949 3094
rect 55995 3048 56065 3094
rect 56111 3048 56181 3094
rect 56227 3048 56297 3094
rect 56343 3048 56413 3094
rect 56459 3048 56529 3094
rect 56575 3048 56586 3094
rect 50834 2978 56586 3048
rect 50834 2932 50845 2978
rect 50891 2932 50961 2978
rect 51007 2932 51077 2978
rect 51123 2932 51193 2978
rect 51239 2932 51309 2978
rect 51355 2932 51425 2978
rect 51471 2932 51541 2978
rect 51587 2932 51657 2978
rect 51703 2932 51773 2978
rect 51819 2932 51889 2978
rect 51935 2932 52005 2978
rect 52051 2932 52121 2978
rect 52167 2932 52237 2978
rect 52283 2932 52353 2978
rect 52399 2932 52469 2978
rect 52515 2932 52585 2978
rect 52631 2932 52701 2978
rect 52747 2932 52817 2978
rect 52863 2932 52933 2978
rect 52979 2932 53049 2978
rect 53095 2932 53165 2978
rect 53211 2932 53281 2978
rect 53327 2932 53397 2978
rect 53443 2932 53513 2978
rect 53559 2932 53629 2978
rect 53675 2932 53745 2978
rect 53791 2932 53861 2978
rect 53907 2932 53977 2978
rect 54023 2932 54093 2978
rect 54139 2932 54209 2978
rect 54255 2932 54325 2978
rect 54371 2932 54441 2978
rect 54487 2932 54557 2978
rect 54603 2932 54673 2978
rect 54719 2932 54789 2978
rect 54835 2932 54905 2978
rect 54951 2932 55021 2978
rect 55067 2932 55137 2978
rect 55183 2932 55253 2978
rect 55299 2932 55369 2978
rect 55415 2932 55485 2978
rect 55531 2932 55601 2978
rect 55647 2932 55717 2978
rect 55763 2932 55833 2978
rect 55879 2932 55949 2978
rect 55995 2932 56065 2978
rect 56111 2932 56181 2978
rect 56227 2932 56297 2978
rect 56343 2932 56413 2978
rect 56459 2932 56529 2978
rect 56575 2932 56586 2978
rect 50834 2862 56586 2932
rect 50834 2816 50845 2862
rect 50891 2816 50961 2862
rect 51007 2816 51077 2862
rect 51123 2816 51193 2862
rect 51239 2816 51309 2862
rect 51355 2816 51425 2862
rect 51471 2816 51541 2862
rect 51587 2816 51657 2862
rect 51703 2816 51773 2862
rect 51819 2816 51889 2862
rect 51935 2816 52005 2862
rect 52051 2816 52121 2862
rect 52167 2816 52237 2862
rect 52283 2816 52353 2862
rect 52399 2816 52469 2862
rect 52515 2816 52585 2862
rect 52631 2816 52701 2862
rect 52747 2816 52817 2862
rect 52863 2816 52933 2862
rect 52979 2816 53049 2862
rect 53095 2816 53165 2862
rect 53211 2816 53281 2862
rect 53327 2816 53397 2862
rect 53443 2816 53513 2862
rect 53559 2816 53629 2862
rect 53675 2816 53745 2862
rect 53791 2816 53861 2862
rect 53907 2816 53977 2862
rect 54023 2816 54093 2862
rect 54139 2816 54209 2862
rect 54255 2816 54325 2862
rect 54371 2816 54441 2862
rect 54487 2816 54557 2862
rect 54603 2816 54673 2862
rect 54719 2816 54789 2862
rect 54835 2816 54905 2862
rect 54951 2816 55021 2862
rect 55067 2816 55137 2862
rect 55183 2816 55253 2862
rect 55299 2816 55369 2862
rect 55415 2816 55485 2862
rect 55531 2816 55601 2862
rect 55647 2816 55717 2862
rect 55763 2816 55833 2862
rect 55879 2816 55949 2862
rect 55995 2816 56065 2862
rect 56111 2816 56181 2862
rect 56227 2816 56297 2862
rect 56343 2816 56413 2862
rect 56459 2816 56529 2862
rect 56575 2816 56586 2862
rect 50834 2746 56586 2816
rect 50834 2700 50845 2746
rect 50891 2700 50961 2746
rect 51007 2700 51077 2746
rect 51123 2700 51193 2746
rect 51239 2700 51309 2746
rect 51355 2700 51425 2746
rect 51471 2700 51541 2746
rect 51587 2700 51657 2746
rect 51703 2700 51773 2746
rect 51819 2700 51889 2746
rect 51935 2700 52005 2746
rect 52051 2700 52121 2746
rect 52167 2700 52237 2746
rect 52283 2700 52353 2746
rect 52399 2700 52469 2746
rect 52515 2700 52585 2746
rect 52631 2700 52701 2746
rect 52747 2700 52817 2746
rect 52863 2700 52933 2746
rect 52979 2700 53049 2746
rect 53095 2700 53165 2746
rect 53211 2700 53281 2746
rect 53327 2700 53397 2746
rect 53443 2700 53513 2746
rect 53559 2700 53629 2746
rect 53675 2700 53745 2746
rect 53791 2700 53861 2746
rect 53907 2700 53977 2746
rect 54023 2700 54093 2746
rect 54139 2700 54209 2746
rect 54255 2700 54325 2746
rect 54371 2700 54441 2746
rect 54487 2700 54557 2746
rect 54603 2700 54673 2746
rect 54719 2700 54789 2746
rect 54835 2700 54905 2746
rect 54951 2700 55021 2746
rect 55067 2700 55137 2746
rect 55183 2700 55253 2746
rect 55299 2700 55369 2746
rect 55415 2700 55485 2746
rect 55531 2700 55601 2746
rect 55647 2700 55717 2746
rect 55763 2700 55833 2746
rect 55879 2700 55949 2746
rect 55995 2700 56065 2746
rect 56111 2700 56181 2746
rect 56227 2700 56297 2746
rect 56343 2700 56413 2746
rect 56459 2700 56529 2746
rect 56575 2700 56586 2746
rect 50834 2630 56586 2700
rect 50834 2584 50845 2630
rect 50891 2584 50961 2630
rect 51007 2584 51077 2630
rect 51123 2584 51193 2630
rect 51239 2584 51309 2630
rect 51355 2584 51425 2630
rect 51471 2584 51541 2630
rect 51587 2584 51657 2630
rect 51703 2584 51773 2630
rect 51819 2584 51889 2630
rect 51935 2584 52005 2630
rect 52051 2584 52121 2630
rect 52167 2584 52237 2630
rect 52283 2584 52353 2630
rect 52399 2584 52469 2630
rect 52515 2584 52585 2630
rect 52631 2584 52701 2630
rect 52747 2584 52817 2630
rect 52863 2584 52933 2630
rect 52979 2584 53049 2630
rect 53095 2584 53165 2630
rect 53211 2584 53281 2630
rect 53327 2584 53397 2630
rect 53443 2584 53513 2630
rect 53559 2584 53629 2630
rect 53675 2584 53745 2630
rect 53791 2584 53861 2630
rect 53907 2584 53977 2630
rect 54023 2584 54093 2630
rect 54139 2584 54209 2630
rect 54255 2584 54325 2630
rect 54371 2584 54441 2630
rect 54487 2584 54557 2630
rect 54603 2584 54673 2630
rect 54719 2584 54789 2630
rect 54835 2584 54905 2630
rect 54951 2584 55021 2630
rect 55067 2584 55137 2630
rect 55183 2584 55253 2630
rect 55299 2584 55369 2630
rect 55415 2584 55485 2630
rect 55531 2584 55601 2630
rect 55647 2584 55717 2630
rect 55763 2584 55833 2630
rect 55879 2584 55949 2630
rect 55995 2584 56065 2630
rect 56111 2584 56181 2630
rect 56227 2584 56297 2630
rect 56343 2584 56413 2630
rect 56459 2584 56529 2630
rect 56575 2584 56586 2630
rect 50834 2514 56586 2584
rect 50834 2468 50845 2514
rect 50891 2468 50961 2514
rect 51007 2468 51077 2514
rect 51123 2468 51193 2514
rect 51239 2468 51309 2514
rect 51355 2468 51425 2514
rect 51471 2468 51541 2514
rect 51587 2468 51657 2514
rect 51703 2468 51773 2514
rect 51819 2468 51889 2514
rect 51935 2468 52005 2514
rect 52051 2468 52121 2514
rect 52167 2468 52237 2514
rect 52283 2468 52353 2514
rect 52399 2468 52469 2514
rect 52515 2468 52585 2514
rect 52631 2468 52701 2514
rect 52747 2468 52817 2514
rect 52863 2468 52933 2514
rect 52979 2468 53049 2514
rect 53095 2468 53165 2514
rect 53211 2468 53281 2514
rect 53327 2468 53397 2514
rect 53443 2468 53513 2514
rect 53559 2468 53629 2514
rect 53675 2468 53745 2514
rect 53791 2468 53861 2514
rect 53907 2468 53977 2514
rect 54023 2468 54093 2514
rect 54139 2468 54209 2514
rect 54255 2468 54325 2514
rect 54371 2468 54441 2514
rect 54487 2468 54557 2514
rect 54603 2468 54673 2514
rect 54719 2468 54789 2514
rect 54835 2468 54905 2514
rect 54951 2468 55021 2514
rect 55067 2468 55137 2514
rect 55183 2468 55253 2514
rect 55299 2468 55369 2514
rect 55415 2468 55485 2514
rect 55531 2468 55601 2514
rect 55647 2468 55717 2514
rect 55763 2468 55833 2514
rect 55879 2468 55949 2514
rect 55995 2468 56065 2514
rect 56111 2468 56181 2514
rect 56227 2468 56297 2514
rect 56343 2468 56413 2514
rect 56459 2468 56529 2514
rect 56575 2468 56586 2514
rect 50834 2398 56586 2468
rect 50834 2352 50845 2398
rect 50891 2352 50961 2398
rect 51007 2352 51077 2398
rect 51123 2352 51193 2398
rect 51239 2352 51309 2398
rect 51355 2352 51425 2398
rect 51471 2352 51541 2398
rect 51587 2352 51657 2398
rect 51703 2352 51773 2398
rect 51819 2352 51889 2398
rect 51935 2352 52005 2398
rect 52051 2352 52121 2398
rect 52167 2352 52237 2398
rect 52283 2352 52353 2398
rect 52399 2352 52469 2398
rect 52515 2352 52585 2398
rect 52631 2352 52701 2398
rect 52747 2352 52817 2398
rect 52863 2352 52933 2398
rect 52979 2352 53049 2398
rect 53095 2352 53165 2398
rect 53211 2352 53281 2398
rect 53327 2352 53397 2398
rect 53443 2352 53513 2398
rect 53559 2352 53629 2398
rect 53675 2352 53745 2398
rect 53791 2352 53861 2398
rect 53907 2352 53977 2398
rect 54023 2352 54093 2398
rect 54139 2352 54209 2398
rect 54255 2352 54325 2398
rect 54371 2352 54441 2398
rect 54487 2352 54557 2398
rect 54603 2352 54673 2398
rect 54719 2352 54789 2398
rect 54835 2352 54905 2398
rect 54951 2352 55021 2398
rect 55067 2352 55137 2398
rect 55183 2352 55253 2398
rect 55299 2352 55369 2398
rect 55415 2352 55485 2398
rect 55531 2352 55601 2398
rect 55647 2352 55717 2398
rect 55763 2352 55833 2398
rect 55879 2352 55949 2398
rect 55995 2352 56065 2398
rect 56111 2352 56181 2398
rect 56227 2352 56297 2398
rect 56343 2352 56413 2398
rect 56459 2352 56529 2398
rect 56575 2352 56586 2398
rect 50834 2282 56586 2352
rect 50834 2236 50845 2282
rect 50891 2236 50961 2282
rect 51007 2236 51077 2282
rect 51123 2236 51193 2282
rect 51239 2236 51309 2282
rect 51355 2236 51425 2282
rect 51471 2236 51541 2282
rect 51587 2236 51657 2282
rect 51703 2236 51773 2282
rect 51819 2236 51889 2282
rect 51935 2236 52005 2282
rect 52051 2236 52121 2282
rect 52167 2236 52237 2282
rect 52283 2236 52353 2282
rect 52399 2236 52469 2282
rect 52515 2236 52585 2282
rect 52631 2236 52701 2282
rect 52747 2236 52817 2282
rect 52863 2236 52933 2282
rect 52979 2236 53049 2282
rect 53095 2236 53165 2282
rect 53211 2236 53281 2282
rect 53327 2236 53397 2282
rect 53443 2236 53513 2282
rect 53559 2236 53629 2282
rect 53675 2236 53745 2282
rect 53791 2236 53861 2282
rect 53907 2236 53977 2282
rect 54023 2236 54093 2282
rect 54139 2236 54209 2282
rect 54255 2236 54325 2282
rect 54371 2236 54441 2282
rect 54487 2236 54557 2282
rect 54603 2236 54673 2282
rect 54719 2236 54789 2282
rect 54835 2236 54905 2282
rect 54951 2236 55021 2282
rect 55067 2236 55137 2282
rect 55183 2236 55253 2282
rect 55299 2236 55369 2282
rect 55415 2236 55485 2282
rect 55531 2236 55601 2282
rect 55647 2236 55717 2282
rect 55763 2236 55833 2282
rect 55879 2236 55949 2282
rect 55995 2236 56065 2282
rect 56111 2236 56181 2282
rect 56227 2236 56297 2282
rect 56343 2236 56413 2282
rect 56459 2236 56529 2282
rect 56575 2236 56586 2282
rect 50834 2166 56586 2236
rect 50834 2120 50845 2166
rect 50891 2120 50961 2166
rect 51007 2120 51077 2166
rect 51123 2120 51193 2166
rect 51239 2120 51309 2166
rect 51355 2120 51425 2166
rect 51471 2120 51541 2166
rect 51587 2120 51657 2166
rect 51703 2120 51773 2166
rect 51819 2120 51889 2166
rect 51935 2120 52005 2166
rect 52051 2120 52121 2166
rect 52167 2120 52237 2166
rect 52283 2120 52353 2166
rect 52399 2120 52469 2166
rect 52515 2120 52585 2166
rect 52631 2120 52701 2166
rect 52747 2120 52817 2166
rect 52863 2120 52933 2166
rect 52979 2120 53049 2166
rect 53095 2120 53165 2166
rect 53211 2120 53281 2166
rect 53327 2120 53397 2166
rect 53443 2120 53513 2166
rect 53559 2120 53629 2166
rect 53675 2120 53745 2166
rect 53791 2120 53861 2166
rect 53907 2120 53977 2166
rect 54023 2120 54093 2166
rect 54139 2120 54209 2166
rect 54255 2120 54325 2166
rect 54371 2120 54441 2166
rect 54487 2120 54557 2166
rect 54603 2120 54673 2166
rect 54719 2120 54789 2166
rect 54835 2120 54905 2166
rect 54951 2120 55021 2166
rect 55067 2120 55137 2166
rect 55183 2120 55253 2166
rect 55299 2120 55369 2166
rect 55415 2120 55485 2166
rect 55531 2120 55601 2166
rect 55647 2120 55717 2166
rect 55763 2120 55833 2166
rect 55879 2120 55949 2166
rect 55995 2120 56065 2166
rect 56111 2120 56181 2166
rect 56227 2120 56297 2166
rect 56343 2120 56413 2166
rect 56459 2120 56529 2166
rect 56575 2120 56586 2166
rect 50834 2050 56586 2120
rect 50834 2004 50845 2050
rect 50891 2004 50961 2050
rect 51007 2004 51077 2050
rect 51123 2004 51193 2050
rect 51239 2004 51309 2050
rect 51355 2004 51425 2050
rect 51471 2004 51541 2050
rect 51587 2004 51657 2050
rect 51703 2004 51773 2050
rect 51819 2004 51889 2050
rect 51935 2004 52005 2050
rect 52051 2004 52121 2050
rect 52167 2004 52237 2050
rect 52283 2004 52353 2050
rect 52399 2004 52469 2050
rect 52515 2004 52585 2050
rect 52631 2004 52701 2050
rect 52747 2004 52817 2050
rect 52863 2004 52933 2050
rect 52979 2004 53049 2050
rect 53095 2004 53165 2050
rect 53211 2004 53281 2050
rect 53327 2004 53397 2050
rect 53443 2004 53513 2050
rect 53559 2004 53629 2050
rect 53675 2004 53745 2050
rect 53791 2004 53861 2050
rect 53907 2004 53977 2050
rect 54023 2004 54093 2050
rect 54139 2004 54209 2050
rect 54255 2004 54325 2050
rect 54371 2004 54441 2050
rect 54487 2004 54557 2050
rect 54603 2004 54673 2050
rect 54719 2004 54789 2050
rect 54835 2004 54905 2050
rect 54951 2004 55021 2050
rect 55067 2004 55137 2050
rect 55183 2004 55253 2050
rect 55299 2004 55369 2050
rect 55415 2004 55485 2050
rect 55531 2004 55601 2050
rect 55647 2004 55717 2050
rect 55763 2004 55833 2050
rect 55879 2004 55949 2050
rect 55995 2004 56065 2050
rect 56111 2004 56181 2050
rect 56227 2004 56297 2050
rect 56343 2004 56413 2050
rect 56459 2004 56529 2050
rect 56575 2004 56586 2050
rect 50834 1934 56586 2004
rect 50834 1925 50845 1934
rect 40169 1888 50845 1925
rect 50891 1888 50961 1934
rect 51007 1888 51077 1934
rect 51123 1888 51193 1934
rect 51239 1888 51309 1934
rect 51355 1888 51425 1934
rect 51471 1888 51541 1934
rect 51587 1888 51657 1934
rect 51703 1888 51773 1934
rect 51819 1888 51889 1934
rect 51935 1888 52005 1934
rect 52051 1888 52121 1934
rect 52167 1888 52237 1934
rect 52283 1888 52353 1934
rect 52399 1888 52469 1934
rect 52515 1888 52585 1934
rect 52631 1888 52701 1934
rect 52747 1888 52817 1934
rect 52863 1888 52933 1934
rect 52979 1888 53049 1934
rect 53095 1888 53165 1934
rect 53211 1888 53281 1934
rect 53327 1888 53397 1934
rect 53443 1888 53513 1934
rect 53559 1888 53629 1934
rect 53675 1888 53745 1934
rect 53791 1888 53861 1934
rect 53907 1888 53977 1934
rect 54023 1888 54093 1934
rect 54139 1888 54209 1934
rect 54255 1888 54325 1934
rect 54371 1888 54441 1934
rect 54487 1888 54557 1934
rect 54603 1888 54673 1934
rect 54719 1888 54789 1934
rect 54835 1888 54905 1934
rect 54951 1888 55021 1934
rect 55067 1888 55137 1934
rect 55183 1888 55253 1934
rect 55299 1888 55369 1934
rect 55415 1888 55485 1934
rect 55531 1888 55601 1934
rect 55647 1888 55717 1934
rect 55763 1888 55833 1934
rect 55879 1888 55949 1934
rect 55995 1888 56065 1934
rect 56111 1888 56181 1934
rect 56227 1888 56297 1934
rect 56343 1888 56413 1934
rect 56459 1888 56529 1934
rect 56575 1925 56586 1934
rect 57295 3882 57383 3934
rect 57435 3882 57595 3934
rect 57647 3882 57736 3934
rect 57295 3717 57736 3882
rect 57295 3665 57383 3717
rect 57435 3665 57595 3717
rect 57647 3665 57736 3717
rect 57295 1925 57736 3665
rect 56575 1888 57736 1925
rect 27387 1818 57736 1888
rect 27387 1772 28639 1818
rect 28685 1772 28755 1818
rect 28801 1772 28871 1818
rect 28917 1772 28987 1818
rect 29033 1772 29103 1818
rect 29149 1772 29219 1818
rect 29265 1772 29335 1818
rect 29381 1772 29451 1818
rect 29497 1772 29567 1818
rect 29613 1772 29683 1818
rect 29729 1772 29799 1818
rect 29845 1772 29915 1818
rect 29961 1772 30031 1818
rect 30077 1772 30147 1818
rect 30193 1772 30263 1818
rect 30309 1772 30379 1818
rect 30425 1772 30495 1818
rect 30541 1772 30611 1818
rect 30657 1772 30727 1818
rect 30773 1772 30843 1818
rect 30889 1772 30959 1818
rect 31005 1772 31075 1818
rect 31121 1772 31191 1818
rect 31237 1772 31307 1818
rect 31353 1772 31423 1818
rect 31469 1772 31539 1818
rect 31585 1772 31655 1818
rect 31701 1772 31771 1818
rect 31817 1772 31887 1818
rect 31933 1772 32003 1818
rect 32049 1772 32119 1818
rect 32165 1772 32235 1818
rect 32281 1772 32351 1818
rect 32397 1772 32467 1818
rect 32513 1772 32583 1818
rect 32629 1772 32699 1818
rect 32745 1772 32815 1818
rect 32861 1772 32931 1818
rect 32977 1772 33047 1818
rect 33093 1772 33163 1818
rect 33209 1772 33279 1818
rect 33325 1772 33395 1818
rect 33441 1772 33511 1818
rect 33557 1772 33627 1818
rect 33673 1772 33743 1818
rect 33789 1772 33859 1818
rect 33905 1772 33975 1818
rect 34021 1772 34091 1818
rect 34137 1772 34207 1818
rect 34253 1772 34323 1818
rect 34369 1772 34439 1818
rect 34485 1772 34555 1818
rect 34601 1772 34671 1818
rect 34717 1772 34787 1818
rect 34833 1772 34903 1818
rect 34949 1772 35019 1818
rect 35065 1772 35135 1818
rect 35181 1772 35251 1818
rect 35297 1772 35367 1818
rect 35413 1772 35483 1818
rect 35529 1772 35599 1818
rect 35645 1772 35715 1818
rect 35761 1772 35831 1818
rect 35877 1772 35947 1818
rect 35993 1772 36063 1818
rect 36109 1772 36179 1818
rect 36225 1772 36295 1818
rect 36341 1772 36411 1818
rect 36457 1772 36527 1818
rect 36573 1772 36643 1818
rect 36689 1772 36759 1818
rect 36805 1772 36875 1818
rect 36921 1772 36991 1818
rect 37037 1772 37107 1818
rect 37153 1772 37223 1818
rect 37269 1772 37339 1818
rect 37385 1772 37455 1818
rect 37501 1772 37571 1818
rect 37617 1772 37687 1818
rect 37733 1772 37803 1818
rect 37849 1772 37919 1818
rect 37965 1772 38035 1818
rect 38081 1772 38151 1818
rect 38197 1772 38267 1818
rect 38313 1772 38383 1818
rect 38429 1772 38499 1818
rect 38545 1772 38615 1818
rect 38661 1772 38731 1818
rect 38777 1772 38847 1818
rect 38893 1772 38963 1818
rect 39009 1772 39079 1818
rect 39125 1772 39195 1818
rect 39241 1772 39311 1818
rect 39357 1772 39427 1818
rect 39473 1772 39543 1818
rect 39589 1772 39659 1818
rect 39705 1772 39775 1818
rect 39821 1772 39891 1818
rect 39937 1772 40007 1818
rect 40053 1772 40123 1818
rect 40169 1772 50845 1818
rect 50891 1772 50961 1818
rect 51007 1772 51077 1818
rect 51123 1772 51193 1818
rect 51239 1772 51309 1818
rect 51355 1772 51425 1818
rect 51471 1772 51541 1818
rect 51587 1772 51657 1818
rect 51703 1772 51773 1818
rect 51819 1772 51889 1818
rect 51935 1772 52005 1818
rect 52051 1772 52121 1818
rect 52167 1772 52237 1818
rect 52283 1772 52353 1818
rect 52399 1772 52469 1818
rect 52515 1772 52585 1818
rect 52631 1772 52701 1818
rect 52747 1772 52817 1818
rect 52863 1772 52933 1818
rect 52979 1772 53049 1818
rect 53095 1772 53165 1818
rect 53211 1772 53281 1818
rect 53327 1772 53397 1818
rect 53443 1772 53513 1818
rect 53559 1772 53629 1818
rect 53675 1772 53745 1818
rect 53791 1772 53861 1818
rect 53907 1772 53977 1818
rect 54023 1772 54093 1818
rect 54139 1772 54209 1818
rect 54255 1772 54325 1818
rect 54371 1772 54441 1818
rect 54487 1772 54557 1818
rect 54603 1772 54673 1818
rect 54719 1772 54789 1818
rect 54835 1772 54905 1818
rect 54951 1772 55021 1818
rect 55067 1772 55137 1818
rect 55183 1772 55253 1818
rect 55299 1772 55369 1818
rect 55415 1772 55485 1818
rect 55531 1772 55601 1818
rect 55647 1772 55717 1818
rect 55763 1772 55833 1818
rect 55879 1772 55949 1818
rect 55995 1772 56065 1818
rect 56111 1772 56181 1818
rect 56227 1772 56297 1818
rect 56343 1772 56413 1818
rect 56459 1772 56529 1818
rect 56575 1772 57736 1818
rect 57909 33432 58351 33519
rect 57909 33380 57998 33432
rect 58050 33380 58210 33432
rect 58262 33380 58351 33432
rect 57909 33215 58351 33380
rect 57909 33163 57998 33215
rect 58050 33163 58210 33215
rect 58262 33163 58351 33215
rect 57909 32997 58351 33163
rect 57909 32945 57998 32997
rect 58050 32945 58210 32997
rect 58262 32945 58351 32997
rect 57909 32779 58351 32945
rect 57909 32727 57998 32779
rect 58050 32727 58210 32779
rect 58262 32727 58351 32779
rect 57909 32562 58351 32727
rect 57909 32510 57998 32562
rect 58050 32510 58210 32562
rect 58262 32510 58351 32562
rect 57909 32344 58351 32510
rect 57909 32292 57998 32344
rect 58050 32292 58210 32344
rect 58262 32292 58351 32344
rect 57909 32127 58351 32292
rect 57909 32075 57998 32127
rect 58050 32075 58210 32127
rect 58262 32075 58351 32127
rect 57909 31909 58351 32075
rect 83398 32048 83834 32122
rect 57909 31857 57998 31909
rect 58050 31857 58210 31909
rect 58262 31857 58351 31909
rect 57909 31691 58351 31857
rect 57909 31639 57998 31691
rect 58050 31639 58210 31691
rect 58262 31639 58351 31691
rect 57909 31474 58351 31639
rect 57909 31422 57998 31474
rect 58050 31422 58210 31474
rect 58262 31422 58351 31474
rect 57909 31256 58351 31422
rect 57909 31204 57998 31256
rect 58050 31204 58210 31256
rect 58262 31204 58351 31256
rect 57909 31038 58351 31204
rect 57909 30986 57998 31038
rect 58050 30986 58210 31038
rect 58262 30986 58351 31038
rect 57909 30821 58351 30986
rect 57909 30769 57998 30821
rect 58050 30769 58210 30821
rect 58262 30769 58351 30821
rect 57909 30603 58351 30769
rect 57909 30551 57998 30603
rect 58050 30551 58210 30603
rect 58262 30551 58351 30603
rect 57909 30386 58351 30551
rect 57909 30334 57998 30386
rect 58050 30334 58210 30386
rect 58262 30334 58351 30386
rect 57909 30168 58351 30334
rect 57909 30116 57998 30168
rect 58050 30116 58210 30168
rect 58262 30116 58351 30168
rect 57909 29950 58351 30116
rect 57909 29898 57998 29950
rect 58050 29898 58210 29950
rect 58262 29898 58351 29950
rect 57909 29733 58351 29898
rect 57909 29681 57998 29733
rect 58050 29681 58210 29733
rect 58262 29681 58351 29733
rect 57909 29515 58351 29681
rect 57909 29463 57998 29515
rect 58050 29463 58210 29515
rect 58262 29463 58351 29515
rect 57909 29297 58351 29463
rect 57909 29245 57998 29297
rect 58050 29245 58210 29297
rect 58262 29245 58351 29297
rect 57909 29080 58351 29245
rect 57909 29028 57998 29080
rect 58050 29028 58210 29080
rect 58262 29028 58351 29080
rect 57909 28862 58351 29028
rect 57909 28810 57998 28862
rect 58050 28810 58210 28862
rect 58262 28810 58351 28862
rect 57909 28644 58351 28810
rect 57909 28592 57998 28644
rect 58050 28592 58210 28644
rect 58262 28592 58351 28644
rect 57909 28427 58351 28592
rect 57909 28375 57998 28427
rect 58050 28375 58210 28427
rect 58262 28375 58351 28427
rect 57909 28209 58351 28375
rect 57909 28157 57998 28209
rect 58050 28157 58210 28209
rect 58262 28157 58351 28209
rect 57909 27992 58351 28157
rect 57909 27940 57998 27992
rect 58050 27940 58210 27992
rect 58262 27940 58351 27992
rect 57909 27774 58351 27940
rect 57909 27722 57998 27774
rect 58050 27722 58210 27774
rect 58262 27722 58351 27774
rect 57909 27556 58351 27722
rect 57909 27504 57998 27556
rect 58050 27504 58210 27556
rect 58262 27504 58351 27556
rect 57909 27339 58351 27504
rect 57909 27287 57998 27339
rect 58050 27287 58210 27339
rect 58262 27287 58351 27339
rect 57909 27121 58351 27287
rect 57909 27069 57998 27121
rect 58050 27069 58210 27121
rect 58262 27069 58351 27121
rect 57909 26903 58351 27069
rect 57909 26851 57998 26903
rect 58050 26851 58210 26903
rect 58262 26851 58351 26903
rect 57909 26686 58351 26851
rect 57909 26634 57998 26686
rect 58050 26634 58210 26686
rect 58262 26634 58351 26686
rect 57909 26468 58351 26634
rect 57909 26416 57998 26468
rect 58050 26416 58210 26468
rect 58262 26416 58351 26468
rect 57909 26250 58351 26416
rect 57909 26198 57998 26250
rect 58050 26198 58210 26250
rect 58262 26198 58351 26250
rect 57909 26033 58351 26198
rect 57909 25981 57998 26033
rect 58050 25981 58210 26033
rect 58262 25981 58351 26033
rect 57909 25815 58351 25981
rect 57909 25763 57998 25815
rect 58050 25763 58210 25815
rect 58262 25763 58351 25815
rect 57909 25598 58351 25763
rect 57909 25546 57998 25598
rect 58050 25546 58210 25598
rect 58262 25546 58351 25598
rect 57909 25380 58351 25546
rect 57909 25328 57998 25380
rect 58050 25328 58210 25380
rect 58262 25328 58351 25380
rect 57909 25162 58351 25328
rect 57909 25110 57998 25162
rect 58050 25110 58210 25162
rect 58262 25110 58351 25162
rect 57909 24945 58351 25110
rect 57909 24893 57998 24945
rect 58050 24893 58210 24945
rect 58262 24893 58351 24945
rect 57909 24727 58351 24893
rect 57909 24675 57998 24727
rect 58050 24675 58210 24727
rect 58262 24675 58351 24727
rect 57909 24509 58351 24675
rect 57909 24457 57998 24509
rect 58050 24457 58210 24509
rect 58262 24457 58351 24509
rect 57909 24292 58351 24457
rect 57909 24240 57998 24292
rect 58050 24240 58210 24292
rect 58262 24240 58351 24292
rect 57909 24074 58351 24240
rect 57909 24022 57998 24074
rect 58050 24022 58210 24074
rect 58262 24022 58351 24074
rect 57909 23857 58351 24022
rect 57909 23805 57998 23857
rect 58050 23805 58210 23857
rect 58262 23805 58351 23857
rect 57909 23639 58351 23805
rect 57909 23587 57998 23639
rect 58050 23587 58210 23639
rect 58262 23587 58351 23639
rect 57909 23421 58351 23587
rect 57909 23369 57998 23421
rect 58050 23369 58210 23421
rect 58262 23369 58351 23421
rect 57909 23204 58351 23369
rect 57909 23152 57998 23204
rect 58050 23152 58210 23204
rect 58262 23152 58351 23204
rect 57909 22986 58351 23152
rect 57909 22934 57998 22986
rect 58050 22934 58210 22986
rect 58262 22934 58351 22986
rect 57909 22768 58351 22934
rect 57909 22716 57998 22768
rect 58050 22716 58210 22768
rect 58262 22716 58351 22768
rect 57909 22551 58351 22716
rect 57909 22499 57998 22551
rect 58050 22499 58210 22551
rect 58262 22499 58351 22551
rect 57909 22333 58351 22499
rect 57909 22281 57998 22333
rect 58050 22281 58210 22333
rect 58262 22281 58351 22333
rect 57909 22115 58351 22281
rect 57909 22063 57998 22115
rect 58050 22063 58210 22115
rect 58262 22063 58351 22115
rect 57909 21898 58351 22063
rect 57909 21846 57998 21898
rect 58050 21846 58210 21898
rect 58262 21846 58351 21898
rect 57909 21680 58351 21846
rect 57909 21628 57998 21680
rect 58050 21628 58210 21680
rect 58262 21628 58351 21680
rect 57909 21463 58351 21628
rect 57909 21411 57998 21463
rect 58050 21411 58210 21463
rect 58262 21411 58351 21463
rect 57909 21245 58351 21411
rect 57909 21193 57998 21245
rect 58050 21193 58210 21245
rect 58262 21193 58351 21245
rect 57909 21027 58351 21193
rect 57909 20975 57998 21027
rect 58050 20975 58210 21027
rect 58262 20975 58351 21027
rect 57909 20810 58351 20975
rect 57909 20758 57998 20810
rect 58050 20758 58210 20810
rect 58262 20758 58351 20810
rect 57909 20592 58351 20758
rect 57909 20540 57998 20592
rect 58050 20540 58210 20592
rect 58262 20540 58351 20592
rect 57909 20374 58351 20540
rect 57909 20322 57998 20374
rect 58050 20322 58210 20374
rect 58262 20322 58351 20374
rect 57909 20157 58351 20322
rect 57909 20105 57998 20157
rect 58050 20105 58210 20157
rect 58262 20105 58351 20157
rect 57909 19939 58351 20105
rect 57909 19887 57998 19939
rect 58050 19887 58210 19939
rect 58262 19887 58351 19939
rect 57909 19722 58351 19887
rect 57909 19670 57998 19722
rect 58050 19670 58210 19722
rect 58262 19670 58351 19722
rect 57909 19504 58351 19670
rect 57909 19452 57998 19504
rect 58050 19452 58210 19504
rect 58262 19452 58351 19504
rect 57909 19286 58351 19452
rect 57909 19234 57998 19286
rect 58050 19234 58210 19286
rect 58262 19234 58351 19286
rect 57909 19068 58351 19234
rect 57909 19016 57998 19068
rect 58050 19016 58210 19068
rect 58262 19016 58351 19068
rect 57909 18851 58351 19016
rect 57909 18799 57998 18851
rect 58050 18799 58210 18851
rect 58262 18799 58351 18851
rect 57909 18633 58351 18799
rect 57909 18581 57998 18633
rect 58050 18581 58210 18633
rect 58262 18581 58351 18633
rect 57909 18416 58351 18581
rect 57909 18364 57998 18416
rect 58050 18364 58210 18416
rect 58262 18364 58351 18416
rect 57909 18198 58351 18364
rect 57909 18146 57998 18198
rect 58050 18146 58210 18198
rect 58262 18146 58351 18198
rect 57909 17980 58351 18146
rect 57909 17928 57998 17980
rect 58050 17928 58210 17980
rect 58262 17928 58351 17980
rect 57909 17763 58351 17928
rect 57909 17711 57998 17763
rect 58050 17711 58210 17763
rect 58262 17711 58351 17763
rect 57909 17545 58351 17711
rect 57909 17493 57998 17545
rect 58050 17493 58210 17545
rect 58262 17493 58351 17545
rect 57909 17327 58351 17493
rect 57909 17275 57998 17327
rect 58050 17275 58210 17327
rect 58262 17275 58351 17327
rect 57909 17110 58351 17275
rect 57909 17058 57998 17110
rect 58050 17058 58210 17110
rect 58262 17058 58351 17110
rect 57909 16892 58351 17058
rect 57909 16840 57998 16892
rect 58050 16840 58210 16892
rect 58262 16840 58351 16892
rect 57909 16675 58351 16840
rect 57909 16623 57998 16675
rect 58050 16623 58210 16675
rect 58262 16623 58351 16675
rect 57909 16457 58351 16623
rect 57909 16405 57998 16457
rect 58050 16405 58210 16457
rect 58262 16405 58351 16457
rect 57909 16239 58351 16405
rect 57909 16187 57998 16239
rect 58050 16187 58210 16239
rect 58262 16187 58351 16239
rect 57909 16022 58351 16187
rect 57909 15970 57998 16022
rect 58050 15970 58210 16022
rect 58262 15970 58351 16022
rect 57909 15804 58351 15970
rect 57909 15752 57998 15804
rect 58050 15752 58210 15804
rect 58262 15752 58351 15804
rect 57909 15586 58351 15752
rect 57909 15534 57998 15586
rect 58050 15534 58210 15586
rect 58262 15534 58351 15586
rect 57909 15369 58351 15534
rect 57909 15317 57998 15369
rect 58050 15317 58210 15369
rect 58262 15317 58351 15369
rect 57909 15151 58351 15317
rect 57909 15099 57998 15151
rect 58050 15099 58210 15151
rect 58262 15099 58351 15151
rect 57909 14933 58351 15099
rect 57909 14881 57998 14933
rect 58050 14881 58210 14933
rect 58262 14881 58351 14933
rect 57909 14716 58351 14881
rect 57909 14664 57998 14716
rect 58050 14664 58210 14716
rect 58262 14664 58351 14716
rect 57909 14498 58351 14664
rect 57909 14446 57998 14498
rect 58050 14446 58210 14498
rect 58262 14446 58351 14498
rect 57909 14281 58351 14446
rect 57909 14229 57998 14281
rect 58050 14229 58210 14281
rect 58262 14229 58351 14281
rect 57909 14063 58351 14229
rect 57909 14011 57998 14063
rect 58050 14011 58210 14063
rect 58262 14011 58351 14063
rect 57909 13845 58351 14011
rect 57909 13793 57998 13845
rect 58050 13793 58210 13845
rect 58262 13793 58351 13845
rect 57909 13628 58351 13793
rect 57909 13576 57998 13628
rect 58050 13576 58210 13628
rect 58262 13576 58351 13628
rect 57909 13410 58351 13576
rect 57909 13358 57998 13410
rect 58050 13358 58210 13410
rect 58262 13358 58351 13410
rect 57909 13192 58351 13358
rect 57909 13140 57998 13192
rect 58050 13140 58210 13192
rect 58262 13140 58351 13192
rect 57909 12975 58351 13140
rect 57909 12923 57998 12975
rect 58050 12923 58210 12975
rect 58262 12923 58351 12975
rect 57909 12757 58351 12923
rect 57909 12705 57998 12757
rect 58050 12705 58210 12757
rect 58262 12705 58351 12757
rect 57909 12540 58351 12705
rect 57909 12488 57998 12540
rect 58050 12488 58210 12540
rect 58262 12488 58351 12540
rect 57909 12322 58351 12488
rect 57909 12270 57998 12322
rect 58050 12270 58210 12322
rect 58262 12270 58351 12322
rect 57909 12104 58351 12270
rect 57909 12052 57998 12104
rect 58050 12052 58210 12104
rect 58262 12052 58351 12104
rect 57909 11887 58351 12052
rect 57909 11835 57998 11887
rect 58050 11835 58210 11887
rect 58262 11835 58351 11887
rect 57909 11669 58351 11835
rect 57909 11617 57998 11669
rect 58050 11617 58210 11669
rect 58262 11617 58351 11669
rect 57909 11451 58351 11617
rect 57909 11399 57998 11451
rect 58050 11399 58210 11451
rect 58262 11399 58351 11451
rect 57909 11234 58351 11399
rect 57909 11182 57998 11234
rect 58050 11182 58210 11234
rect 58262 11182 58351 11234
rect 57909 11016 58351 11182
rect 57909 10964 57998 11016
rect 58050 10964 58210 11016
rect 58262 10964 58351 11016
rect 57909 10798 58351 10964
rect 57909 10746 57998 10798
rect 58050 10746 58210 10798
rect 58262 10746 58351 10798
rect 57909 10581 58351 10746
rect 57909 10529 57998 10581
rect 58050 10529 58210 10581
rect 58262 10529 58351 10581
rect 57909 10363 58351 10529
rect 57909 10311 57998 10363
rect 58050 10311 58210 10363
rect 58262 10311 58351 10363
rect 57909 10146 58351 10311
rect 57909 10094 57998 10146
rect 58050 10094 58210 10146
rect 58262 10094 58351 10146
rect 57909 9928 58351 10094
rect 57909 9876 57998 9928
rect 58050 9876 58210 9928
rect 58262 9876 58351 9928
rect 57909 9710 58351 9876
rect 57909 9658 57998 9710
rect 58050 9658 58210 9710
rect 58262 9658 58351 9710
rect 57909 9493 58351 9658
rect 57909 9441 57998 9493
rect 58050 9441 58210 9493
rect 58262 9441 58351 9493
rect 57909 9275 58351 9441
rect 57909 9223 57998 9275
rect 58050 9223 58210 9275
rect 58262 9223 58351 9275
rect 57909 9057 58351 9223
rect 57909 9005 57998 9057
rect 58050 9005 58210 9057
rect 58262 9005 58351 9057
rect 57909 8840 58351 9005
rect 57909 8788 57998 8840
rect 58050 8788 58210 8840
rect 58262 8788 58351 8840
rect 57909 8622 58351 8788
rect 57909 8570 57998 8622
rect 58050 8570 58210 8622
rect 58262 8570 58351 8622
rect 57909 8404 58351 8570
rect 57909 8352 57998 8404
rect 58050 8352 58210 8404
rect 58262 8352 58351 8404
rect 57909 8187 58351 8352
rect 57909 8135 57998 8187
rect 58050 8135 58210 8187
rect 58262 8135 58351 8187
rect 57909 7969 58351 8135
rect 57909 7917 57998 7969
rect 58050 7917 58210 7969
rect 58262 7917 58351 7969
rect 57909 7752 58351 7917
rect 57909 7700 57998 7752
rect 58050 7700 58210 7752
rect 58262 7700 58351 7752
rect 57909 7534 58351 7700
rect 57909 7482 57998 7534
rect 58050 7482 58210 7534
rect 58262 7482 58351 7534
rect 57909 7316 58351 7482
rect 57909 7264 57998 7316
rect 58050 7264 58210 7316
rect 58262 7264 58351 7316
rect 57909 7099 58351 7264
rect 57909 7047 57998 7099
rect 58050 7047 58210 7099
rect 58262 7047 58351 7099
rect 57909 6881 58351 7047
rect 57909 6829 57998 6881
rect 58050 6829 58210 6881
rect 58262 6829 58351 6881
rect 57909 6663 58351 6829
rect 57909 6611 57998 6663
rect 58050 6611 58210 6663
rect 58262 6611 58351 6663
rect 57909 6446 58351 6611
rect 57909 6394 57998 6446
rect 58050 6394 58210 6446
rect 58262 6394 58351 6446
rect 57909 6228 58351 6394
rect 57909 6176 57998 6228
rect 58050 6176 58210 6228
rect 58262 6176 58351 6228
rect 57909 6011 58351 6176
rect 57909 5959 57998 6011
rect 58050 5959 58210 6011
rect 58262 5959 58351 6011
rect 57909 5793 58351 5959
rect 57909 5741 57998 5793
rect 58050 5741 58210 5793
rect 58262 5741 58351 5793
rect 57909 5575 58351 5741
rect 57909 5523 57998 5575
rect 58050 5523 58210 5575
rect 58262 5523 58351 5575
rect 57909 5358 58351 5523
rect 57909 5306 57998 5358
rect 58050 5306 58210 5358
rect 58262 5306 58351 5358
rect 61277 5479 61457 5491
rect 61277 5323 61289 5479
rect 61445 5323 61457 5479
rect 61277 5311 61457 5323
rect 57909 4587 58351 5306
rect 57909 4535 57998 4587
rect 58050 4535 58210 4587
rect 58262 4535 58351 4587
rect 57909 4370 58351 4535
rect 57909 4318 57998 4370
rect 58050 4318 58210 4370
rect 58262 4318 58351 4370
rect 57909 4152 58351 4318
rect 57909 4100 57998 4152
rect 58050 4100 58210 4152
rect 58262 4100 58351 4152
rect 57909 3934 58351 4100
rect 57909 3882 57998 3934
rect 58050 3882 58210 3934
rect 58262 3882 58351 3934
rect 57909 3717 58351 3882
rect 57909 3665 57998 3717
rect 58050 3665 58210 3717
rect 58262 3665 58351 3717
rect 57909 1777 58351 3665
rect 27387 1702 57736 1772
rect 2562 1689 2742 1701
rect 2562 1637 2574 1689
rect 2730 1637 2742 1689
rect 2562 1625 2742 1637
rect 12627 1689 12807 1701
rect 12627 1637 12639 1689
rect 12795 1637 12807 1689
rect 12627 1625 12807 1637
rect 13077 1689 13257 1701
rect 13077 1637 13089 1689
rect 13245 1637 13257 1689
rect 13077 1625 13257 1637
rect 23427 1689 23607 1701
rect 23427 1637 23439 1689
rect 23595 1637 23607 1689
rect 23427 1625 23607 1637
rect 27387 1656 28639 1702
rect 28685 1656 28755 1702
rect 28801 1656 28871 1702
rect 28917 1656 28987 1702
rect 29033 1656 29103 1702
rect 29149 1656 29219 1702
rect 29265 1656 29335 1702
rect 29381 1656 29451 1702
rect 29497 1656 29567 1702
rect 29613 1656 29683 1702
rect 29729 1656 29799 1702
rect 29845 1656 29915 1702
rect 29961 1656 30031 1702
rect 30077 1656 30147 1702
rect 30193 1656 30263 1702
rect 30309 1656 30379 1702
rect 30425 1656 30495 1702
rect 30541 1656 30611 1702
rect 30657 1656 30727 1702
rect 30773 1656 30843 1702
rect 30889 1656 30959 1702
rect 31005 1656 31075 1702
rect 31121 1656 31191 1702
rect 31237 1656 31307 1702
rect 31353 1656 31423 1702
rect 31469 1656 31539 1702
rect 31585 1656 31655 1702
rect 31701 1656 31771 1702
rect 31817 1656 31887 1702
rect 31933 1656 32003 1702
rect 32049 1656 32119 1702
rect 32165 1656 32235 1702
rect 32281 1656 32351 1702
rect 32397 1656 32467 1702
rect 32513 1656 32583 1702
rect 32629 1656 32699 1702
rect 32745 1656 32815 1702
rect 32861 1656 32931 1702
rect 32977 1656 33047 1702
rect 33093 1656 33163 1702
rect 33209 1656 33279 1702
rect 33325 1656 33395 1702
rect 33441 1656 33511 1702
rect 33557 1656 33627 1702
rect 33673 1656 33743 1702
rect 33789 1656 33859 1702
rect 33905 1656 33975 1702
rect 34021 1656 34091 1702
rect 34137 1656 34207 1702
rect 34253 1656 34323 1702
rect 34369 1656 34439 1702
rect 34485 1656 34555 1702
rect 34601 1656 34671 1702
rect 34717 1656 34787 1702
rect 34833 1656 34903 1702
rect 34949 1656 35019 1702
rect 35065 1656 35135 1702
rect 35181 1656 35251 1702
rect 35297 1656 35367 1702
rect 35413 1656 35483 1702
rect 35529 1656 35599 1702
rect 35645 1656 35715 1702
rect 35761 1656 35831 1702
rect 35877 1656 35947 1702
rect 35993 1656 36063 1702
rect 36109 1656 36179 1702
rect 36225 1656 36295 1702
rect 36341 1656 36411 1702
rect 36457 1656 36527 1702
rect 36573 1656 36643 1702
rect 36689 1656 36759 1702
rect 36805 1656 36875 1702
rect 36921 1656 36991 1702
rect 37037 1656 37107 1702
rect 37153 1656 37223 1702
rect 37269 1656 37339 1702
rect 37385 1656 37455 1702
rect 37501 1656 37571 1702
rect 37617 1656 37687 1702
rect 37733 1656 37803 1702
rect 37849 1656 37919 1702
rect 37965 1656 38035 1702
rect 38081 1656 38151 1702
rect 38197 1656 38267 1702
rect 38313 1656 38383 1702
rect 38429 1656 38499 1702
rect 38545 1656 38615 1702
rect 38661 1656 38731 1702
rect 38777 1656 38847 1702
rect 38893 1656 38963 1702
rect 39009 1656 39079 1702
rect 39125 1656 39195 1702
rect 39241 1656 39311 1702
rect 39357 1656 39427 1702
rect 39473 1656 39543 1702
rect 39589 1656 39659 1702
rect 39705 1656 39775 1702
rect 39821 1656 39891 1702
rect 39937 1656 40007 1702
rect 40053 1656 40123 1702
rect 40169 1656 50845 1702
rect 50891 1656 50961 1702
rect 51007 1656 51077 1702
rect 51123 1656 51193 1702
rect 51239 1656 51309 1702
rect 51355 1656 51425 1702
rect 51471 1656 51541 1702
rect 51587 1656 51657 1702
rect 51703 1656 51773 1702
rect 51819 1656 51889 1702
rect 51935 1656 52005 1702
rect 52051 1656 52121 1702
rect 52167 1656 52237 1702
rect 52283 1656 52353 1702
rect 52399 1656 52469 1702
rect 52515 1656 52585 1702
rect 52631 1656 52701 1702
rect 52747 1656 52817 1702
rect 52863 1656 52933 1702
rect 52979 1656 53049 1702
rect 53095 1656 53165 1702
rect 53211 1656 53281 1702
rect 53327 1656 53397 1702
rect 53443 1656 53513 1702
rect 53559 1656 53629 1702
rect 53675 1656 53745 1702
rect 53791 1656 53861 1702
rect 53907 1656 53977 1702
rect 54023 1656 54093 1702
rect 54139 1656 54209 1702
rect 54255 1656 54325 1702
rect 54371 1656 54441 1702
rect 54487 1656 54557 1702
rect 54603 1656 54673 1702
rect 54719 1656 54789 1702
rect 54835 1656 54905 1702
rect 54951 1656 55021 1702
rect 55067 1656 55137 1702
rect 55183 1656 55253 1702
rect 55299 1656 55369 1702
rect 55415 1656 55485 1702
rect 55531 1656 55601 1702
rect 55647 1656 55717 1702
rect 55763 1656 55833 1702
rect 55879 1656 55949 1702
rect 55995 1656 56065 1702
rect 56111 1656 56181 1702
rect 56227 1656 56297 1702
rect 56343 1656 56413 1702
rect 56459 1656 56529 1702
rect 56575 1656 57736 1702
rect 27387 1282 57736 1656
rect 62137 1689 62317 1701
rect 62137 1637 62149 1689
rect 62305 1637 62317 1689
rect 62137 1625 62317 1637
rect 72203 1689 72383 1701
rect 72203 1637 72215 1689
rect 72371 1637 72383 1689
rect 72203 1625 72383 1637
rect 72653 1689 72833 1701
rect 72653 1637 72665 1689
rect 72821 1637 72833 1689
rect 72653 1625 72833 1637
rect 82718 1689 82898 1701
rect 82718 1637 82730 1689
rect 82886 1637 82898 1689
rect 82718 1625 82898 1637
rect 282 917 86090 1282
rect 282 657 29092 917
rect 29144 657 86090 917
rect 282 282 86090 657
<< via1 >>
rect 25380 65862 25432 65914
rect 25504 65862 25556 65914
rect 25628 65862 25680 65914
rect 25752 65862 25804 65914
rect 25876 65862 25928 65914
rect 25380 65738 25432 65790
rect 25504 65738 25556 65790
rect 25628 65738 25680 65790
rect 25752 65738 25804 65790
rect 25876 65738 25928 65790
rect 27790 65801 27842 65853
rect 28001 65801 28053 65853
rect 28212 65801 28264 65853
rect 28423 65801 28475 65853
rect 28634 65801 28686 65853
rect 28845 65801 28897 65853
rect 29056 65801 29108 65853
rect 29582 65801 29634 65853
rect 29793 65850 29845 65853
rect 29793 65804 29798 65850
rect 29798 65804 29844 65850
rect 29844 65804 29845 65850
rect 29793 65801 29845 65804
rect 30005 65801 30057 65853
rect 30216 65801 30268 65853
rect 30807 65836 30859 65853
rect 31018 65836 31070 65853
rect 30807 65801 30854 65836
rect 30854 65801 30859 65836
rect 31018 65801 31058 65836
rect 31058 65801 31070 65836
rect 31229 65801 31281 65853
rect 31440 65836 31492 65853
rect 31651 65836 31703 65853
rect 31440 65801 31487 65836
rect 31487 65801 31492 65836
rect 31651 65801 31691 65836
rect 31691 65801 31703 65836
rect 31861 65801 31913 65853
rect 32072 65836 32124 65853
rect 32283 65836 32335 65853
rect 32072 65801 32119 65836
rect 32119 65801 32124 65836
rect 32283 65801 32323 65836
rect 32323 65801 32335 65836
rect 32494 65801 32546 65853
rect 30807 65627 30854 65635
rect 30854 65627 30859 65635
rect 31018 65627 31058 65635
rect 31058 65627 31070 65635
rect 30807 65583 30859 65627
rect 31018 65583 31070 65627
rect 31229 65583 31281 65635
rect 31440 65627 31487 65635
rect 31487 65627 31492 65635
rect 31651 65627 31691 65635
rect 31691 65627 31703 65635
rect 31440 65583 31492 65627
rect 31651 65583 31703 65627
rect 31861 65583 31913 65635
rect 32072 65627 32119 65635
rect 32119 65627 32124 65635
rect 32283 65627 32323 65635
rect 32323 65627 32335 65635
rect 32072 65583 32124 65627
rect 32283 65583 32335 65627
rect 32494 65583 32546 65635
rect 34290 65801 34342 65853
rect 34501 65801 34553 65853
rect 34712 65801 34764 65853
rect 34923 65801 34975 65853
rect 35443 65818 35495 65833
rect 35654 65818 35706 65833
rect 35865 65818 35917 65833
rect 36076 65818 36128 65833
rect 36287 65818 36339 65833
rect 35443 65781 35495 65818
rect 35654 65781 35706 65818
rect 35865 65781 35917 65818
rect 36076 65781 36128 65818
rect 36287 65781 36339 65818
rect 40252 65806 40304 65858
rect 40432 65806 40484 65858
rect 42710 65863 42717 65905
rect 42717 65863 42762 65905
rect 42710 65853 42762 65863
rect 42921 65853 42973 65905
rect 43132 65853 43184 65905
rect 34290 65583 34342 65635
rect 34501 65594 34553 65635
rect 34712 65594 34764 65635
rect 34923 65594 34975 65635
rect 34501 65583 34552 65594
rect 34552 65583 34553 65594
rect 34712 65583 34758 65594
rect 34758 65583 34764 65594
rect 34923 65583 34964 65594
rect 34964 65583 34975 65594
rect 30807 65366 30859 65418
rect 31018 65366 31070 65418
rect 31229 65366 31281 65418
rect 31440 65366 31492 65418
rect 31651 65366 31703 65418
rect 31861 65366 31913 65418
rect 32072 65366 32124 65418
rect 32283 65366 32335 65418
rect 32494 65366 32546 65418
rect 39053 65594 39105 65601
rect 39264 65594 39316 65601
rect 39475 65594 39527 65601
rect 42246 65792 42298 65844
rect 42458 65843 42510 65844
rect 42458 65797 42459 65843
rect 42459 65797 42510 65843
rect 43777 65853 43829 65905
rect 43988 65853 44040 65905
rect 44199 65853 44251 65905
rect 44410 65853 44462 65905
rect 42458 65792 42510 65797
rect 40252 65594 40304 65640
rect 40432 65594 40484 65640
rect 39053 65549 39102 65594
rect 39102 65549 39105 65594
rect 39264 65549 39310 65594
rect 39310 65549 39316 65594
rect 39475 65549 39518 65594
rect 39518 65549 39527 65594
rect 40252 65588 40303 65594
rect 40303 65588 40304 65594
rect 40432 65588 40463 65594
rect 40463 65588 40484 65594
rect 33050 65370 33102 65372
rect 33261 65370 33313 65372
rect 33472 65370 33524 65372
rect 33683 65370 33735 65372
rect 33894 65370 33946 65372
rect 48828 65818 48880 65833
rect 49039 65818 49091 65833
rect 49250 65818 49302 65833
rect 49461 65818 49513 65833
rect 48828 65781 48880 65818
rect 49039 65781 49053 65818
rect 49053 65781 49091 65818
rect 49250 65781 49259 65818
rect 49259 65781 49302 65818
rect 49461 65781 49465 65818
rect 49465 65781 49511 65818
rect 49511 65781 49513 65818
rect 50137 65801 50189 65853
rect 50348 65801 50400 65853
rect 50559 65801 50611 65853
rect 50770 65801 50822 65853
rect 50137 65594 50189 65635
rect 50348 65594 50400 65635
rect 50559 65594 50611 65635
rect 50770 65594 50822 65635
rect 33050 65324 33102 65370
rect 33261 65324 33313 65370
rect 33472 65324 33524 65370
rect 33683 65324 33735 65370
rect 33894 65324 33934 65370
rect 33934 65324 33946 65370
rect 35443 65324 35495 65370
rect 35654 65324 35706 65370
rect 35865 65324 35917 65370
rect 36076 65324 36128 65370
rect 36287 65324 36339 65370
rect 41010 65325 41022 65370
rect 41022 65325 41062 65370
rect 41221 65325 41228 65370
rect 41228 65325 41273 65370
rect 41432 65325 41436 65370
rect 41436 65325 41484 65370
rect 41643 65325 41644 65370
rect 41644 65325 41695 65370
rect 33050 65320 33102 65324
rect 33261 65320 33313 65324
rect 33472 65320 33524 65324
rect 33683 65320 33735 65324
rect 33894 65320 33946 65324
rect 35443 65318 35495 65324
rect 35654 65318 35706 65324
rect 35865 65318 35917 65324
rect 36076 65318 36128 65324
rect 36287 65318 36339 65324
rect 41010 65318 41062 65325
rect 41221 65318 41273 65325
rect 41432 65318 41484 65325
rect 41643 65318 41695 65325
rect 41854 65318 41906 65370
rect 42064 65318 42116 65370
rect 50137 65583 50189 65594
rect 50348 65583 50400 65594
rect 50559 65583 50611 65594
rect 50770 65583 50774 65594
rect 50774 65583 50822 65594
rect 52576 65801 52628 65853
rect 52787 65836 52839 65853
rect 52998 65836 53050 65853
rect 52787 65801 52799 65836
rect 52799 65801 52839 65836
rect 52998 65801 53003 65836
rect 53003 65801 53050 65836
rect 53209 65801 53261 65853
rect 53419 65836 53471 65853
rect 53630 65836 53682 65853
rect 53419 65801 53431 65836
rect 53431 65801 53471 65836
rect 53630 65801 53635 65836
rect 53635 65801 53682 65836
rect 53841 65801 53893 65853
rect 54052 65836 54104 65853
rect 54263 65836 54315 65853
rect 54052 65801 54064 65836
rect 54064 65801 54104 65836
rect 54263 65801 54268 65836
rect 54268 65801 54315 65836
rect 54855 65801 54907 65853
rect 55066 65801 55118 65853
rect 55278 65850 55330 65853
rect 55278 65804 55279 65850
rect 55279 65804 55325 65850
rect 55325 65804 55330 65850
rect 55278 65801 55330 65804
rect 55489 65801 55541 65853
rect 56015 65801 56067 65853
rect 56226 65801 56278 65853
rect 56437 65801 56489 65853
rect 56648 65801 56700 65853
rect 56859 65801 56911 65853
rect 57070 65801 57122 65853
rect 57281 65801 57333 65853
rect 52576 65583 52628 65635
rect 52787 65627 52799 65635
rect 52799 65627 52839 65635
rect 52998 65627 53003 65635
rect 53003 65627 53050 65635
rect 52787 65583 52839 65627
rect 52998 65583 53050 65627
rect 53209 65583 53261 65635
rect 53419 65627 53431 65635
rect 53431 65627 53471 65635
rect 53630 65627 53635 65635
rect 53635 65627 53682 65635
rect 53419 65583 53471 65627
rect 53630 65583 53682 65627
rect 53841 65583 53893 65635
rect 54052 65627 54064 65635
rect 54064 65627 54104 65635
rect 54263 65627 54268 65635
rect 54268 65627 54315 65635
rect 54052 65583 54104 65627
rect 54263 65583 54315 65627
rect 48828 65324 48880 65370
rect 49039 65324 49053 65370
rect 49053 65324 49091 65370
rect 49250 65324 49259 65370
rect 49259 65324 49302 65370
rect 49461 65324 49465 65370
rect 49465 65324 49511 65370
rect 49511 65324 49513 65370
rect 51081 65324 51083 65370
rect 51083 65324 51133 65370
rect 48828 65318 48880 65324
rect 49039 65318 49091 65324
rect 49250 65318 49302 65324
rect 49461 65318 49513 65324
rect 51081 65318 51133 65324
rect 51292 65318 51344 65370
rect 51503 65324 51552 65370
rect 51552 65324 51555 65370
rect 51714 65324 51758 65370
rect 51758 65324 51766 65370
rect 51925 65324 51964 65370
rect 51964 65324 51977 65370
rect 52576 65366 52628 65418
rect 52787 65366 52839 65418
rect 52998 65366 53050 65418
rect 53209 65366 53261 65418
rect 53419 65366 53471 65418
rect 53630 65366 53682 65418
rect 53841 65366 53893 65418
rect 54052 65366 54104 65418
rect 54263 65366 54315 65418
rect 51503 65318 51555 65324
rect 51714 65318 51766 65324
rect 51925 65318 51977 65324
rect 29582 64901 29634 64953
rect 29793 64950 29845 64953
rect 29793 64904 29798 64950
rect 29798 64904 29844 64950
rect 29844 64904 29845 64950
rect 29793 64901 29845 64904
rect 30005 64901 30057 64953
rect 30216 64901 30268 64953
rect 30854 64901 30906 64953
rect 31065 64901 31117 64953
rect 31276 64901 31328 64953
rect 31486 64950 31538 64953
rect 31697 64950 31749 64953
rect 31909 64950 31961 64953
rect 32120 64950 32172 64953
rect 32330 64950 32382 64953
rect 32541 64950 32593 64953
rect 32752 64950 32804 64953
rect 34284 64950 34336 64953
rect 34495 64950 34547 64953
rect 31486 64904 31538 64950
rect 31697 64904 31749 64950
rect 31909 64904 31961 64950
rect 32120 64904 32172 64950
rect 32330 64904 32382 64950
rect 32541 64904 32593 64950
rect 32752 64904 32804 64950
rect 34284 64904 34302 64950
rect 34302 64904 34336 64950
rect 34495 64904 34508 64950
rect 34508 64904 34547 64950
rect 31486 64901 31538 64904
rect 31697 64901 31749 64904
rect 31909 64901 31961 64904
rect 32120 64901 32172 64904
rect 32330 64901 32382 64904
rect 32541 64901 32593 64904
rect 32752 64901 32804 64904
rect 34284 64901 34336 64904
rect 34495 64901 34547 64904
rect 34707 64901 34759 64953
rect 34918 64901 34970 64953
rect 35220 64901 35272 64953
rect 35430 64901 35482 64953
rect 35641 64901 35693 64953
rect 35853 64901 35905 64953
rect 36064 64901 36116 64953
rect 36274 64901 36326 64953
rect 38330 64950 38382 64953
rect 38330 64904 38382 64950
rect 38330 64901 38382 64904
rect 38541 64901 38593 64953
rect 38752 64901 38804 64953
rect 58858 65862 58910 65914
rect 58982 65862 59034 65914
rect 59106 65862 59158 65914
rect 59230 65862 59282 65914
rect 59354 65862 59406 65914
rect 58858 65738 58910 65790
rect 58982 65738 59034 65790
rect 59106 65738 59158 65790
rect 59230 65738 59282 65790
rect 59354 65738 59406 65790
rect 39052 64950 39104 64953
rect 39232 64950 39284 64953
rect 39052 64904 39062 64950
rect 39062 64904 39104 64950
rect 39232 64904 39266 64950
rect 39266 64904 39284 64950
rect 39052 64901 39104 64904
rect 39232 64901 39284 64904
rect 33057 64726 33109 64729
rect 33237 64726 33289 64729
rect 33057 64680 33109 64726
rect 33237 64680 33289 64726
rect 33057 64677 33109 64680
rect 33237 64677 33289 64680
rect 33819 64726 33871 64737
rect 33999 64726 34051 64737
rect 33819 64685 33833 64726
rect 33833 64685 33871 64726
rect 33999 64685 34039 64726
rect 34039 64685 34051 64726
rect 35332 64639 35384 64651
rect 35543 64639 35595 64651
rect 35754 64639 35806 64651
rect 35965 64639 36017 64651
rect 36176 64639 36228 64651
rect 37891 64639 37943 64663
rect 38071 64639 38123 64663
rect 35332 64599 35384 64639
rect 35543 64599 35580 64639
rect 35580 64599 35595 64639
rect 35754 64599 35786 64639
rect 35786 64599 35806 64639
rect 35965 64599 35992 64639
rect 35992 64599 36017 64639
rect 36176 64599 36198 64639
rect 36198 64599 36228 64639
rect 37891 64611 37909 64639
rect 37909 64611 37943 64639
rect 38071 64611 38072 64639
rect 38072 64611 38123 64639
rect 34267 64456 34302 64491
rect 34302 64456 34319 64491
rect 34447 64456 34451 64491
rect 34451 64456 34499 64491
rect 34627 64456 34658 64491
rect 34658 64456 34679 64491
rect 34267 64439 34319 64456
rect 34447 64439 34499 64456
rect 34627 64439 34679 64456
rect 33057 64278 33109 64281
rect 33237 64278 33289 64281
rect 33057 64232 33109 64278
rect 33237 64232 33289 64278
rect 33057 64229 33109 64232
rect 33237 64229 33289 64232
rect 36678 64364 36697 64416
rect 36697 64364 36730 64416
rect 36961 64415 37013 64423
rect 37172 64415 37224 64423
rect 36961 64371 36971 64415
rect 36971 64371 37013 64415
rect 37172 64371 37206 64415
rect 37206 64371 37224 64415
rect 37384 64371 37436 64423
rect 37595 64371 37647 64423
rect 40253 64901 40305 64953
rect 40433 64901 40485 64953
rect 43790 64901 43842 64953
rect 44001 64901 44053 64953
rect 44213 64950 44265 64953
rect 44213 64904 44236 64950
rect 44236 64904 44265 64950
rect 44213 64901 44265 64904
rect 44424 64901 44476 64953
rect 44834 64950 44886 64953
rect 45045 64950 45097 64953
rect 45256 64950 45308 64953
rect 44834 64904 44858 64950
rect 44858 64904 44886 64950
rect 45045 64904 45084 64950
rect 45084 64904 45097 64950
rect 45256 64904 45264 64950
rect 45264 64904 45308 64950
rect 44834 64901 44886 64904
rect 45045 64901 45097 64904
rect 45256 64901 45308 64904
rect 48838 64901 48890 64953
rect 49048 64901 49100 64953
rect 49259 64901 49311 64953
rect 49471 64901 49523 64953
rect 49682 64901 49734 64953
rect 49892 64901 49944 64953
rect 50346 64901 50398 64953
rect 50557 64950 50609 64953
rect 50768 64950 50820 64953
rect 52316 64950 52368 64953
rect 52527 64950 52579 64953
rect 52738 64950 52790 64953
rect 52948 64950 53000 64953
rect 53159 64950 53211 64953
rect 53371 64950 53423 64953
rect 53582 64950 53634 64953
rect 50557 64904 50571 64950
rect 50571 64904 50609 64950
rect 50768 64904 50777 64950
rect 50777 64904 50820 64950
rect 52316 64904 52368 64950
rect 52527 64904 52579 64950
rect 52738 64904 52790 64950
rect 52948 64904 53000 64950
rect 53159 64904 53211 64950
rect 53371 64904 53423 64950
rect 53582 64904 53634 64950
rect 50557 64901 50609 64904
rect 50768 64901 50820 64904
rect 39775 64680 39786 64715
rect 39786 64680 39827 64715
rect 39775 64663 39827 64680
rect 39994 64448 40046 64500
rect 39994 64262 40046 64314
rect 52316 64901 52368 64904
rect 52527 64901 52579 64904
rect 52738 64901 52790 64904
rect 52948 64901 53000 64904
rect 53159 64901 53211 64904
rect 53371 64901 53423 64904
rect 53582 64901 53634 64904
rect 53792 64901 53844 64953
rect 54003 64901 54055 64953
rect 54214 64901 54266 64953
rect 54855 64901 54907 64953
rect 55066 64901 55118 64953
rect 55278 64950 55330 64953
rect 55278 64904 55279 64950
rect 55279 64904 55325 64950
rect 55325 64904 55330 64950
rect 55278 64901 55330 64904
rect 55489 64901 55541 64953
rect 41935 64663 41987 64715
rect 51073 64726 51125 64729
rect 51253 64726 51305 64729
rect 42312 64432 42364 64484
rect 51073 64680 51086 64726
rect 51086 64680 51125 64726
rect 51253 64680 51292 64726
rect 51292 64680 51305 64726
rect 48943 64639 48995 64654
rect 49154 64639 49206 64654
rect 49365 64639 49417 64654
rect 49576 64639 49628 64654
rect 49787 64639 49839 64654
rect 48943 64602 48984 64639
rect 48984 64602 48995 64639
rect 49154 64602 49190 64639
rect 49190 64602 49206 64639
rect 49365 64602 49396 64639
rect 49396 64602 49417 64639
rect 49576 64602 49602 64639
rect 49602 64602 49628 64639
rect 49787 64602 49839 64639
rect 51073 64677 51125 64680
rect 51253 64677 51305 64680
rect 44939 64456 44971 64491
rect 44971 64456 44991 64491
rect 45151 64456 45197 64491
rect 45197 64456 45203 64491
rect 48596 64495 48648 64547
rect 44939 64439 44991 64456
rect 45151 64439 45203 64456
rect 45597 64337 45604 64375
rect 45604 64337 45649 64375
rect 45597 64323 45649 64337
rect 50300 64439 50352 64491
rect 50511 64456 50513 64491
rect 50513 64456 50563 64491
rect 50511 64439 50563 64456
rect 50722 64439 50774 64491
rect 48596 64277 48648 64329
rect 51835 64680 51887 64722
rect 52015 64680 52067 64722
rect 51835 64670 51887 64680
rect 52015 64670 52067 64680
rect 35332 64145 35384 64191
rect 35543 64145 35580 64191
rect 35580 64145 35595 64191
rect 35754 64145 35786 64191
rect 35786 64145 35806 64191
rect 35965 64145 35992 64191
rect 35992 64145 36017 64191
rect 36176 64145 36198 64191
rect 36198 64145 36228 64191
rect 37891 64145 37909 64189
rect 37909 64145 37943 64189
rect 38071 64145 38072 64189
rect 38072 64145 38123 64189
rect 48943 64145 48984 64191
rect 48984 64145 48995 64191
rect 49154 64145 49190 64191
rect 49190 64145 49206 64191
rect 49365 64145 49396 64191
rect 49396 64145 49417 64191
rect 49576 64145 49602 64191
rect 49602 64145 49628 64191
rect 49787 64145 49839 64191
rect 51835 64232 51887 64259
rect 52015 64232 52067 64259
rect 51835 64207 51887 64232
rect 52015 64207 52067 64232
rect 35332 64139 35384 64145
rect 35543 64139 35595 64145
rect 35754 64139 35806 64145
rect 35965 64139 36017 64145
rect 36176 64139 36228 64145
rect 37891 64137 37943 64145
rect 38071 64137 38123 64145
rect 27790 64001 27842 64053
rect 28001 64001 28053 64053
rect 28212 64001 28264 64053
rect 28423 64001 28475 64053
rect 28634 64001 28686 64053
rect 28845 64050 28897 64053
rect 28845 64004 28856 64050
rect 28856 64004 28897 64050
rect 28845 64001 28897 64004
rect 29056 64001 29108 64053
rect 29582 64001 29634 64053
rect 29793 64050 29845 64053
rect 29793 64004 29798 64050
rect 29798 64004 29844 64050
rect 29844 64004 29845 64050
rect 29793 64001 29845 64004
rect 30005 64001 30057 64053
rect 30216 64001 30268 64053
rect 30854 64001 30906 64053
rect 31065 64001 31117 64053
rect 31276 64001 31328 64053
rect 31486 64001 31538 64053
rect 31697 64001 31749 64053
rect 31909 64001 31961 64053
rect 32120 64001 32172 64053
rect 32330 64001 32382 64053
rect 32541 64001 32593 64053
rect 32752 64001 32804 64053
rect 48943 64139 48995 64145
rect 49154 64139 49206 64145
rect 49365 64139 49417 64145
rect 49576 64139 49628 64145
rect 49787 64139 49839 64145
rect 34755 64001 34807 64053
rect 34935 64050 34987 64053
rect 34935 64004 34962 64050
rect 34962 64004 34987 64050
rect 34935 64001 34987 64004
rect 50138 64050 50190 64053
rect 50138 64004 50160 64050
rect 50160 64004 50190 64050
rect 50138 64001 50190 64004
rect 50318 64001 50370 64053
rect 35332 63909 35384 63915
rect 35543 63909 35595 63915
rect 35754 63909 35806 63915
rect 35965 63909 36017 63915
rect 36176 63909 36228 63915
rect 37891 63909 37943 63917
rect 38071 63909 38123 63917
rect 52316 64001 52368 64053
rect 52527 64001 52579 64053
rect 52738 64001 52790 64053
rect 52948 64001 53000 64053
rect 53159 64001 53211 64053
rect 53371 64001 53423 64053
rect 53582 64001 53634 64053
rect 53792 64001 53844 64053
rect 54003 64001 54055 64053
rect 54214 64001 54266 64053
rect 54855 64001 54907 64053
rect 55066 64001 55118 64053
rect 55278 64050 55330 64053
rect 55278 64004 55279 64050
rect 55279 64004 55325 64050
rect 55325 64004 55330 64050
rect 55278 64001 55330 64004
rect 55489 64001 55541 64053
rect 56015 64001 56067 64053
rect 56226 64050 56278 64053
rect 56226 64004 56267 64050
rect 56267 64004 56278 64050
rect 56226 64001 56278 64004
rect 56437 64001 56489 64053
rect 56648 64001 56700 64053
rect 56859 64001 56911 64053
rect 57070 64001 57122 64053
rect 57281 64001 57333 64053
rect 48943 63909 48995 63915
rect 49154 63909 49206 63915
rect 49365 63909 49417 63915
rect 49576 63909 49628 63915
rect 49787 63909 49839 63915
rect 33057 63822 33109 63825
rect 33237 63822 33289 63825
rect 35332 63863 35384 63909
rect 35543 63863 35580 63909
rect 35580 63863 35595 63909
rect 35754 63863 35786 63909
rect 35786 63863 35806 63909
rect 35965 63863 35992 63909
rect 35992 63863 36017 63909
rect 36176 63863 36198 63909
rect 36198 63863 36228 63909
rect 37891 63865 37909 63909
rect 37909 63865 37943 63909
rect 38071 63865 38072 63909
rect 38072 63865 38123 63909
rect 33057 63776 33109 63822
rect 33237 63776 33289 63822
rect 33057 63773 33109 63776
rect 33237 63773 33289 63776
rect 33057 63374 33109 63377
rect 33237 63374 33289 63377
rect 33057 63328 33109 63374
rect 33237 63328 33289 63374
rect 33057 63325 33109 63328
rect 33237 63325 33289 63328
rect 29582 63101 29634 63153
rect 29793 63150 29845 63153
rect 29793 63104 29798 63150
rect 29798 63104 29844 63150
rect 29844 63104 29845 63150
rect 29793 63101 29845 63104
rect 30005 63101 30057 63153
rect 30216 63101 30268 63153
rect 34267 63598 34319 63615
rect 34447 63598 34499 63615
rect 34627 63598 34679 63615
rect 34267 63563 34302 63598
rect 34302 63563 34319 63598
rect 34447 63563 34451 63598
rect 34451 63563 34499 63598
rect 34627 63563 34658 63598
rect 34658 63563 34679 63598
rect 36678 63638 36697 63690
rect 36697 63638 36730 63690
rect 48943 63863 48984 63909
rect 48984 63863 48995 63909
rect 49154 63863 49190 63909
rect 49190 63863 49206 63909
rect 49365 63863 49396 63909
rect 49396 63863 49417 63909
rect 49576 63863 49602 63909
rect 49602 63863 49628 63909
rect 49787 63863 49839 63909
rect 39994 63740 40046 63792
rect 36961 63639 36971 63683
rect 36971 63639 37013 63683
rect 37172 63639 37206 63683
rect 37206 63639 37224 63683
rect 36961 63631 37013 63639
rect 37172 63631 37224 63639
rect 37384 63631 37436 63683
rect 37595 63631 37647 63683
rect 35332 63415 35384 63455
rect 35543 63415 35580 63455
rect 35580 63415 35595 63455
rect 35754 63415 35786 63455
rect 35786 63415 35806 63455
rect 35965 63415 35992 63455
rect 35992 63415 36017 63455
rect 36176 63415 36198 63455
rect 36198 63415 36228 63455
rect 37891 63415 37909 63443
rect 37909 63415 37943 63443
rect 38071 63415 38072 63443
rect 38072 63415 38123 63443
rect 35332 63403 35384 63415
rect 35543 63403 35595 63415
rect 35754 63403 35806 63415
rect 35965 63403 36017 63415
rect 36176 63403 36228 63415
rect 33819 63328 33833 63369
rect 33833 63328 33871 63369
rect 33999 63328 34039 63369
rect 34039 63328 34051 63369
rect 37891 63391 37943 63415
rect 38071 63391 38123 63415
rect 33819 63317 33871 63328
rect 33999 63317 34051 63328
rect 30854 63101 30906 63153
rect 31065 63101 31117 63153
rect 31276 63101 31328 63153
rect 31486 63150 31538 63153
rect 31697 63150 31749 63153
rect 31909 63150 31961 63153
rect 32120 63150 32172 63153
rect 32330 63150 32382 63153
rect 32541 63150 32593 63153
rect 32752 63150 32804 63153
rect 34284 63150 34336 63153
rect 34495 63150 34547 63153
rect 31486 63104 31538 63150
rect 31697 63104 31749 63150
rect 31909 63104 31961 63150
rect 32120 63104 32172 63150
rect 32330 63104 32382 63150
rect 32541 63104 32593 63150
rect 32752 63104 32804 63150
rect 34284 63104 34302 63150
rect 34302 63104 34336 63150
rect 34495 63104 34508 63150
rect 34508 63104 34547 63150
rect 31486 63101 31538 63104
rect 31697 63101 31749 63104
rect 31909 63101 31961 63104
rect 32120 63101 32172 63104
rect 32330 63101 32382 63104
rect 32541 63101 32593 63104
rect 32752 63101 32804 63104
rect 34284 63101 34336 63104
rect 34495 63101 34547 63104
rect 34707 63101 34759 63153
rect 34918 63101 34970 63153
rect 35220 63101 35272 63153
rect 35430 63101 35482 63153
rect 35641 63101 35693 63153
rect 35853 63101 35905 63153
rect 36064 63101 36116 63153
rect 36274 63101 36326 63153
rect 38330 63150 38382 63153
rect 38330 63104 38382 63150
rect 38330 63101 38382 63104
rect 38541 63101 38593 63153
rect 38752 63101 38804 63153
rect 39052 63150 39104 63153
rect 39232 63150 39284 63153
rect 39052 63104 39062 63150
rect 39062 63104 39104 63150
rect 39232 63104 39266 63150
rect 39266 63104 39284 63150
rect 39052 63101 39104 63104
rect 39232 63101 39284 63104
rect 33057 62926 33109 62929
rect 33237 62926 33289 62929
rect 33057 62880 33109 62926
rect 33237 62880 33289 62926
rect 33057 62877 33109 62880
rect 33237 62877 33289 62880
rect 33819 62926 33871 62937
rect 33999 62926 34051 62937
rect 33819 62885 33833 62926
rect 33833 62885 33871 62926
rect 33999 62885 34039 62926
rect 34039 62885 34051 62926
rect 35332 62839 35384 62851
rect 35543 62839 35595 62851
rect 35754 62839 35806 62851
rect 35965 62839 36017 62851
rect 36176 62839 36228 62851
rect 37891 62839 37943 62863
rect 38071 62839 38123 62863
rect 35332 62799 35384 62839
rect 35543 62799 35580 62839
rect 35580 62799 35595 62839
rect 35754 62799 35786 62839
rect 35786 62799 35806 62839
rect 35965 62799 35992 62839
rect 35992 62799 36017 62839
rect 36176 62799 36198 62839
rect 36198 62799 36228 62839
rect 37891 62811 37909 62839
rect 37909 62811 37943 62839
rect 38071 62811 38072 62839
rect 38072 62811 38123 62839
rect 34267 62656 34302 62691
rect 34302 62656 34319 62691
rect 34447 62656 34451 62691
rect 34451 62656 34499 62691
rect 34627 62656 34658 62691
rect 34658 62656 34679 62691
rect 34267 62639 34319 62656
rect 34447 62639 34499 62656
rect 34627 62639 34679 62656
rect 33057 62478 33109 62481
rect 33237 62478 33289 62481
rect 33057 62432 33109 62478
rect 33237 62432 33289 62478
rect 33057 62429 33109 62432
rect 33237 62429 33289 62432
rect 36678 62564 36697 62616
rect 36697 62564 36730 62616
rect 36961 62615 37013 62623
rect 37172 62615 37224 62623
rect 36961 62571 36971 62615
rect 36971 62571 37013 62615
rect 37172 62571 37206 62615
rect 37206 62571 37224 62615
rect 37384 62571 37436 62623
rect 37595 62571 37647 62623
rect 39994 63554 40046 63606
rect 39775 63374 39827 63391
rect 39775 63339 39786 63374
rect 39786 63339 39827 63374
rect 42312 63570 42364 63622
rect 41935 63339 41987 63391
rect 45975 63679 46027 63731
rect 48596 63725 48648 63777
rect 51835 63822 51887 63847
rect 52015 63822 52067 63847
rect 51835 63795 51887 63822
rect 52015 63795 52067 63822
rect 44939 63598 44991 63615
rect 45151 63598 45203 63615
rect 44939 63563 44971 63598
rect 44971 63563 44991 63598
rect 45151 63563 45197 63598
rect 45197 63563 45203 63598
rect 48596 63507 48648 63559
rect 50300 63563 50352 63615
rect 50511 63598 50563 63615
rect 50511 63563 50513 63598
rect 50513 63563 50563 63598
rect 50722 63563 50774 63615
rect 48943 63415 48984 63452
rect 48984 63415 48995 63452
rect 49154 63415 49190 63452
rect 49190 63415 49206 63452
rect 49365 63415 49396 63452
rect 49396 63415 49417 63452
rect 49576 63415 49602 63452
rect 49602 63415 49628 63452
rect 49787 63415 49839 63452
rect 48943 63400 48995 63415
rect 49154 63400 49206 63415
rect 49365 63400 49417 63415
rect 49576 63400 49628 63415
rect 49787 63400 49839 63415
rect 51073 63374 51125 63377
rect 51253 63374 51305 63377
rect 51073 63328 51086 63374
rect 51086 63328 51125 63374
rect 51253 63328 51292 63374
rect 51292 63328 51305 63374
rect 51073 63325 51125 63328
rect 51253 63325 51305 63328
rect 51835 63374 51887 63384
rect 52015 63374 52067 63384
rect 51835 63332 51887 63374
rect 52015 63332 52067 63374
rect 40253 63101 40305 63153
rect 40433 63101 40485 63153
rect 43790 63101 43842 63153
rect 44001 63101 44053 63153
rect 44213 63150 44265 63153
rect 44213 63104 44236 63150
rect 44236 63104 44265 63150
rect 44213 63101 44265 63104
rect 44424 63101 44476 63153
rect 44834 63150 44886 63153
rect 45045 63150 45097 63153
rect 45256 63150 45308 63153
rect 44834 63104 44858 63150
rect 44858 63104 44886 63150
rect 45045 63104 45084 63150
rect 45084 63104 45097 63150
rect 45256 63104 45264 63150
rect 45264 63104 45308 63150
rect 44834 63101 44886 63104
rect 45045 63101 45097 63104
rect 45256 63101 45308 63104
rect 48838 63101 48890 63153
rect 49048 63101 49100 63153
rect 49259 63101 49311 63153
rect 49471 63101 49523 63153
rect 49682 63101 49734 63153
rect 49892 63101 49944 63153
rect 50346 63101 50398 63153
rect 50557 63150 50609 63153
rect 50768 63150 50820 63153
rect 52316 63150 52368 63153
rect 52527 63150 52579 63153
rect 52738 63150 52790 63153
rect 52948 63150 53000 63153
rect 53159 63150 53211 63153
rect 53371 63150 53423 63153
rect 53582 63150 53634 63153
rect 50557 63104 50571 63150
rect 50571 63104 50609 63150
rect 50768 63104 50777 63150
rect 50777 63104 50820 63150
rect 52316 63104 52368 63150
rect 52527 63104 52579 63150
rect 52738 63104 52790 63150
rect 52948 63104 53000 63150
rect 53159 63104 53211 63150
rect 53371 63104 53423 63150
rect 53582 63104 53634 63150
rect 50557 63101 50609 63104
rect 50768 63101 50820 63104
rect 39775 62880 39786 62915
rect 39786 62880 39827 62915
rect 39775 62863 39827 62880
rect 39994 62648 40046 62700
rect 39994 62462 40046 62514
rect 52316 63101 52368 63104
rect 52527 63101 52579 63104
rect 52738 63101 52790 63104
rect 52948 63101 53000 63104
rect 53159 63101 53211 63104
rect 53371 63101 53423 63104
rect 53582 63101 53634 63104
rect 53792 63101 53844 63153
rect 54003 63101 54055 63153
rect 54214 63101 54266 63153
rect 54855 63101 54907 63153
rect 55066 63101 55118 63153
rect 55278 63150 55330 63153
rect 55278 63104 55279 63150
rect 55279 63104 55325 63150
rect 55325 63104 55330 63150
rect 55278 63101 55330 63104
rect 55489 63101 55541 63153
rect 41935 62863 41987 62915
rect 51073 62926 51125 62929
rect 51253 62926 51305 62929
rect 42312 62632 42364 62684
rect 51073 62880 51086 62926
rect 51086 62880 51125 62926
rect 51253 62880 51292 62926
rect 51292 62880 51305 62926
rect 48943 62839 48995 62854
rect 49154 62839 49206 62854
rect 49365 62839 49417 62854
rect 49576 62839 49628 62854
rect 49787 62839 49839 62854
rect 48943 62802 48984 62839
rect 48984 62802 48995 62839
rect 49154 62802 49190 62839
rect 49190 62802 49206 62839
rect 49365 62802 49396 62839
rect 49396 62802 49417 62839
rect 49576 62802 49602 62839
rect 49602 62802 49628 62839
rect 49787 62802 49839 62839
rect 51073 62877 51125 62880
rect 51253 62877 51305 62880
rect 44939 62656 44971 62691
rect 44971 62656 44991 62691
rect 45151 62656 45197 62691
rect 45197 62656 45203 62691
rect 48596 62695 48648 62747
rect 44939 62639 44991 62656
rect 45151 62639 45203 62656
rect 46353 62523 46405 62575
rect 50300 62639 50352 62691
rect 50511 62656 50513 62691
rect 50513 62656 50563 62691
rect 50511 62639 50563 62656
rect 50722 62639 50774 62691
rect 48596 62477 48648 62529
rect 51835 62880 51887 62922
rect 52015 62880 52067 62922
rect 51835 62870 51887 62880
rect 52015 62870 52067 62880
rect 35332 62345 35384 62391
rect 35543 62345 35580 62391
rect 35580 62345 35595 62391
rect 35754 62345 35786 62391
rect 35786 62345 35806 62391
rect 35965 62345 35992 62391
rect 35992 62345 36017 62391
rect 36176 62345 36198 62391
rect 36198 62345 36228 62391
rect 37891 62345 37909 62389
rect 37909 62345 37943 62389
rect 38071 62345 38072 62389
rect 38072 62345 38123 62389
rect 48943 62345 48984 62391
rect 48984 62345 48995 62391
rect 49154 62345 49190 62391
rect 49190 62345 49206 62391
rect 49365 62345 49396 62391
rect 49396 62345 49417 62391
rect 49576 62345 49602 62391
rect 49602 62345 49628 62391
rect 49787 62345 49839 62391
rect 51835 62432 51887 62459
rect 52015 62432 52067 62459
rect 51835 62407 51887 62432
rect 52015 62407 52067 62432
rect 35332 62339 35384 62345
rect 35543 62339 35595 62345
rect 35754 62339 35806 62345
rect 35965 62339 36017 62345
rect 36176 62339 36228 62345
rect 37891 62337 37943 62345
rect 38071 62337 38123 62345
rect 27790 62201 27842 62253
rect 28001 62201 28053 62253
rect 28212 62201 28264 62253
rect 28423 62201 28475 62253
rect 28634 62201 28686 62253
rect 28845 62250 28897 62253
rect 28845 62204 28856 62250
rect 28856 62204 28897 62250
rect 28845 62201 28897 62204
rect 29056 62201 29108 62253
rect 29582 62201 29634 62253
rect 29793 62250 29845 62253
rect 29793 62204 29798 62250
rect 29798 62204 29844 62250
rect 29844 62204 29845 62250
rect 29793 62201 29845 62204
rect 30005 62201 30057 62253
rect 30216 62201 30268 62253
rect 30854 62201 30906 62253
rect 31065 62201 31117 62253
rect 31276 62201 31328 62253
rect 31486 62201 31538 62253
rect 31697 62201 31749 62253
rect 31909 62201 31961 62253
rect 32120 62201 32172 62253
rect 32330 62201 32382 62253
rect 32541 62201 32593 62253
rect 32752 62201 32804 62253
rect 48943 62339 48995 62345
rect 49154 62339 49206 62345
rect 49365 62339 49417 62345
rect 49576 62339 49628 62345
rect 49787 62339 49839 62345
rect 34755 62201 34807 62253
rect 34935 62250 34987 62253
rect 34935 62204 34962 62250
rect 34962 62204 34987 62250
rect 34935 62201 34987 62204
rect 50138 62250 50190 62253
rect 50138 62204 50160 62250
rect 50160 62204 50190 62250
rect 50138 62201 50190 62204
rect 50318 62201 50370 62253
rect 35332 62109 35384 62115
rect 35543 62109 35595 62115
rect 35754 62109 35806 62115
rect 35965 62109 36017 62115
rect 36176 62109 36228 62115
rect 37891 62109 37943 62117
rect 38071 62109 38123 62117
rect 52316 62201 52368 62253
rect 52527 62201 52579 62253
rect 52738 62201 52790 62253
rect 52948 62201 53000 62253
rect 53159 62201 53211 62253
rect 53371 62201 53423 62253
rect 53582 62201 53634 62253
rect 53792 62201 53844 62253
rect 54003 62201 54055 62253
rect 54214 62201 54266 62253
rect 54855 62201 54907 62253
rect 55066 62201 55118 62253
rect 55278 62250 55330 62253
rect 55278 62204 55279 62250
rect 55279 62204 55325 62250
rect 55325 62204 55330 62250
rect 55278 62201 55330 62204
rect 55489 62201 55541 62253
rect 56015 62201 56067 62253
rect 56226 62250 56278 62253
rect 56226 62204 56267 62250
rect 56267 62204 56278 62250
rect 56226 62201 56278 62204
rect 56437 62201 56489 62253
rect 56648 62201 56700 62253
rect 56859 62201 56911 62253
rect 57070 62201 57122 62253
rect 57281 62201 57333 62253
rect 48943 62109 48995 62115
rect 49154 62109 49206 62115
rect 49365 62109 49417 62115
rect 49576 62109 49628 62115
rect 49787 62109 49839 62115
rect 33057 62022 33109 62025
rect 33237 62022 33289 62025
rect 35332 62063 35384 62109
rect 35543 62063 35580 62109
rect 35580 62063 35595 62109
rect 35754 62063 35786 62109
rect 35786 62063 35806 62109
rect 35965 62063 35992 62109
rect 35992 62063 36017 62109
rect 36176 62063 36198 62109
rect 36198 62063 36228 62109
rect 37891 62065 37909 62109
rect 37909 62065 37943 62109
rect 38071 62065 38072 62109
rect 38072 62065 38123 62109
rect 33057 61976 33109 62022
rect 33237 61976 33289 62022
rect 33057 61973 33109 61976
rect 33237 61973 33289 61976
rect 33057 61574 33109 61577
rect 33237 61574 33289 61577
rect 33057 61528 33109 61574
rect 33237 61528 33289 61574
rect 33057 61525 33109 61528
rect 33237 61525 33289 61528
rect 29582 61301 29634 61353
rect 29793 61350 29845 61353
rect 29793 61304 29798 61350
rect 29798 61304 29844 61350
rect 29844 61304 29845 61350
rect 29793 61301 29845 61304
rect 30005 61301 30057 61353
rect 30216 61301 30268 61353
rect 34267 61798 34319 61815
rect 34447 61798 34499 61815
rect 34627 61798 34679 61815
rect 34267 61763 34302 61798
rect 34302 61763 34319 61798
rect 34447 61763 34451 61798
rect 34451 61763 34499 61798
rect 34627 61763 34658 61798
rect 34658 61763 34679 61798
rect 36678 61838 36697 61890
rect 36697 61838 36730 61890
rect 48943 62063 48984 62109
rect 48984 62063 48995 62109
rect 49154 62063 49190 62109
rect 49190 62063 49206 62109
rect 49365 62063 49396 62109
rect 49396 62063 49417 62109
rect 49576 62063 49602 62109
rect 49602 62063 49628 62109
rect 49787 62063 49839 62109
rect 39994 61940 40046 61992
rect 36961 61839 36971 61883
rect 36971 61839 37013 61883
rect 37172 61839 37206 61883
rect 37206 61839 37224 61883
rect 36961 61831 37013 61839
rect 37172 61831 37224 61839
rect 37384 61831 37436 61883
rect 37595 61831 37647 61883
rect 35332 61615 35384 61655
rect 35543 61615 35580 61655
rect 35580 61615 35595 61655
rect 35754 61615 35786 61655
rect 35786 61615 35806 61655
rect 35965 61615 35992 61655
rect 35992 61615 36017 61655
rect 36176 61615 36198 61655
rect 36198 61615 36228 61655
rect 37891 61615 37909 61643
rect 37909 61615 37943 61643
rect 38071 61615 38072 61643
rect 38072 61615 38123 61643
rect 35332 61603 35384 61615
rect 35543 61603 35595 61615
rect 35754 61603 35806 61615
rect 35965 61603 36017 61615
rect 36176 61603 36228 61615
rect 33819 61528 33833 61569
rect 33833 61528 33871 61569
rect 33999 61528 34039 61569
rect 34039 61528 34051 61569
rect 37891 61591 37943 61615
rect 38071 61591 38123 61615
rect 33819 61517 33871 61528
rect 33999 61517 34051 61528
rect 30854 61301 30906 61353
rect 31065 61301 31117 61353
rect 31276 61301 31328 61353
rect 31486 61350 31538 61353
rect 31697 61350 31749 61353
rect 31909 61350 31961 61353
rect 32120 61350 32172 61353
rect 32330 61350 32382 61353
rect 32541 61350 32593 61353
rect 32752 61350 32804 61353
rect 34284 61350 34336 61353
rect 34495 61350 34547 61353
rect 31486 61304 31538 61350
rect 31697 61304 31749 61350
rect 31909 61304 31961 61350
rect 32120 61304 32172 61350
rect 32330 61304 32382 61350
rect 32541 61304 32593 61350
rect 32752 61304 32804 61350
rect 34284 61304 34302 61350
rect 34302 61304 34336 61350
rect 34495 61304 34508 61350
rect 34508 61304 34547 61350
rect 31486 61301 31538 61304
rect 31697 61301 31749 61304
rect 31909 61301 31961 61304
rect 32120 61301 32172 61304
rect 32330 61301 32382 61304
rect 32541 61301 32593 61304
rect 32752 61301 32804 61304
rect 34284 61301 34336 61304
rect 34495 61301 34547 61304
rect 34707 61301 34759 61353
rect 34918 61301 34970 61353
rect 35220 61301 35272 61353
rect 35430 61301 35482 61353
rect 35641 61301 35693 61353
rect 35853 61301 35905 61353
rect 36064 61301 36116 61353
rect 36274 61301 36326 61353
rect 38330 61350 38382 61353
rect 38330 61304 38382 61350
rect 38330 61301 38382 61304
rect 38541 61301 38593 61353
rect 38752 61301 38804 61353
rect 39052 61350 39104 61353
rect 39232 61350 39284 61353
rect 39052 61304 39062 61350
rect 39062 61304 39104 61350
rect 39232 61304 39266 61350
rect 39266 61304 39284 61350
rect 39052 61301 39104 61304
rect 39232 61301 39284 61304
rect 33057 61126 33109 61129
rect 33237 61126 33289 61129
rect 33057 61080 33109 61126
rect 33237 61080 33289 61126
rect 33057 61077 33109 61080
rect 33237 61077 33289 61080
rect 33819 61126 33871 61137
rect 33999 61126 34051 61137
rect 33819 61085 33833 61126
rect 33833 61085 33871 61126
rect 33999 61085 34039 61126
rect 34039 61085 34051 61126
rect 35332 61039 35384 61051
rect 35543 61039 35595 61051
rect 35754 61039 35806 61051
rect 35965 61039 36017 61051
rect 36176 61039 36228 61051
rect 37891 61039 37943 61063
rect 38071 61039 38123 61063
rect 35332 60999 35384 61039
rect 35543 60999 35580 61039
rect 35580 60999 35595 61039
rect 35754 60999 35786 61039
rect 35786 60999 35806 61039
rect 35965 60999 35992 61039
rect 35992 60999 36017 61039
rect 36176 60999 36198 61039
rect 36198 60999 36228 61039
rect 37891 61011 37909 61039
rect 37909 61011 37943 61039
rect 38071 61011 38072 61039
rect 38072 61011 38123 61039
rect 34267 60856 34302 60891
rect 34302 60856 34319 60891
rect 34447 60856 34451 60891
rect 34451 60856 34499 60891
rect 34627 60856 34658 60891
rect 34658 60856 34679 60891
rect 34267 60839 34319 60856
rect 34447 60839 34499 60856
rect 34627 60839 34679 60856
rect 33057 60678 33109 60681
rect 33237 60678 33289 60681
rect 33057 60632 33109 60678
rect 33237 60632 33289 60678
rect 33057 60629 33109 60632
rect 33237 60629 33289 60632
rect 36678 60764 36697 60816
rect 36697 60764 36730 60816
rect 36961 60815 37013 60823
rect 37172 60815 37224 60823
rect 36961 60771 36971 60815
rect 36971 60771 37013 60815
rect 37172 60771 37206 60815
rect 37206 60771 37224 60815
rect 37384 60771 37436 60823
rect 37595 60771 37647 60823
rect 39994 61754 40046 61806
rect 39775 61574 39827 61591
rect 39775 61539 39786 61574
rect 39786 61539 39827 61574
rect 42312 61770 42364 61822
rect 41935 61539 41987 61591
rect 46731 61879 46783 61931
rect 48596 61925 48648 61977
rect 51835 62022 51887 62047
rect 52015 62022 52067 62047
rect 51835 61995 51887 62022
rect 52015 61995 52067 62022
rect 44939 61798 44991 61815
rect 45151 61798 45203 61815
rect 44939 61763 44971 61798
rect 44971 61763 44991 61798
rect 45151 61763 45197 61798
rect 45197 61763 45203 61798
rect 48596 61707 48648 61759
rect 50300 61763 50352 61815
rect 50511 61798 50563 61815
rect 50511 61763 50513 61798
rect 50513 61763 50563 61798
rect 50722 61763 50774 61815
rect 48943 61615 48984 61652
rect 48984 61615 48995 61652
rect 49154 61615 49190 61652
rect 49190 61615 49206 61652
rect 49365 61615 49396 61652
rect 49396 61615 49417 61652
rect 49576 61615 49602 61652
rect 49602 61615 49628 61652
rect 49787 61615 49839 61652
rect 48943 61600 48995 61615
rect 49154 61600 49206 61615
rect 49365 61600 49417 61615
rect 49576 61600 49628 61615
rect 49787 61600 49839 61615
rect 51073 61574 51125 61577
rect 51253 61574 51305 61577
rect 51073 61528 51086 61574
rect 51086 61528 51125 61574
rect 51253 61528 51292 61574
rect 51292 61528 51305 61574
rect 51073 61525 51125 61528
rect 51253 61525 51305 61528
rect 51835 61574 51887 61584
rect 52015 61574 52067 61584
rect 51835 61532 51887 61574
rect 52015 61532 52067 61574
rect 40253 61301 40305 61353
rect 40433 61301 40485 61353
rect 43790 61301 43842 61353
rect 44001 61301 44053 61353
rect 44213 61350 44265 61353
rect 44213 61304 44236 61350
rect 44236 61304 44265 61350
rect 44213 61301 44265 61304
rect 44424 61301 44476 61353
rect 44834 61350 44886 61353
rect 45045 61350 45097 61353
rect 45256 61350 45308 61353
rect 44834 61304 44858 61350
rect 44858 61304 44886 61350
rect 45045 61304 45084 61350
rect 45084 61304 45097 61350
rect 45256 61304 45264 61350
rect 45264 61304 45308 61350
rect 44834 61301 44886 61304
rect 45045 61301 45097 61304
rect 45256 61301 45308 61304
rect 48838 61301 48890 61353
rect 49048 61301 49100 61353
rect 49259 61301 49311 61353
rect 49471 61301 49523 61353
rect 49682 61301 49734 61353
rect 49892 61301 49944 61353
rect 50346 61301 50398 61353
rect 50557 61350 50609 61353
rect 50768 61350 50820 61353
rect 52316 61350 52368 61353
rect 52527 61350 52579 61353
rect 52738 61350 52790 61353
rect 52948 61350 53000 61353
rect 53159 61350 53211 61353
rect 53371 61350 53423 61353
rect 53582 61350 53634 61353
rect 50557 61304 50571 61350
rect 50571 61304 50609 61350
rect 50768 61304 50777 61350
rect 50777 61304 50820 61350
rect 52316 61304 52368 61350
rect 52527 61304 52579 61350
rect 52738 61304 52790 61350
rect 52948 61304 53000 61350
rect 53159 61304 53211 61350
rect 53371 61304 53423 61350
rect 53582 61304 53634 61350
rect 50557 61301 50609 61304
rect 50768 61301 50820 61304
rect 39775 61080 39786 61115
rect 39786 61080 39827 61115
rect 39775 61063 39827 61080
rect 39994 60848 40046 60900
rect 39994 60662 40046 60714
rect 52316 61301 52368 61304
rect 52527 61301 52579 61304
rect 52738 61301 52790 61304
rect 52948 61301 53000 61304
rect 53159 61301 53211 61304
rect 53371 61301 53423 61304
rect 53582 61301 53634 61304
rect 53792 61301 53844 61353
rect 54003 61301 54055 61353
rect 54214 61301 54266 61353
rect 54855 61301 54907 61353
rect 55066 61301 55118 61353
rect 55278 61350 55330 61353
rect 55278 61304 55279 61350
rect 55279 61304 55325 61350
rect 55325 61304 55330 61350
rect 55278 61301 55330 61304
rect 55489 61301 55541 61353
rect 41935 61063 41987 61115
rect 51073 61126 51125 61129
rect 51253 61126 51305 61129
rect 42312 60832 42364 60884
rect 51073 61080 51086 61126
rect 51086 61080 51125 61126
rect 51253 61080 51292 61126
rect 51292 61080 51305 61126
rect 48943 61039 48995 61054
rect 49154 61039 49206 61054
rect 49365 61039 49417 61054
rect 49576 61039 49628 61054
rect 49787 61039 49839 61054
rect 48943 61002 48984 61039
rect 48984 61002 48995 61039
rect 49154 61002 49190 61039
rect 49190 61002 49206 61039
rect 49365 61002 49396 61039
rect 49396 61002 49417 61039
rect 49576 61002 49602 61039
rect 49602 61002 49628 61039
rect 49787 61002 49839 61039
rect 51073 61077 51125 61080
rect 51253 61077 51305 61080
rect 44939 60856 44971 60891
rect 44971 60856 44991 60891
rect 45151 60856 45197 60891
rect 45197 60856 45203 60891
rect 48596 60895 48648 60947
rect 44939 60839 44991 60856
rect 45151 60839 45203 60856
rect 47108 60723 47160 60775
rect 50300 60839 50352 60891
rect 50511 60856 50513 60891
rect 50513 60856 50563 60891
rect 50511 60839 50563 60856
rect 50722 60839 50774 60891
rect 48596 60677 48648 60729
rect 51835 61080 51887 61122
rect 52015 61080 52067 61122
rect 51835 61070 51887 61080
rect 52015 61070 52067 61080
rect 35332 60545 35384 60591
rect 35543 60545 35580 60591
rect 35580 60545 35595 60591
rect 35754 60545 35786 60591
rect 35786 60545 35806 60591
rect 35965 60545 35992 60591
rect 35992 60545 36017 60591
rect 36176 60545 36198 60591
rect 36198 60545 36228 60591
rect 37891 60545 37909 60589
rect 37909 60545 37943 60589
rect 38071 60545 38072 60589
rect 38072 60545 38123 60589
rect 48943 60545 48984 60591
rect 48984 60545 48995 60591
rect 49154 60545 49190 60591
rect 49190 60545 49206 60591
rect 49365 60545 49396 60591
rect 49396 60545 49417 60591
rect 49576 60545 49602 60591
rect 49602 60545 49628 60591
rect 49787 60545 49839 60591
rect 51835 60632 51887 60659
rect 52015 60632 52067 60659
rect 51835 60607 51887 60632
rect 52015 60607 52067 60632
rect 35332 60539 35384 60545
rect 35543 60539 35595 60545
rect 35754 60539 35806 60545
rect 35965 60539 36017 60545
rect 36176 60539 36228 60545
rect 37891 60537 37943 60545
rect 38071 60537 38123 60545
rect 27790 60401 27842 60453
rect 28001 60401 28053 60453
rect 28212 60401 28264 60453
rect 28423 60401 28475 60453
rect 28634 60401 28686 60453
rect 28845 60450 28897 60453
rect 28845 60404 28856 60450
rect 28856 60404 28897 60450
rect 28845 60401 28897 60404
rect 29056 60401 29108 60453
rect 29582 60401 29634 60453
rect 29793 60450 29845 60453
rect 29793 60404 29798 60450
rect 29798 60404 29844 60450
rect 29844 60404 29845 60450
rect 29793 60401 29845 60404
rect 30005 60401 30057 60453
rect 30216 60401 30268 60453
rect 30854 60401 30906 60453
rect 31065 60401 31117 60453
rect 31276 60401 31328 60453
rect 31486 60401 31538 60453
rect 31697 60401 31749 60453
rect 31909 60401 31961 60453
rect 32120 60401 32172 60453
rect 32330 60401 32382 60453
rect 32541 60401 32593 60453
rect 32752 60401 32804 60453
rect 48943 60539 48995 60545
rect 49154 60539 49206 60545
rect 49365 60539 49417 60545
rect 49576 60539 49628 60545
rect 49787 60539 49839 60545
rect 34755 60401 34807 60453
rect 34935 60450 34987 60453
rect 34935 60404 34962 60450
rect 34962 60404 34987 60450
rect 34935 60401 34987 60404
rect 50138 60450 50190 60453
rect 50138 60404 50160 60450
rect 50160 60404 50190 60450
rect 50138 60401 50190 60404
rect 50318 60401 50370 60453
rect 35332 60309 35384 60315
rect 35543 60309 35595 60315
rect 35754 60309 35806 60315
rect 35965 60309 36017 60315
rect 36176 60309 36228 60315
rect 37891 60309 37943 60317
rect 38071 60309 38123 60317
rect 52316 60401 52368 60453
rect 52527 60401 52579 60453
rect 52738 60401 52790 60453
rect 52948 60401 53000 60453
rect 53159 60401 53211 60453
rect 53371 60401 53423 60453
rect 53582 60401 53634 60453
rect 53792 60401 53844 60453
rect 54003 60401 54055 60453
rect 54214 60401 54266 60453
rect 54855 60401 54907 60453
rect 55066 60401 55118 60453
rect 55278 60450 55330 60453
rect 55278 60404 55279 60450
rect 55279 60404 55325 60450
rect 55325 60404 55330 60450
rect 55278 60401 55330 60404
rect 55489 60401 55541 60453
rect 56015 60401 56067 60453
rect 56226 60450 56278 60453
rect 56226 60404 56267 60450
rect 56267 60404 56278 60450
rect 56226 60401 56278 60404
rect 56437 60401 56489 60453
rect 56648 60401 56700 60453
rect 56859 60401 56911 60453
rect 57070 60401 57122 60453
rect 57281 60401 57333 60453
rect 48943 60309 48995 60315
rect 49154 60309 49206 60315
rect 49365 60309 49417 60315
rect 49576 60309 49628 60315
rect 49787 60309 49839 60315
rect 33057 60222 33109 60225
rect 33237 60222 33289 60225
rect 35332 60263 35384 60309
rect 35543 60263 35580 60309
rect 35580 60263 35595 60309
rect 35754 60263 35786 60309
rect 35786 60263 35806 60309
rect 35965 60263 35992 60309
rect 35992 60263 36017 60309
rect 36176 60263 36198 60309
rect 36198 60263 36228 60309
rect 37891 60265 37909 60309
rect 37909 60265 37943 60309
rect 38071 60265 38072 60309
rect 38072 60265 38123 60309
rect 33057 60176 33109 60222
rect 33237 60176 33289 60222
rect 33057 60173 33109 60176
rect 33237 60173 33289 60176
rect 33057 59774 33109 59777
rect 33237 59774 33289 59777
rect 33057 59728 33109 59774
rect 33237 59728 33289 59774
rect 33057 59725 33109 59728
rect 33237 59725 33289 59728
rect 29582 59501 29634 59553
rect 29793 59550 29845 59553
rect 29793 59504 29798 59550
rect 29798 59504 29844 59550
rect 29844 59504 29845 59550
rect 29793 59501 29845 59504
rect 30005 59501 30057 59553
rect 30216 59501 30268 59553
rect 34267 59998 34319 60015
rect 34447 59998 34499 60015
rect 34627 59998 34679 60015
rect 34267 59963 34302 59998
rect 34302 59963 34319 59998
rect 34447 59963 34451 59998
rect 34451 59963 34499 59998
rect 34627 59963 34658 59998
rect 34658 59963 34679 59998
rect 36678 60038 36697 60090
rect 36697 60038 36730 60090
rect 48943 60263 48984 60309
rect 48984 60263 48995 60309
rect 49154 60263 49190 60309
rect 49190 60263 49206 60309
rect 49365 60263 49396 60309
rect 49396 60263 49417 60309
rect 49576 60263 49602 60309
rect 49602 60263 49628 60309
rect 49787 60263 49839 60309
rect 39994 60140 40046 60192
rect 36961 60039 36971 60083
rect 36971 60039 37013 60083
rect 37172 60039 37206 60083
rect 37206 60039 37224 60083
rect 36961 60031 37013 60039
rect 37172 60031 37224 60039
rect 37384 60031 37436 60083
rect 37595 60031 37647 60083
rect 35332 59815 35384 59855
rect 35543 59815 35580 59855
rect 35580 59815 35595 59855
rect 35754 59815 35786 59855
rect 35786 59815 35806 59855
rect 35965 59815 35992 59855
rect 35992 59815 36017 59855
rect 36176 59815 36198 59855
rect 36198 59815 36228 59855
rect 37891 59815 37909 59843
rect 37909 59815 37943 59843
rect 38071 59815 38072 59843
rect 38072 59815 38123 59843
rect 35332 59803 35384 59815
rect 35543 59803 35595 59815
rect 35754 59803 35806 59815
rect 35965 59803 36017 59815
rect 36176 59803 36228 59815
rect 33819 59728 33833 59769
rect 33833 59728 33871 59769
rect 33999 59728 34039 59769
rect 34039 59728 34051 59769
rect 37891 59791 37943 59815
rect 38071 59791 38123 59815
rect 33819 59717 33871 59728
rect 33999 59717 34051 59728
rect 30854 59501 30906 59553
rect 31065 59501 31117 59553
rect 31276 59501 31328 59553
rect 31486 59550 31538 59553
rect 31697 59550 31749 59553
rect 31909 59550 31961 59553
rect 32120 59550 32172 59553
rect 32330 59550 32382 59553
rect 32541 59550 32593 59553
rect 32752 59550 32804 59553
rect 34284 59550 34336 59553
rect 34495 59550 34547 59553
rect 31486 59504 31538 59550
rect 31697 59504 31749 59550
rect 31909 59504 31961 59550
rect 32120 59504 32172 59550
rect 32330 59504 32382 59550
rect 32541 59504 32593 59550
rect 32752 59504 32804 59550
rect 34284 59504 34302 59550
rect 34302 59504 34336 59550
rect 34495 59504 34508 59550
rect 34508 59504 34547 59550
rect 31486 59501 31538 59504
rect 31697 59501 31749 59504
rect 31909 59501 31961 59504
rect 32120 59501 32172 59504
rect 32330 59501 32382 59504
rect 32541 59501 32593 59504
rect 32752 59501 32804 59504
rect 34284 59501 34336 59504
rect 34495 59501 34547 59504
rect 34707 59501 34759 59553
rect 34918 59501 34970 59553
rect 35220 59501 35272 59553
rect 35430 59501 35482 59553
rect 35641 59501 35693 59553
rect 35853 59501 35905 59553
rect 36064 59501 36116 59553
rect 36274 59501 36326 59553
rect 38330 59550 38382 59553
rect 38330 59504 38382 59550
rect 38330 59501 38382 59504
rect 38541 59501 38593 59553
rect 38752 59501 38804 59553
rect 39052 59550 39104 59553
rect 39232 59550 39284 59553
rect 39052 59504 39062 59550
rect 39062 59504 39104 59550
rect 39232 59504 39266 59550
rect 39266 59504 39284 59550
rect 39052 59501 39104 59504
rect 39232 59501 39284 59504
rect 33057 59326 33109 59329
rect 33237 59326 33289 59329
rect 33057 59280 33109 59326
rect 33237 59280 33289 59326
rect 33057 59277 33109 59280
rect 33237 59277 33289 59280
rect 33819 59326 33871 59337
rect 33999 59326 34051 59337
rect 33819 59285 33833 59326
rect 33833 59285 33871 59326
rect 33999 59285 34039 59326
rect 34039 59285 34051 59326
rect 35332 59239 35384 59251
rect 35543 59239 35595 59251
rect 35754 59239 35806 59251
rect 35965 59239 36017 59251
rect 36176 59239 36228 59251
rect 37891 59239 37943 59263
rect 38071 59239 38123 59263
rect 35332 59199 35384 59239
rect 35543 59199 35580 59239
rect 35580 59199 35595 59239
rect 35754 59199 35786 59239
rect 35786 59199 35806 59239
rect 35965 59199 35992 59239
rect 35992 59199 36017 59239
rect 36176 59199 36198 59239
rect 36198 59199 36228 59239
rect 37891 59211 37909 59239
rect 37909 59211 37943 59239
rect 38071 59211 38072 59239
rect 38072 59211 38123 59239
rect 34267 59056 34302 59091
rect 34302 59056 34319 59091
rect 34447 59056 34451 59091
rect 34451 59056 34499 59091
rect 34627 59056 34658 59091
rect 34658 59056 34679 59091
rect 34267 59039 34319 59056
rect 34447 59039 34499 59056
rect 34627 59039 34679 59056
rect 33057 58878 33109 58881
rect 33237 58878 33289 58881
rect 33057 58832 33109 58878
rect 33237 58832 33289 58878
rect 33057 58829 33109 58832
rect 33237 58829 33289 58832
rect 36678 58964 36697 59016
rect 36697 58964 36730 59016
rect 36961 59015 37013 59023
rect 37172 59015 37224 59023
rect 36961 58971 36971 59015
rect 36971 58971 37013 59015
rect 37172 58971 37206 59015
rect 37206 58971 37224 59015
rect 37384 58971 37436 59023
rect 37595 58971 37647 59023
rect 39994 59954 40046 60006
rect 39775 59774 39827 59791
rect 39775 59739 39786 59774
rect 39786 59739 39827 59774
rect 42312 59970 42364 60022
rect 41935 59739 41987 59791
rect 47486 60079 47538 60131
rect 48596 60125 48648 60177
rect 51835 60222 51887 60247
rect 52015 60222 52067 60247
rect 51835 60195 51887 60222
rect 52015 60195 52067 60222
rect 44939 59998 44991 60015
rect 45151 59998 45203 60015
rect 44939 59963 44971 59998
rect 44971 59963 44991 59998
rect 45151 59963 45197 59998
rect 45197 59963 45203 59998
rect 48596 59907 48648 59959
rect 50300 59963 50352 60015
rect 50511 59998 50563 60015
rect 50511 59963 50513 59998
rect 50513 59963 50563 59998
rect 50722 59963 50774 60015
rect 48943 59815 48984 59852
rect 48984 59815 48995 59852
rect 49154 59815 49190 59852
rect 49190 59815 49206 59852
rect 49365 59815 49396 59852
rect 49396 59815 49417 59852
rect 49576 59815 49602 59852
rect 49602 59815 49628 59852
rect 49787 59815 49839 59852
rect 48943 59800 48995 59815
rect 49154 59800 49206 59815
rect 49365 59800 49417 59815
rect 49576 59800 49628 59815
rect 49787 59800 49839 59815
rect 51073 59774 51125 59777
rect 51253 59774 51305 59777
rect 51073 59728 51086 59774
rect 51086 59728 51125 59774
rect 51253 59728 51292 59774
rect 51292 59728 51305 59774
rect 51073 59725 51125 59728
rect 51253 59725 51305 59728
rect 51835 59774 51887 59784
rect 52015 59774 52067 59784
rect 51835 59732 51887 59774
rect 52015 59732 52067 59774
rect 40253 59501 40305 59553
rect 40433 59501 40485 59553
rect 43790 59501 43842 59553
rect 44001 59501 44053 59553
rect 44213 59550 44265 59553
rect 44213 59504 44236 59550
rect 44236 59504 44265 59550
rect 44213 59501 44265 59504
rect 44424 59501 44476 59553
rect 44834 59550 44886 59553
rect 45045 59550 45097 59553
rect 45256 59550 45308 59553
rect 44834 59504 44858 59550
rect 44858 59504 44886 59550
rect 45045 59504 45084 59550
rect 45084 59504 45097 59550
rect 45256 59504 45264 59550
rect 45264 59504 45308 59550
rect 44834 59501 44886 59504
rect 45045 59501 45097 59504
rect 45256 59501 45308 59504
rect 48838 59501 48890 59553
rect 49048 59501 49100 59553
rect 49259 59501 49311 59553
rect 49471 59501 49523 59553
rect 49682 59501 49734 59553
rect 49892 59501 49944 59553
rect 50346 59501 50398 59553
rect 50557 59550 50609 59553
rect 50768 59550 50820 59553
rect 52316 59550 52368 59553
rect 52527 59550 52579 59553
rect 52738 59550 52790 59553
rect 52948 59550 53000 59553
rect 53159 59550 53211 59553
rect 53371 59550 53423 59553
rect 53582 59550 53634 59553
rect 50557 59504 50571 59550
rect 50571 59504 50609 59550
rect 50768 59504 50777 59550
rect 50777 59504 50820 59550
rect 52316 59504 52368 59550
rect 52527 59504 52579 59550
rect 52738 59504 52790 59550
rect 52948 59504 53000 59550
rect 53159 59504 53211 59550
rect 53371 59504 53423 59550
rect 53582 59504 53634 59550
rect 50557 59501 50609 59504
rect 50768 59501 50820 59504
rect 39775 59280 39786 59315
rect 39786 59280 39827 59315
rect 39775 59263 39827 59280
rect 39994 59048 40046 59100
rect 39994 58862 40046 58914
rect 52316 59501 52368 59504
rect 52527 59501 52579 59504
rect 52738 59501 52790 59504
rect 52948 59501 53000 59504
rect 53159 59501 53211 59504
rect 53371 59501 53423 59504
rect 53582 59501 53634 59504
rect 53792 59501 53844 59553
rect 54003 59501 54055 59553
rect 54214 59501 54266 59553
rect 54855 59501 54907 59553
rect 55066 59501 55118 59553
rect 55278 59550 55330 59553
rect 55278 59504 55279 59550
rect 55279 59504 55325 59550
rect 55325 59504 55330 59550
rect 55278 59501 55330 59504
rect 55489 59501 55541 59553
rect 41935 59263 41987 59315
rect 51073 59326 51125 59329
rect 51253 59326 51305 59329
rect 42312 59032 42364 59084
rect 51073 59280 51086 59326
rect 51086 59280 51125 59326
rect 51253 59280 51292 59326
rect 51292 59280 51305 59326
rect 48943 59239 48995 59254
rect 49154 59239 49206 59254
rect 49365 59239 49417 59254
rect 49576 59239 49628 59254
rect 49787 59239 49839 59254
rect 48943 59202 48984 59239
rect 48984 59202 48995 59239
rect 49154 59202 49190 59239
rect 49190 59202 49206 59239
rect 49365 59202 49396 59239
rect 49396 59202 49417 59239
rect 49576 59202 49602 59239
rect 49602 59202 49628 59239
rect 49787 59202 49839 59239
rect 51073 59277 51125 59280
rect 51253 59277 51305 59280
rect 44939 59056 44971 59091
rect 44971 59056 44991 59091
rect 45151 59056 45197 59091
rect 45197 59056 45203 59091
rect 48596 59095 48648 59147
rect 44939 59039 44991 59056
rect 45151 59039 45203 59056
rect 47864 58923 47916 58975
rect 50300 59039 50352 59091
rect 50511 59056 50513 59091
rect 50513 59056 50563 59091
rect 50511 59039 50563 59056
rect 50722 59039 50774 59091
rect 48596 58877 48648 58929
rect 51835 59280 51887 59322
rect 52015 59280 52067 59322
rect 51835 59270 51887 59280
rect 52015 59270 52067 59280
rect 35332 58745 35384 58791
rect 35543 58745 35580 58791
rect 35580 58745 35595 58791
rect 35754 58745 35786 58791
rect 35786 58745 35806 58791
rect 35965 58745 35992 58791
rect 35992 58745 36017 58791
rect 36176 58745 36198 58791
rect 36198 58745 36228 58791
rect 37891 58745 37909 58789
rect 37909 58745 37943 58789
rect 38071 58745 38072 58789
rect 38072 58745 38123 58789
rect 48943 58745 48984 58791
rect 48984 58745 48995 58791
rect 49154 58745 49190 58791
rect 49190 58745 49206 58791
rect 49365 58745 49396 58791
rect 49396 58745 49417 58791
rect 49576 58745 49602 58791
rect 49602 58745 49628 58791
rect 49787 58745 49839 58791
rect 51835 58832 51887 58859
rect 52015 58832 52067 58859
rect 51835 58807 51887 58832
rect 52015 58807 52067 58832
rect 35332 58739 35384 58745
rect 35543 58739 35595 58745
rect 35754 58739 35806 58745
rect 35965 58739 36017 58745
rect 36176 58739 36228 58745
rect 37891 58737 37943 58745
rect 38071 58737 38123 58745
rect 27790 58601 27842 58653
rect 28001 58601 28053 58653
rect 28212 58601 28264 58653
rect 28423 58601 28475 58653
rect 28634 58601 28686 58653
rect 28845 58650 28897 58653
rect 28845 58604 28856 58650
rect 28856 58604 28897 58650
rect 28845 58601 28897 58604
rect 29056 58601 29108 58653
rect 29582 58601 29634 58653
rect 29793 58650 29845 58653
rect 29793 58604 29798 58650
rect 29798 58604 29844 58650
rect 29844 58604 29845 58650
rect 29793 58601 29845 58604
rect 30005 58601 30057 58653
rect 30216 58601 30268 58653
rect 30854 58601 30906 58653
rect 31065 58601 31117 58653
rect 31276 58601 31328 58653
rect 31486 58601 31538 58653
rect 31697 58601 31749 58653
rect 31909 58601 31961 58653
rect 32120 58601 32172 58653
rect 32330 58601 32382 58653
rect 32541 58601 32593 58653
rect 32752 58601 32804 58653
rect 48943 58739 48995 58745
rect 49154 58739 49206 58745
rect 49365 58739 49417 58745
rect 49576 58739 49628 58745
rect 49787 58739 49839 58745
rect 34755 58601 34807 58653
rect 34935 58650 34987 58653
rect 34935 58604 34962 58650
rect 34962 58604 34987 58650
rect 34935 58601 34987 58604
rect 50138 58650 50190 58653
rect 50138 58604 50160 58650
rect 50160 58604 50190 58650
rect 50138 58601 50190 58604
rect 50318 58601 50370 58653
rect 35332 58509 35384 58515
rect 35543 58509 35595 58515
rect 35754 58509 35806 58515
rect 35965 58509 36017 58515
rect 36176 58509 36228 58515
rect 37891 58509 37943 58517
rect 38071 58509 38123 58517
rect 52316 58601 52368 58653
rect 52527 58601 52579 58653
rect 52738 58601 52790 58653
rect 52948 58601 53000 58653
rect 53159 58601 53211 58653
rect 53371 58601 53423 58653
rect 53582 58601 53634 58653
rect 53792 58601 53844 58653
rect 54003 58601 54055 58653
rect 54214 58601 54266 58653
rect 54855 58601 54907 58653
rect 55066 58601 55118 58653
rect 55278 58650 55330 58653
rect 55278 58604 55279 58650
rect 55279 58604 55325 58650
rect 55325 58604 55330 58650
rect 55278 58601 55330 58604
rect 55489 58601 55541 58653
rect 56015 58601 56067 58653
rect 56226 58650 56278 58653
rect 56226 58604 56267 58650
rect 56267 58604 56278 58650
rect 56226 58601 56278 58604
rect 56437 58601 56489 58653
rect 56648 58601 56700 58653
rect 56859 58601 56911 58653
rect 57070 58601 57122 58653
rect 57281 58601 57333 58653
rect 48943 58509 48995 58515
rect 49154 58509 49206 58515
rect 49365 58509 49417 58515
rect 49576 58509 49628 58515
rect 49787 58509 49839 58515
rect 33057 58422 33109 58425
rect 33237 58422 33289 58425
rect 35332 58463 35384 58509
rect 35543 58463 35580 58509
rect 35580 58463 35595 58509
rect 35754 58463 35786 58509
rect 35786 58463 35806 58509
rect 35965 58463 35992 58509
rect 35992 58463 36017 58509
rect 36176 58463 36198 58509
rect 36198 58463 36228 58509
rect 37891 58465 37909 58509
rect 37909 58465 37943 58509
rect 38071 58465 38072 58509
rect 38072 58465 38123 58509
rect 33057 58376 33109 58422
rect 33237 58376 33289 58422
rect 33057 58373 33109 58376
rect 33237 58373 33289 58376
rect 33057 57974 33109 57977
rect 33237 57974 33289 57977
rect 33057 57928 33109 57974
rect 33237 57928 33289 57974
rect 33057 57925 33109 57928
rect 33237 57925 33289 57928
rect 29582 57701 29634 57753
rect 29793 57750 29845 57753
rect 29793 57704 29798 57750
rect 29798 57704 29844 57750
rect 29844 57704 29845 57750
rect 29793 57701 29845 57704
rect 30005 57701 30057 57753
rect 30216 57701 30268 57753
rect 34267 58198 34319 58215
rect 34447 58198 34499 58215
rect 34627 58198 34679 58215
rect 34267 58163 34302 58198
rect 34302 58163 34319 58198
rect 34447 58163 34451 58198
rect 34451 58163 34499 58198
rect 34627 58163 34658 58198
rect 34658 58163 34679 58198
rect 36678 58238 36697 58290
rect 36697 58238 36730 58290
rect 48943 58463 48984 58509
rect 48984 58463 48995 58509
rect 49154 58463 49190 58509
rect 49190 58463 49206 58509
rect 49365 58463 49396 58509
rect 49396 58463 49417 58509
rect 49576 58463 49602 58509
rect 49602 58463 49628 58509
rect 49787 58463 49839 58509
rect 39994 58340 40046 58392
rect 36961 58239 36971 58283
rect 36971 58239 37013 58283
rect 37172 58239 37206 58283
rect 37206 58239 37224 58283
rect 36961 58231 37013 58239
rect 37172 58231 37224 58239
rect 37384 58231 37436 58283
rect 37595 58231 37647 58283
rect 35332 58015 35384 58055
rect 35543 58015 35580 58055
rect 35580 58015 35595 58055
rect 35754 58015 35786 58055
rect 35786 58015 35806 58055
rect 35965 58015 35992 58055
rect 35992 58015 36017 58055
rect 36176 58015 36198 58055
rect 36198 58015 36228 58055
rect 37891 58015 37909 58043
rect 37909 58015 37943 58043
rect 38071 58015 38072 58043
rect 38072 58015 38123 58043
rect 35332 58003 35384 58015
rect 35543 58003 35595 58015
rect 35754 58003 35806 58015
rect 35965 58003 36017 58015
rect 36176 58003 36228 58015
rect 33819 57928 33833 57969
rect 33833 57928 33871 57969
rect 33999 57928 34039 57969
rect 34039 57928 34051 57969
rect 37891 57991 37943 58015
rect 38071 57991 38123 58015
rect 33819 57917 33871 57928
rect 33999 57917 34051 57928
rect 30854 57701 30906 57753
rect 31065 57701 31117 57753
rect 31276 57701 31328 57753
rect 31486 57750 31538 57753
rect 31697 57750 31749 57753
rect 31909 57750 31961 57753
rect 32120 57750 32172 57753
rect 32330 57750 32382 57753
rect 32541 57750 32593 57753
rect 32752 57750 32804 57753
rect 34284 57750 34336 57753
rect 34495 57750 34547 57753
rect 31486 57704 31538 57750
rect 31697 57704 31749 57750
rect 31909 57704 31961 57750
rect 32120 57704 32172 57750
rect 32330 57704 32382 57750
rect 32541 57704 32593 57750
rect 32752 57704 32804 57750
rect 34284 57704 34302 57750
rect 34302 57704 34336 57750
rect 34495 57704 34508 57750
rect 34508 57704 34547 57750
rect 31486 57701 31538 57704
rect 31697 57701 31749 57704
rect 31909 57701 31961 57704
rect 32120 57701 32172 57704
rect 32330 57701 32382 57704
rect 32541 57701 32593 57704
rect 32752 57701 32804 57704
rect 34284 57701 34336 57704
rect 34495 57701 34547 57704
rect 34707 57701 34759 57753
rect 34918 57701 34970 57753
rect 35220 57701 35272 57753
rect 35430 57701 35482 57753
rect 35641 57701 35693 57753
rect 35853 57701 35905 57753
rect 36064 57701 36116 57753
rect 36274 57701 36326 57753
rect 38330 57750 38382 57753
rect 38330 57704 38382 57750
rect 38330 57701 38382 57704
rect 38541 57701 38593 57753
rect 38752 57701 38804 57753
rect 39052 57750 39104 57753
rect 39232 57750 39284 57753
rect 39052 57704 39062 57750
rect 39062 57704 39104 57750
rect 39232 57704 39266 57750
rect 39266 57704 39284 57750
rect 39052 57701 39104 57704
rect 39232 57701 39284 57704
rect 33057 57526 33109 57529
rect 33237 57526 33289 57529
rect 33057 57480 33109 57526
rect 33237 57480 33289 57526
rect 33057 57477 33109 57480
rect 33237 57477 33289 57480
rect 33819 57526 33871 57537
rect 33999 57526 34051 57537
rect 33819 57485 33833 57526
rect 33833 57485 33871 57526
rect 33999 57485 34039 57526
rect 34039 57485 34051 57526
rect 35332 57439 35384 57451
rect 35543 57439 35595 57451
rect 35754 57439 35806 57451
rect 35965 57439 36017 57451
rect 36176 57439 36228 57451
rect 37891 57439 37943 57463
rect 38071 57439 38123 57463
rect 35332 57399 35384 57439
rect 35543 57399 35580 57439
rect 35580 57399 35595 57439
rect 35754 57399 35786 57439
rect 35786 57399 35806 57439
rect 35965 57399 35992 57439
rect 35992 57399 36017 57439
rect 36176 57399 36198 57439
rect 36198 57399 36228 57439
rect 37891 57411 37909 57439
rect 37909 57411 37943 57439
rect 38071 57411 38072 57439
rect 38072 57411 38123 57439
rect 34267 57256 34302 57291
rect 34302 57256 34319 57291
rect 34447 57256 34451 57291
rect 34451 57256 34499 57291
rect 34627 57256 34658 57291
rect 34658 57256 34679 57291
rect 34267 57239 34319 57256
rect 34447 57239 34499 57256
rect 34627 57239 34679 57256
rect 33057 57078 33109 57081
rect 33237 57078 33289 57081
rect 33057 57032 33109 57078
rect 33237 57032 33289 57078
rect 33057 57029 33109 57032
rect 33237 57029 33289 57032
rect 36678 57164 36697 57216
rect 36697 57164 36730 57216
rect 36961 57215 37013 57223
rect 37172 57215 37224 57223
rect 36961 57171 36971 57215
rect 36971 57171 37013 57215
rect 37172 57171 37206 57215
rect 37206 57171 37224 57215
rect 37384 57171 37436 57223
rect 37595 57171 37647 57223
rect 39994 58154 40046 58206
rect 39775 57974 39827 57991
rect 39775 57939 39786 57974
rect 39786 57939 39827 57974
rect 42312 58170 42364 58222
rect 41935 57939 41987 57991
rect 48241 58279 48293 58331
rect 48596 58325 48648 58377
rect 51835 58422 51887 58447
rect 52015 58422 52067 58447
rect 51835 58395 51887 58422
rect 52015 58395 52067 58422
rect 44939 58198 44991 58215
rect 45151 58198 45203 58215
rect 44939 58163 44971 58198
rect 44971 58163 44991 58198
rect 45151 58163 45197 58198
rect 45197 58163 45203 58198
rect 48596 58107 48648 58159
rect 50300 58163 50352 58215
rect 50511 58198 50563 58215
rect 50511 58163 50513 58198
rect 50513 58163 50563 58198
rect 50722 58163 50774 58215
rect 48943 58015 48984 58052
rect 48984 58015 48995 58052
rect 49154 58015 49190 58052
rect 49190 58015 49206 58052
rect 49365 58015 49396 58052
rect 49396 58015 49417 58052
rect 49576 58015 49602 58052
rect 49602 58015 49628 58052
rect 49787 58015 49839 58052
rect 48943 58000 48995 58015
rect 49154 58000 49206 58015
rect 49365 58000 49417 58015
rect 49576 58000 49628 58015
rect 49787 58000 49839 58015
rect 51073 57974 51125 57977
rect 51253 57974 51305 57977
rect 51073 57928 51086 57974
rect 51086 57928 51125 57974
rect 51253 57928 51292 57974
rect 51292 57928 51305 57974
rect 51073 57925 51125 57928
rect 51253 57925 51305 57928
rect 51835 57974 51887 57984
rect 52015 57974 52067 57984
rect 51835 57932 51887 57974
rect 52015 57932 52067 57974
rect 40253 57701 40305 57753
rect 40433 57701 40485 57753
rect 43790 57701 43842 57753
rect 44001 57701 44053 57753
rect 44213 57750 44265 57753
rect 44213 57704 44236 57750
rect 44236 57704 44265 57750
rect 44213 57701 44265 57704
rect 44424 57701 44476 57753
rect 44834 57750 44886 57753
rect 45045 57750 45097 57753
rect 45256 57750 45308 57753
rect 44834 57704 44858 57750
rect 44858 57704 44886 57750
rect 45045 57704 45084 57750
rect 45084 57704 45097 57750
rect 45256 57704 45264 57750
rect 45264 57704 45308 57750
rect 44834 57701 44886 57704
rect 45045 57701 45097 57704
rect 45256 57701 45308 57704
rect 48838 57701 48890 57753
rect 49048 57701 49100 57753
rect 49259 57701 49311 57753
rect 49471 57701 49523 57753
rect 49682 57701 49734 57753
rect 49892 57701 49944 57753
rect 50346 57701 50398 57753
rect 50557 57750 50609 57753
rect 50768 57750 50820 57753
rect 52316 57750 52368 57753
rect 52527 57750 52579 57753
rect 52738 57750 52790 57753
rect 52948 57750 53000 57753
rect 53159 57750 53211 57753
rect 53371 57750 53423 57753
rect 53582 57750 53634 57753
rect 50557 57704 50571 57750
rect 50571 57704 50609 57750
rect 50768 57704 50777 57750
rect 50777 57704 50820 57750
rect 52316 57704 52368 57750
rect 52527 57704 52579 57750
rect 52738 57704 52790 57750
rect 52948 57704 53000 57750
rect 53159 57704 53211 57750
rect 53371 57704 53423 57750
rect 53582 57704 53634 57750
rect 50557 57701 50609 57704
rect 50768 57701 50820 57704
rect 39775 57480 39786 57515
rect 39786 57480 39827 57515
rect 39775 57463 39827 57480
rect 39994 57248 40046 57300
rect 39994 57062 40046 57114
rect 52316 57701 52368 57704
rect 52527 57701 52579 57704
rect 52738 57701 52790 57704
rect 52948 57701 53000 57704
rect 53159 57701 53211 57704
rect 53371 57701 53423 57704
rect 53582 57701 53634 57704
rect 53792 57701 53844 57753
rect 54003 57701 54055 57753
rect 54214 57701 54266 57753
rect 54855 57701 54907 57753
rect 55066 57701 55118 57753
rect 55278 57750 55330 57753
rect 55278 57704 55279 57750
rect 55279 57704 55325 57750
rect 55325 57704 55330 57750
rect 55278 57701 55330 57704
rect 55489 57701 55541 57753
rect 41935 57463 41987 57515
rect 51073 57526 51125 57529
rect 51253 57526 51305 57529
rect 42690 57232 42742 57284
rect 51073 57480 51086 57526
rect 51086 57480 51125 57526
rect 51253 57480 51292 57526
rect 51292 57480 51305 57526
rect 48943 57439 48995 57454
rect 49154 57439 49206 57454
rect 49365 57439 49417 57454
rect 49576 57439 49628 57454
rect 49787 57439 49839 57454
rect 48943 57402 48984 57439
rect 48984 57402 48995 57439
rect 49154 57402 49190 57439
rect 49190 57402 49206 57439
rect 49365 57402 49396 57439
rect 49396 57402 49417 57439
rect 49576 57402 49602 57439
rect 49602 57402 49628 57439
rect 49787 57402 49839 57439
rect 51073 57477 51125 57480
rect 51253 57477 51305 57480
rect 44939 57256 44971 57291
rect 44971 57256 44991 57291
rect 45151 57256 45197 57291
rect 45197 57256 45203 57291
rect 48596 57295 48648 57347
rect 44939 57239 44991 57256
rect 45151 57239 45203 57256
rect 45597 57137 45604 57175
rect 45604 57137 45649 57175
rect 45597 57123 45649 57137
rect 50300 57239 50352 57291
rect 50511 57256 50513 57291
rect 50513 57256 50563 57291
rect 50511 57239 50563 57256
rect 50722 57239 50774 57291
rect 48596 57077 48648 57129
rect 51835 57480 51887 57522
rect 52015 57480 52067 57522
rect 51835 57470 51887 57480
rect 52015 57470 52067 57480
rect 35332 56945 35384 56991
rect 35543 56945 35580 56991
rect 35580 56945 35595 56991
rect 35754 56945 35786 56991
rect 35786 56945 35806 56991
rect 35965 56945 35992 56991
rect 35992 56945 36017 56991
rect 36176 56945 36198 56991
rect 36198 56945 36228 56991
rect 37891 56945 37909 56989
rect 37909 56945 37943 56989
rect 38071 56945 38072 56989
rect 38072 56945 38123 56989
rect 48943 56945 48984 56991
rect 48984 56945 48995 56991
rect 49154 56945 49190 56991
rect 49190 56945 49206 56991
rect 49365 56945 49396 56991
rect 49396 56945 49417 56991
rect 49576 56945 49602 56991
rect 49602 56945 49628 56991
rect 49787 56945 49839 56991
rect 51835 57032 51887 57059
rect 52015 57032 52067 57059
rect 51835 57007 51887 57032
rect 52015 57007 52067 57032
rect 35332 56939 35384 56945
rect 35543 56939 35595 56945
rect 35754 56939 35806 56945
rect 35965 56939 36017 56945
rect 36176 56939 36228 56945
rect 37891 56937 37943 56945
rect 38071 56937 38123 56945
rect 27790 56801 27842 56853
rect 28001 56801 28053 56853
rect 28212 56801 28264 56853
rect 28423 56801 28475 56853
rect 28634 56801 28686 56853
rect 28845 56850 28897 56853
rect 28845 56804 28856 56850
rect 28856 56804 28897 56850
rect 28845 56801 28897 56804
rect 29056 56801 29108 56853
rect 29582 56801 29634 56853
rect 29793 56850 29845 56853
rect 29793 56804 29798 56850
rect 29798 56804 29844 56850
rect 29844 56804 29845 56850
rect 29793 56801 29845 56804
rect 30005 56801 30057 56853
rect 30216 56801 30268 56853
rect 30854 56801 30906 56853
rect 31065 56801 31117 56853
rect 31276 56801 31328 56853
rect 31486 56801 31538 56853
rect 31697 56801 31749 56853
rect 31909 56801 31961 56853
rect 32120 56801 32172 56853
rect 32330 56801 32382 56853
rect 32541 56801 32593 56853
rect 32752 56801 32804 56853
rect 48943 56939 48995 56945
rect 49154 56939 49206 56945
rect 49365 56939 49417 56945
rect 49576 56939 49628 56945
rect 49787 56939 49839 56945
rect 34755 56801 34807 56853
rect 34935 56850 34987 56853
rect 34935 56804 34962 56850
rect 34962 56804 34987 56850
rect 34935 56801 34987 56804
rect 50138 56850 50190 56853
rect 50138 56804 50160 56850
rect 50160 56804 50190 56850
rect 50138 56801 50190 56804
rect 50318 56801 50370 56853
rect 35332 56709 35384 56715
rect 35543 56709 35595 56715
rect 35754 56709 35806 56715
rect 35965 56709 36017 56715
rect 36176 56709 36228 56715
rect 37891 56709 37943 56717
rect 38071 56709 38123 56717
rect 52316 56801 52368 56853
rect 52527 56801 52579 56853
rect 52738 56801 52790 56853
rect 52948 56801 53000 56853
rect 53159 56801 53211 56853
rect 53371 56801 53423 56853
rect 53582 56801 53634 56853
rect 53792 56801 53844 56853
rect 54003 56801 54055 56853
rect 54214 56801 54266 56853
rect 54855 56801 54907 56853
rect 55066 56801 55118 56853
rect 55278 56850 55330 56853
rect 55278 56804 55279 56850
rect 55279 56804 55325 56850
rect 55325 56804 55330 56850
rect 55278 56801 55330 56804
rect 55489 56801 55541 56853
rect 56015 56801 56067 56853
rect 56226 56850 56278 56853
rect 56226 56804 56267 56850
rect 56267 56804 56278 56850
rect 56226 56801 56278 56804
rect 56437 56801 56489 56853
rect 56648 56801 56700 56853
rect 56859 56801 56911 56853
rect 57070 56801 57122 56853
rect 57281 56801 57333 56853
rect 48943 56709 48995 56715
rect 49154 56709 49206 56715
rect 49365 56709 49417 56715
rect 49576 56709 49628 56715
rect 49787 56709 49839 56715
rect 33057 56622 33109 56625
rect 33237 56622 33289 56625
rect 35332 56663 35384 56709
rect 35543 56663 35580 56709
rect 35580 56663 35595 56709
rect 35754 56663 35786 56709
rect 35786 56663 35806 56709
rect 35965 56663 35992 56709
rect 35992 56663 36017 56709
rect 36176 56663 36198 56709
rect 36198 56663 36228 56709
rect 37891 56665 37909 56709
rect 37909 56665 37943 56709
rect 38071 56665 38072 56709
rect 38072 56665 38123 56709
rect 33057 56576 33109 56622
rect 33237 56576 33289 56622
rect 33057 56573 33109 56576
rect 33237 56573 33289 56576
rect 33057 56174 33109 56177
rect 33237 56174 33289 56177
rect 33057 56128 33109 56174
rect 33237 56128 33289 56174
rect 33057 56125 33109 56128
rect 33237 56125 33289 56128
rect 29582 55901 29634 55953
rect 29793 55950 29845 55953
rect 29793 55904 29798 55950
rect 29798 55904 29844 55950
rect 29844 55904 29845 55950
rect 29793 55901 29845 55904
rect 30005 55901 30057 55953
rect 30216 55901 30268 55953
rect 34267 56398 34319 56415
rect 34447 56398 34499 56415
rect 34627 56398 34679 56415
rect 34267 56363 34302 56398
rect 34302 56363 34319 56398
rect 34447 56363 34451 56398
rect 34451 56363 34499 56398
rect 34627 56363 34658 56398
rect 34658 56363 34679 56398
rect 36678 56438 36697 56490
rect 36697 56438 36730 56490
rect 48943 56663 48984 56709
rect 48984 56663 48995 56709
rect 49154 56663 49190 56709
rect 49190 56663 49206 56709
rect 49365 56663 49396 56709
rect 49396 56663 49417 56709
rect 49576 56663 49602 56709
rect 49602 56663 49628 56709
rect 49787 56663 49839 56709
rect 39994 56540 40046 56592
rect 36961 56439 36971 56483
rect 36971 56439 37013 56483
rect 37172 56439 37206 56483
rect 37206 56439 37224 56483
rect 36961 56431 37013 56439
rect 37172 56431 37224 56439
rect 37384 56431 37436 56483
rect 37595 56431 37647 56483
rect 35332 56215 35384 56255
rect 35543 56215 35580 56255
rect 35580 56215 35595 56255
rect 35754 56215 35786 56255
rect 35786 56215 35806 56255
rect 35965 56215 35992 56255
rect 35992 56215 36017 56255
rect 36176 56215 36198 56255
rect 36198 56215 36228 56255
rect 37891 56215 37909 56243
rect 37909 56215 37943 56243
rect 38071 56215 38072 56243
rect 38072 56215 38123 56243
rect 35332 56203 35384 56215
rect 35543 56203 35595 56215
rect 35754 56203 35806 56215
rect 35965 56203 36017 56215
rect 36176 56203 36228 56215
rect 33819 56128 33833 56169
rect 33833 56128 33871 56169
rect 33999 56128 34039 56169
rect 34039 56128 34051 56169
rect 37891 56191 37943 56215
rect 38071 56191 38123 56215
rect 33819 56117 33871 56128
rect 33999 56117 34051 56128
rect 30854 55901 30906 55953
rect 31065 55901 31117 55953
rect 31276 55901 31328 55953
rect 31486 55950 31538 55953
rect 31697 55950 31749 55953
rect 31909 55950 31961 55953
rect 32120 55950 32172 55953
rect 32330 55950 32382 55953
rect 32541 55950 32593 55953
rect 32752 55950 32804 55953
rect 34284 55950 34336 55953
rect 34495 55950 34547 55953
rect 31486 55904 31538 55950
rect 31697 55904 31749 55950
rect 31909 55904 31961 55950
rect 32120 55904 32172 55950
rect 32330 55904 32382 55950
rect 32541 55904 32593 55950
rect 32752 55904 32804 55950
rect 34284 55904 34302 55950
rect 34302 55904 34336 55950
rect 34495 55904 34508 55950
rect 34508 55904 34547 55950
rect 31486 55901 31538 55904
rect 31697 55901 31749 55904
rect 31909 55901 31961 55904
rect 32120 55901 32172 55904
rect 32330 55901 32382 55904
rect 32541 55901 32593 55904
rect 32752 55901 32804 55904
rect 34284 55901 34336 55904
rect 34495 55901 34547 55904
rect 34707 55901 34759 55953
rect 34918 55901 34970 55953
rect 35220 55901 35272 55953
rect 35430 55901 35482 55953
rect 35641 55901 35693 55953
rect 35853 55901 35905 55953
rect 36064 55901 36116 55953
rect 36274 55901 36326 55953
rect 38330 55950 38382 55953
rect 38330 55904 38382 55950
rect 38330 55901 38382 55904
rect 38541 55901 38593 55953
rect 38752 55901 38804 55953
rect 39052 55950 39104 55953
rect 39232 55950 39284 55953
rect 39052 55904 39062 55950
rect 39062 55904 39104 55950
rect 39232 55904 39266 55950
rect 39266 55904 39284 55950
rect 39052 55901 39104 55904
rect 39232 55901 39284 55904
rect 33057 55726 33109 55729
rect 33237 55726 33289 55729
rect 33057 55680 33109 55726
rect 33237 55680 33289 55726
rect 33057 55677 33109 55680
rect 33237 55677 33289 55680
rect 33819 55726 33871 55737
rect 33999 55726 34051 55737
rect 33819 55685 33833 55726
rect 33833 55685 33871 55726
rect 33999 55685 34039 55726
rect 34039 55685 34051 55726
rect 35332 55639 35384 55651
rect 35543 55639 35595 55651
rect 35754 55639 35806 55651
rect 35965 55639 36017 55651
rect 36176 55639 36228 55651
rect 37891 55639 37943 55663
rect 38071 55639 38123 55663
rect 35332 55599 35384 55639
rect 35543 55599 35580 55639
rect 35580 55599 35595 55639
rect 35754 55599 35786 55639
rect 35786 55599 35806 55639
rect 35965 55599 35992 55639
rect 35992 55599 36017 55639
rect 36176 55599 36198 55639
rect 36198 55599 36228 55639
rect 37891 55611 37909 55639
rect 37909 55611 37943 55639
rect 38071 55611 38072 55639
rect 38072 55611 38123 55639
rect 34267 55456 34302 55491
rect 34302 55456 34319 55491
rect 34447 55456 34451 55491
rect 34451 55456 34499 55491
rect 34627 55456 34658 55491
rect 34658 55456 34679 55491
rect 34267 55439 34319 55456
rect 34447 55439 34499 55456
rect 34627 55439 34679 55456
rect 33057 55278 33109 55281
rect 33237 55278 33289 55281
rect 33057 55232 33109 55278
rect 33237 55232 33289 55278
rect 33057 55229 33109 55232
rect 33237 55229 33289 55232
rect 36678 55364 36697 55416
rect 36697 55364 36730 55416
rect 36961 55415 37013 55423
rect 37172 55415 37224 55423
rect 36961 55371 36971 55415
rect 36971 55371 37013 55415
rect 37172 55371 37206 55415
rect 37206 55371 37224 55415
rect 37384 55371 37436 55423
rect 37595 55371 37647 55423
rect 39994 56354 40046 56406
rect 39775 56174 39827 56191
rect 39775 56139 39786 56174
rect 39786 56139 39827 56174
rect 42690 56370 42742 56422
rect 41935 56139 41987 56191
rect 45975 56479 46027 56531
rect 48596 56525 48648 56577
rect 51835 56622 51887 56647
rect 52015 56622 52067 56647
rect 51835 56595 51887 56622
rect 52015 56595 52067 56622
rect 44939 56398 44991 56415
rect 45151 56398 45203 56415
rect 44939 56363 44971 56398
rect 44971 56363 44991 56398
rect 45151 56363 45197 56398
rect 45197 56363 45203 56398
rect 48596 56307 48648 56359
rect 50300 56363 50352 56415
rect 50511 56398 50563 56415
rect 50511 56363 50513 56398
rect 50513 56363 50563 56398
rect 50722 56363 50774 56415
rect 48943 56215 48984 56252
rect 48984 56215 48995 56252
rect 49154 56215 49190 56252
rect 49190 56215 49206 56252
rect 49365 56215 49396 56252
rect 49396 56215 49417 56252
rect 49576 56215 49602 56252
rect 49602 56215 49628 56252
rect 49787 56215 49839 56252
rect 48943 56200 48995 56215
rect 49154 56200 49206 56215
rect 49365 56200 49417 56215
rect 49576 56200 49628 56215
rect 49787 56200 49839 56215
rect 51073 56174 51125 56177
rect 51253 56174 51305 56177
rect 51073 56128 51086 56174
rect 51086 56128 51125 56174
rect 51253 56128 51292 56174
rect 51292 56128 51305 56174
rect 51073 56125 51125 56128
rect 51253 56125 51305 56128
rect 51835 56174 51887 56184
rect 52015 56174 52067 56184
rect 51835 56132 51887 56174
rect 52015 56132 52067 56174
rect 40253 55901 40305 55953
rect 40433 55901 40485 55953
rect 43790 55901 43842 55953
rect 44001 55901 44053 55953
rect 44213 55950 44265 55953
rect 44213 55904 44236 55950
rect 44236 55904 44265 55950
rect 44213 55901 44265 55904
rect 44424 55901 44476 55953
rect 44834 55950 44886 55953
rect 45045 55950 45097 55953
rect 45256 55950 45308 55953
rect 44834 55904 44858 55950
rect 44858 55904 44886 55950
rect 45045 55904 45084 55950
rect 45084 55904 45097 55950
rect 45256 55904 45264 55950
rect 45264 55904 45308 55950
rect 44834 55901 44886 55904
rect 45045 55901 45097 55904
rect 45256 55901 45308 55904
rect 48838 55901 48890 55953
rect 49048 55901 49100 55953
rect 49259 55901 49311 55953
rect 49471 55901 49523 55953
rect 49682 55901 49734 55953
rect 49892 55901 49944 55953
rect 50346 55901 50398 55953
rect 50557 55950 50609 55953
rect 50768 55950 50820 55953
rect 52316 55950 52368 55953
rect 52527 55950 52579 55953
rect 52738 55950 52790 55953
rect 52948 55950 53000 55953
rect 53159 55950 53211 55953
rect 53371 55950 53423 55953
rect 53582 55950 53634 55953
rect 50557 55904 50571 55950
rect 50571 55904 50609 55950
rect 50768 55904 50777 55950
rect 50777 55904 50820 55950
rect 52316 55904 52368 55950
rect 52527 55904 52579 55950
rect 52738 55904 52790 55950
rect 52948 55904 53000 55950
rect 53159 55904 53211 55950
rect 53371 55904 53423 55950
rect 53582 55904 53634 55950
rect 50557 55901 50609 55904
rect 50768 55901 50820 55904
rect 39775 55680 39786 55715
rect 39786 55680 39827 55715
rect 39775 55663 39827 55680
rect 39994 55448 40046 55500
rect 39994 55262 40046 55314
rect 52316 55901 52368 55904
rect 52527 55901 52579 55904
rect 52738 55901 52790 55904
rect 52948 55901 53000 55904
rect 53159 55901 53211 55904
rect 53371 55901 53423 55904
rect 53582 55901 53634 55904
rect 53792 55901 53844 55953
rect 54003 55901 54055 55953
rect 54214 55901 54266 55953
rect 54855 55901 54907 55953
rect 55066 55901 55118 55953
rect 55278 55950 55330 55953
rect 55278 55904 55279 55950
rect 55279 55904 55325 55950
rect 55325 55904 55330 55950
rect 55278 55901 55330 55904
rect 55489 55901 55541 55953
rect 41935 55663 41987 55715
rect 51073 55726 51125 55729
rect 51253 55726 51305 55729
rect 42690 55432 42742 55484
rect 51073 55680 51086 55726
rect 51086 55680 51125 55726
rect 51253 55680 51292 55726
rect 51292 55680 51305 55726
rect 48943 55639 48995 55654
rect 49154 55639 49206 55654
rect 49365 55639 49417 55654
rect 49576 55639 49628 55654
rect 49787 55639 49839 55654
rect 48943 55602 48984 55639
rect 48984 55602 48995 55639
rect 49154 55602 49190 55639
rect 49190 55602 49206 55639
rect 49365 55602 49396 55639
rect 49396 55602 49417 55639
rect 49576 55602 49602 55639
rect 49602 55602 49628 55639
rect 49787 55602 49839 55639
rect 51073 55677 51125 55680
rect 51253 55677 51305 55680
rect 44939 55456 44971 55491
rect 44971 55456 44991 55491
rect 45151 55456 45197 55491
rect 45197 55456 45203 55491
rect 48596 55495 48648 55547
rect 44939 55439 44991 55456
rect 45151 55439 45203 55456
rect 46353 55323 46405 55375
rect 50300 55439 50352 55491
rect 50511 55456 50513 55491
rect 50513 55456 50563 55491
rect 50511 55439 50563 55456
rect 50722 55439 50774 55491
rect 48596 55277 48648 55329
rect 51835 55680 51887 55722
rect 52015 55680 52067 55722
rect 51835 55670 51887 55680
rect 52015 55670 52067 55680
rect 35332 55145 35384 55191
rect 35543 55145 35580 55191
rect 35580 55145 35595 55191
rect 35754 55145 35786 55191
rect 35786 55145 35806 55191
rect 35965 55145 35992 55191
rect 35992 55145 36017 55191
rect 36176 55145 36198 55191
rect 36198 55145 36228 55191
rect 37891 55145 37909 55189
rect 37909 55145 37943 55189
rect 38071 55145 38072 55189
rect 38072 55145 38123 55189
rect 48943 55145 48984 55191
rect 48984 55145 48995 55191
rect 49154 55145 49190 55191
rect 49190 55145 49206 55191
rect 49365 55145 49396 55191
rect 49396 55145 49417 55191
rect 49576 55145 49602 55191
rect 49602 55145 49628 55191
rect 49787 55145 49839 55191
rect 51835 55232 51887 55259
rect 52015 55232 52067 55259
rect 51835 55207 51887 55232
rect 52015 55207 52067 55232
rect 35332 55139 35384 55145
rect 35543 55139 35595 55145
rect 35754 55139 35806 55145
rect 35965 55139 36017 55145
rect 36176 55139 36228 55145
rect 37891 55137 37943 55145
rect 38071 55137 38123 55145
rect 27790 55001 27842 55053
rect 28001 55001 28053 55053
rect 28212 55001 28264 55053
rect 28423 55001 28475 55053
rect 28634 55001 28686 55053
rect 28845 55050 28897 55053
rect 28845 55004 28856 55050
rect 28856 55004 28897 55050
rect 28845 55001 28897 55004
rect 29056 55001 29108 55053
rect 29582 55001 29634 55053
rect 29793 55050 29845 55053
rect 29793 55004 29798 55050
rect 29798 55004 29844 55050
rect 29844 55004 29845 55050
rect 29793 55001 29845 55004
rect 30005 55001 30057 55053
rect 30216 55001 30268 55053
rect 30854 55001 30906 55053
rect 31065 55001 31117 55053
rect 31276 55001 31328 55053
rect 31486 55001 31538 55053
rect 31697 55001 31749 55053
rect 31909 55001 31961 55053
rect 32120 55001 32172 55053
rect 32330 55001 32382 55053
rect 32541 55001 32593 55053
rect 32752 55001 32804 55053
rect 48943 55139 48995 55145
rect 49154 55139 49206 55145
rect 49365 55139 49417 55145
rect 49576 55139 49628 55145
rect 49787 55139 49839 55145
rect 34755 55001 34807 55053
rect 34935 55050 34987 55053
rect 34935 55004 34962 55050
rect 34962 55004 34987 55050
rect 34935 55001 34987 55004
rect 50138 55050 50190 55053
rect 50138 55004 50160 55050
rect 50160 55004 50190 55050
rect 50138 55001 50190 55004
rect 50318 55001 50370 55053
rect 35332 54909 35384 54915
rect 35543 54909 35595 54915
rect 35754 54909 35806 54915
rect 35965 54909 36017 54915
rect 36176 54909 36228 54915
rect 37891 54909 37943 54917
rect 38071 54909 38123 54917
rect 52316 55001 52368 55053
rect 52527 55001 52579 55053
rect 52738 55001 52790 55053
rect 52948 55001 53000 55053
rect 53159 55001 53211 55053
rect 53371 55001 53423 55053
rect 53582 55001 53634 55053
rect 53792 55001 53844 55053
rect 54003 55001 54055 55053
rect 54214 55001 54266 55053
rect 54855 55001 54907 55053
rect 55066 55001 55118 55053
rect 55278 55050 55330 55053
rect 55278 55004 55279 55050
rect 55279 55004 55325 55050
rect 55325 55004 55330 55050
rect 55278 55001 55330 55004
rect 55489 55001 55541 55053
rect 56015 55001 56067 55053
rect 56226 55050 56278 55053
rect 56226 55004 56267 55050
rect 56267 55004 56278 55050
rect 56226 55001 56278 55004
rect 56437 55001 56489 55053
rect 56648 55001 56700 55053
rect 56859 55001 56911 55053
rect 57070 55001 57122 55053
rect 57281 55001 57333 55053
rect 48943 54909 48995 54915
rect 49154 54909 49206 54915
rect 49365 54909 49417 54915
rect 49576 54909 49628 54915
rect 49787 54909 49839 54915
rect 33057 54822 33109 54825
rect 33237 54822 33289 54825
rect 35332 54863 35384 54909
rect 35543 54863 35580 54909
rect 35580 54863 35595 54909
rect 35754 54863 35786 54909
rect 35786 54863 35806 54909
rect 35965 54863 35992 54909
rect 35992 54863 36017 54909
rect 36176 54863 36198 54909
rect 36198 54863 36228 54909
rect 37891 54865 37909 54909
rect 37909 54865 37943 54909
rect 38071 54865 38072 54909
rect 38072 54865 38123 54909
rect 33057 54776 33109 54822
rect 33237 54776 33289 54822
rect 33057 54773 33109 54776
rect 33237 54773 33289 54776
rect 33057 54374 33109 54377
rect 33237 54374 33289 54377
rect 33057 54328 33109 54374
rect 33237 54328 33289 54374
rect 33057 54325 33109 54328
rect 33237 54325 33289 54328
rect 29582 54101 29634 54153
rect 29793 54150 29845 54153
rect 29793 54104 29798 54150
rect 29798 54104 29844 54150
rect 29844 54104 29845 54150
rect 29793 54101 29845 54104
rect 30005 54101 30057 54153
rect 30216 54101 30268 54153
rect 34267 54598 34319 54615
rect 34447 54598 34499 54615
rect 34627 54598 34679 54615
rect 34267 54563 34302 54598
rect 34302 54563 34319 54598
rect 34447 54563 34451 54598
rect 34451 54563 34499 54598
rect 34627 54563 34658 54598
rect 34658 54563 34679 54598
rect 36678 54638 36697 54690
rect 36697 54638 36730 54690
rect 48943 54863 48984 54909
rect 48984 54863 48995 54909
rect 49154 54863 49190 54909
rect 49190 54863 49206 54909
rect 49365 54863 49396 54909
rect 49396 54863 49417 54909
rect 49576 54863 49602 54909
rect 49602 54863 49628 54909
rect 49787 54863 49839 54909
rect 39994 54740 40046 54792
rect 36961 54639 36971 54683
rect 36971 54639 37013 54683
rect 37172 54639 37206 54683
rect 37206 54639 37224 54683
rect 36961 54631 37013 54639
rect 37172 54631 37224 54639
rect 37384 54631 37436 54683
rect 37595 54631 37647 54683
rect 35332 54415 35384 54455
rect 35543 54415 35580 54455
rect 35580 54415 35595 54455
rect 35754 54415 35786 54455
rect 35786 54415 35806 54455
rect 35965 54415 35992 54455
rect 35992 54415 36017 54455
rect 36176 54415 36198 54455
rect 36198 54415 36228 54455
rect 37891 54415 37909 54443
rect 37909 54415 37943 54443
rect 38071 54415 38072 54443
rect 38072 54415 38123 54443
rect 35332 54403 35384 54415
rect 35543 54403 35595 54415
rect 35754 54403 35806 54415
rect 35965 54403 36017 54415
rect 36176 54403 36228 54415
rect 33819 54328 33833 54369
rect 33833 54328 33871 54369
rect 33999 54328 34039 54369
rect 34039 54328 34051 54369
rect 37891 54391 37943 54415
rect 38071 54391 38123 54415
rect 33819 54317 33871 54328
rect 33999 54317 34051 54328
rect 30854 54101 30906 54153
rect 31065 54101 31117 54153
rect 31276 54101 31328 54153
rect 31486 54150 31538 54153
rect 31697 54150 31749 54153
rect 31909 54150 31961 54153
rect 32120 54150 32172 54153
rect 32330 54150 32382 54153
rect 32541 54150 32593 54153
rect 32752 54150 32804 54153
rect 34284 54150 34336 54153
rect 34495 54150 34547 54153
rect 31486 54104 31538 54150
rect 31697 54104 31749 54150
rect 31909 54104 31961 54150
rect 32120 54104 32172 54150
rect 32330 54104 32382 54150
rect 32541 54104 32593 54150
rect 32752 54104 32804 54150
rect 34284 54104 34302 54150
rect 34302 54104 34336 54150
rect 34495 54104 34508 54150
rect 34508 54104 34547 54150
rect 31486 54101 31538 54104
rect 31697 54101 31749 54104
rect 31909 54101 31961 54104
rect 32120 54101 32172 54104
rect 32330 54101 32382 54104
rect 32541 54101 32593 54104
rect 32752 54101 32804 54104
rect 34284 54101 34336 54104
rect 34495 54101 34547 54104
rect 34707 54101 34759 54153
rect 34918 54101 34970 54153
rect 35220 54101 35272 54153
rect 35430 54101 35482 54153
rect 35641 54101 35693 54153
rect 35853 54101 35905 54153
rect 36064 54101 36116 54153
rect 36274 54101 36326 54153
rect 38330 54150 38382 54153
rect 38330 54104 38382 54150
rect 38330 54101 38382 54104
rect 38541 54101 38593 54153
rect 38752 54101 38804 54153
rect 39052 54150 39104 54153
rect 39232 54150 39284 54153
rect 39052 54104 39062 54150
rect 39062 54104 39104 54150
rect 39232 54104 39266 54150
rect 39266 54104 39284 54150
rect 39052 54101 39104 54104
rect 39232 54101 39284 54104
rect 33057 53926 33109 53929
rect 33237 53926 33289 53929
rect 33057 53880 33109 53926
rect 33237 53880 33289 53926
rect 33057 53877 33109 53880
rect 33237 53877 33289 53880
rect 33819 53926 33871 53937
rect 33999 53926 34051 53937
rect 33819 53885 33833 53926
rect 33833 53885 33871 53926
rect 33999 53885 34039 53926
rect 34039 53885 34051 53926
rect 35332 53839 35384 53851
rect 35543 53839 35595 53851
rect 35754 53839 35806 53851
rect 35965 53839 36017 53851
rect 36176 53839 36228 53851
rect 37891 53839 37943 53863
rect 38071 53839 38123 53863
rect 35332 53799 35384 53839
rect 35543 53799 35580 53839
rect 35580 53799 35595 53839
rect 35754 53799 35786 53839
rect 35786 53799 35806 53839
rect 35965 53799 35992 53839
rect 35992 53799 36017 53839
rect 36176 53799 36198 53839
rect 36198 53799 36228 53839
rect 37891 53811 37909 53839
rect 37909 53811 37943 53839
rect 38071 53811 38072 53839
rect 38072 53811 38123 53839
rect 34267 53656 34302 53691
rect 34302 53656 34319 53691
rect 34447 53656 34451 53691
rect 34451 53656 34499 53691
rect 34627 53656 34658 53691
rect 34658 53656 34679 53691
rect 34267 53639 34319 53656
rect 34447 53639 34499 53656
rect 34627 53639 34679 53656
rect 33057 53478 33109 53481
rect 33237 53478 33289 53481
rect 33057 53432 33109 53478
rect 33237 53432 33289 53478
rect 33057 53429 33109 53432
rect 33237 53429 33289 53432
rect 36678 53564 36697 53616
rect 36697 53564 36730 53616
rect 36961 53615 37013 53623
rect 37172 53615 37224 53623
rect 36961 53571 36971 53615
rect 36971 53571 37013 53615
rect 37172 53571 37206 53615
rect 37206 53571 37224 53615
rect 37384 53571 37436 53623
rect 37595 53571 37647 53623
rect 39994 54554 40046 54606
rect 39775 54374 39827 54391
rect 39775 54339 39786 54374
rect 39786 54339 39827 54374
rect 42690 54570 42742 54622
rect 41935 54339 41987 54391
rect 46731 54679 46783 54731
rect 48596 54725 48648 54777
rect 51835 54822 51887 54847
rect 52015 54822 52067 54847
rect 51835 54795 51887 54822
rect 52015 54795 52067 54822
rect 44939 54598 44991 54615
rect 45151 54598 45203 54615
rect 44939 54563 44971 54598
rect 44971 54563 44991 54598
rect 45151 54563 45197 54598
rect 45197 54563 45203 54598
rect 48596 54507 48648 54559
rect 50300 54563 50352 54615
rect 50511 54598 50563 54615
rect 50511 54563 50513 54598
rect 50513 54563 50563 54598
rect 50722 54563 50774 54615
rect 48943 54415 48984 54452
rect 48984 54415 48995 54452
rect 49154 54415 49190 54452
rect 49190 54415 49206 54452
rect 49365 54415 49396 54452
rect 49396 54415 49417 54452
rect 49576 54415 49602 54452
rect 49602 54415 49628 54452
rect 49787 54415 49839 54452
rect 48943 54400 48995 54415
rect 49154 54400 49206 54415
rect 49365 54400 49417 54415
rect 49576 54400 49628 54415
rect 49787 54400 49839 54415
rect 51073 54374 51125 54377
rect 51253 54374 51305 54377
rect 51073 54328 51086 54374
rect 51086 54328 51125 54374
rect 51253 54328 51292 54374
rect 51292 54328 51305 54374
rect 51073 54325 51125 54328
rect 51253 54325 51305 54328
rect 51835 54374 51887 54384
rect 52015 54374 52067 54384
rect 51835 54332 51887 54374
rect 52015 54332 52067 54374
rect 40253 54101 40305 54153
rect 40433 54101 40485 54153
rect 43790 54101 43842 54153
rect 44001 54101 44053 54153
rect 44213 54150 44265 54153
rect 44213 54104 44236 54150
rect 44236 54104 44265 54150
rect 44213 54101 44265 54104
rect 44424 54101 44476 54153
rect 44834 54150 44886 54153
rect 45045 54150 45097 54153
rect 45256 54150 45308 54153
rect 44834 54104 44858 54150
rect 44858 54104 44886 54150
rect 45045 54104 45084 54150
rect 45084 54104 45097 54150
rect 45256 54104 45264 54150
rect 45264 54104 45308 54150
rect 44834 54101 44886 54104
rect 45045 54101 45097 54104
rect 45256 54101 45308 54104
rect 48838 54101 48890 54153
rect 49048 54101 49100 54153
rect 49259 54101 49311 54153
rect 49471 54101 49523 54153
rect 49682 54101 49734 54153
rect 49892 54101 49944 54153
rect 50346 54101 50398 54153
rect 50557 54150 50609 54153
rect 50768 54150 50820 54153
rect 52316 54150 52368 54153
rect 52527 54150 52579 54153
rect 52738 54150 52790 54153
rect 52948 54150 53000 54153
rect 53159 54150 53211 54153
rect 53371 54150 53423 54153
rect 53582 54150 53634 54153
rect 50557 54104 50571 54150
rect 50571 54104 50609 54150
rect 50768 54104 50777 54150
rect 50777 54104 50820 54150
rect 52316 54104 52368 54150
rect 52527 54104 52579 54150
rect 52738 54104 52790 54150
rect 52948 54104 53000 54150
rect 53159 54104 53211 54150
rect 53371 54104 53423 54150
rect 53582 54104 53634 54150
rect 50557 54101 50609 54104
rect 50768 54101 50820 54104
rect 39775 53880 39786 53915
rect 39786 53880 39827 53915
rect 39775 53863 39827 53880
rect 39994 53648 40046 53700
rect 39994 53462 40046 53514
rect 52316 54101 52368 54104
rect 52527 54101 52579 54104
rect 52738 54101 52790 54104
rect 52948 54101 53000 54104
rect 53159 54101 53211 54104
rect 53371 54101 53423 54104
rect 53582 54101 53634 54104
rect 53792 54101 53844 54153
rect 54003 54101 54055 54153
rect 54214 54101 54266 54153
rect 54855 54101 54907 54153
rect 55066 54101 55118 54153
rect 55278 54150 55330 54153
rect 55278 54104 55279 54150
rect 55279 54104 55325 54150
rect 55325 54104 55330 54150
rect 55278 54101 55330 54104
rect 55489 54101 55541 54153
rect 41935 53863 41987 53915
rect 51073 53926 51125 53929
rect 51253 53926 51305 53929
rect 42690 53632 42742 53684
rect 51073 53880 51086 53926
rect 51086 53880 51125 53926
rect 51253 53880 51292 53926
rect 51292 53880 51305 53926
rect 48943 53839 48995 53854
rect 49154 53839 49206 53854
rect 49365 53839 49417 53854
rect 49576 53839 49628 53854
rect 49787 53839 49839 53854
rect 48943 53802 48984 53839
rect 48984 53802 48995 53839
rect 49154 53802 49190 53839
rect 49190 53802 49206 53839
rect 49365 53802 49396 53839
rect 49396 53802 49417 53839
rect 49576 53802 49602 53839
rect 49602 53802 49628 53839
rect 49787 53802 49839 53839
rect 51073 53877 51125 53880
rect 51253 53877 51305 53880
rect 44939 53656 44971 53691
rect 44971 53656 44991 53691
rect 45151 53656 45197 53691
rect 45197 53656 45203 53691
rect 48596 53695 48648 53747
rect 44939 53639 44991 53656
rect 45151 53639 45203 53656
rect 47108 53523 47160 53575
rect 50300 53639 50352 53691
rect 50511 53656 50513 53691
rect 50513 53656 50563 53691
rect 50511 53639 50563 53656
rect 50722 53639 50774 53691
rect 48596 53477 48648 53529
rect 51835 53880 51887 53922
rect 52015 53880 52067 53922
rect 51835 53870 51887 53880
rect 52015 53870 52067 53880
rect 35332 53345 35384 53391
rect 35543 53345 35580 53391
rect 35580 53345 35595 53391
rect 35754 53345 35786 53391
rect 35786 53345 35806 53391
rect 35965 53345 35992 53391
rect 35992 53345 36017 53391
rect 36176 53345 36198 53391
rect 36198 53345 36228 53391
rect 37891 53345 37909 53389
rect 37909 53345 37943 53389
rect 38071 53345 38072 53389
rect 38072 53345 38123 53389
rect 48943 53345 48984 53391
rect 48984 53345 48995 53391
rect 49154 53345 49190 53391
rect 49190 53345 49206 53391
rect 49365 53345 49396 53391
rect 49396 53345 49417 53391
rect 49576 53345 49602 53391
rect 49602 53345 49628 53391
rect 49787 53345 49839 53391
rect 51835 53432 51887 53459
rect 52015 53432 52067 53459
rect 51835 53407 51887 53432
rect 52015 53407 52067 53432
rect 35332 53339 35384 53345
rect 35543 53339 35595 53345
rect 35754 53339 35806 53345
rect 35965 53339 36017 53345
rect 36176 53339 36228 53345
rect 37891 53337 37943 53345
rect 38071 53337 38123 53345
rect 27790 53201 27842 53253
rect 28001 53201 28053 53253
rect 28212 53201 28264 53253
rect 28423 53201 28475 53253
rect 28634 53201 28686 53253
rect 28845 53250 28897 53253
rect 28845 53204 28856 53250
rect 28856 53204 28897 53250
rect 28845 53201 28897 53204
rect 29056 53201 29108 53253
rect 29582 53201 29634 53253
rect 29793 53250 29845 53253
rect 29793 53204 29798 53250
rect 29798 53204 29844 53250
rect 29844 53204 29845 53250
rect 29793 53201 29845 53204
rect 30005 53201 30057 53253
rect 30216 53201 30268 53253
rect 30854 53201 30906 53253
rect 31065 53201 31117 53253
rect 31276 53201 31328 53253
rect 31486 53201 31538 53253
rect 31697 53201 31749 53253
rect 31909 53201 31961 53253
rect 32120 53201 32172 53253
rect 32330 53201 32382 53253
rect 32541 53201 32593 53253
rect 32752 53201 32804 53253
rect 48943 53339 48995 53345
rect 49154 53339 49206 53345
rect 49365 53339 49417 53345
rect 49576 53339 49628 53345
rect 49787 53339 49839 53345
rect 34755 53201 34807 53253
rect 34935 53250 34987 53253
rect 34935 53204 34962 53250
rect 34962 53204 34987 53250
rect 34935 53201 34987 53204
rect 50138 53250 50190 53253
rect 50138 53204 50160 53250
rect 50160 53204 50190 53250
rect 50138 53201 50190 53204
rect 50318 53201 50370 53253
rect 35332 53109 35384 53115
rect 35543 53109 35595 53115
rect 35754 53109 35806 53115
rect 35965 53109 36017 53115
rect 36176 53109 36228 53115
rect 37891 53109 37943 53117
rect 38071 53109 38123 53117
rect 52316 53201 52368 53253
rect 52527 53201 52579 53253
rect 52738 53201 52790 53253
rect 52948 53201 53000 53253
rect 53159 53201 53211 53253
rect 53371 53201 53423 53253
rect 53582 53201 53634 53253
rect 53792 53201 53844 53253
rect 54003 53201 54055 53253
rect 54214 53201 54266 53253
rect 54855 53201 54907 53253
rect 55066 53201 55118 53253
rect 55278 53250 55330 53253
rect 55278 53204 55279 53250
rect 55279 53204 55325 53250
rect 55325 53204 55330 53250
rect 55278 53201 55330 53204
rect 55489 53201 55541 53253
rect 56015 53201 56067 53253
rect 56226 53250 56278 53253
rect 56226 53204 56267 53250
rect 56267 53204 56278 53250
rect 56226 53201 56278 53204
rect 56437 53201 56489 53253
rect 56648 53201 56700 53253
rect 56859 53201 56911 53253
rect 57070 53201 57122 53253
rect 57281 53201 57333 53253
rect 48943 53109 48995 53115
rect 49154 53109 49206 53115
rect 49365 53109 49417 53115
rect 49576 53109 49628 53115
rect 49787 53109 49839 53115
rect 33057 53022 33109 53025
rect 33237 53022 33289 53025
rect 35332 53063 35384 53109
rect 35543 53063 35580 53109
rect 35580 53063 35595 53109
rect 35754 53063 35786 53109
rect 35786 53063 35806 53109
rect 35965 53063 35992 53109
rect 35992 53063 36017 53109
rect 36176 53063 36198 53109
rect 36198 53063 36228 53109
rect 37891 53065 37909 53109
rect 37909 53065 37943 53109
rect 38071 53065 38072 53109
rect 38072 53065 38123 53109
rect 33057 52976 33109 53022
rect 33237 52976 33289 53022
rect 33057 52973 33109 52976
rect 33237 52973 33289 52976
rect 33057 52574 33109 52577
rect 33237 52574 33289 52577
rect 33057 52528 33109 52574
rect 33237 52528 33289 52574
rect 33057 52525 33109 52528
rect 33237 52525 33289 52528
rect 29582 52301 29634 52353
rect 29793 52350 29845 52353
rect 29793 52304 29798 52350
rect 29798 52304 29844 52350
rect 29844 52304 29845 52350
rect 29793 52301 29845 52304
rect 30005 52301 30057 52353
rect 30216 52301 30268 52353
rect 34267 52798 34319 52815
rect 34447 52798 34499 52815
rect 34627 52798 34679 52815
rect 34267 52763 34302 52798
rect 34302 52763 34319 52798
rect 34447 52763 34451 52798
rect 34451 52763 34499 52798
rect 34627 52763 34658 52798
rect 34658 52763 34679 52798
rect 36678 52838 36697 52890
rect 36697 52838 36730 52890
rect 48943 53063 48984 53109
rect 48984 53063 48995 53109
rect 49154 53063 49190 53109
rect 49190 53063 49206 53109
rect 49365 53063 49396 53109
rect 49396 53063 49417 53109
rect 49576 53063 49602 53109
rect 49602 53063 49628 53109
rect 49787 53063 49839 53109
rect 39994 52940 40046 52992
rect 36961 52839 36971 52883
rect 36971 52839 37013 52883
rect 37172 52839 37206 52883
rect 37206 52839 37224 52883
rect 36961 52831 37013 52839
rect 37172 52831 37224 52839
rect 37384 52831 37436 52883
rect 37595 52831 37647 52883
rect 35332 52615 35384 52655
rect 35543 52615 35580 52655
rect 35580 52615 35595 52655
rect 35754 52615 35786 52655
rect 35786 52615 35806 52655
rect 35965 52615 35992 52655
rect 35992 52615 36017 52655
rect 36176 52615 36198 52655
rect 36198 52615 36228 52655
rect 37891 52615 37909 52643
rect 37909 52615 37943 52643
rect 38071 52615 38072 52643
rect 38072 52615 38123 52643
rect 35332 52603 35384 52615
rect 35543 52603 35595 52615
rect 35754 52603 35806 52615
rect 35965 52603 36017 52615
rect 36176 52603 36228 52615
rect 33819 52528 33833 52569
rect 33833 52528 33871 52569
rect 33999 52528 34039 52569
rect 34039 52528 34051 52569
rect 37891 52591 37943 52615
rect 38071 52591 38123 52615
rect 33819 52517 33871 52528
rect 33999 52517 34051 52528
rect 30854 52301 30906 52353
rect 31065 52301 31117 52353
rect 31276 52301 31328 52353
rect 31486 52350 31538 52353
rect 31697 52350 31749 52353
rect 31909 52350 31961 52353
rect 32120 52350 32172 52353
rect 32330 52350 32382 52353
rect 32541 52350 32593 52353
rect 32752 52350 32804 52353
rect 34284 52350 34336 52353
rect 34495 52350 34547 52353
rect 31486 52304 31538 52350
rect 31697 52304 31749 52350
rect 31909 52304 31961 52350
rect 32120 52304 32172 52350
rect 32330 52304 32382 52350
rect 32541 52304 32593 52350
rect 32752 52304 32804 52350
rect 34284 52304 34302 52350
rect 34302 52304 34336 52350
rect 34495 52304 34508 52350
rect 34508 52304 34547 52350
rect 31486 52301 31538 52304
rect 31697 52301 31749 52304
rect 31909 52301 31961 52304
rect 32120 52301 32172 52304
rect 32330 52301 32382 52304
rect 32541 52301 32593 52304
rect 32752 52301 32804 52304
rect 34284 52301 34336 52304
rect 34495 52301 34547 52304
rect 34707 52301 34759 52353
rect 34918 52301 34970 52353
rect 35220 52301 35272 52353
rect 35430 52301 35482 52353
rect 35641 52301 35693 52353
rect 35853 52301 35905 52353
rect 36064 52301 36116 52353
rect 36274 52301 36326 52353
rect 38330 52350 38382 52353
rect 38330 52304 38382 52350
rect 38330 52301 38382 52304
rect 38541 52301 38593 52353
rect 38752 52301 38804 52353
rect 39052 52350 39104 52353
rect 39232 52350 39284 52353
rect 39052 52304 39062 52350
rect 39062 52304 39104 52350
rect 39232 52304 39266 52350
rect 39266 52304 39284 52350
rect 39052 52301 39104 52304
rect 39232 52301 39284 52304
rect 33057 52126 33109 52129
rect 33237 52126 33289 52129
rect 33057 52080 33109 52126
rect 33237 52080 33289 52126
rect 33057 52077 33109 52080
rect 33237 52077 33289 52080
rect 33819 52126 33871 52137
rect 33999 52126 34051 52137
rect 33819 52085 33833 52126
rect 33833 52085 33871 52126
rect 33999 52085 34039 52126
rect 34039 52085 34051 52126
rect 35332 52039 35384 52051
rect 35543 52039 35595 52051
rect 35754 52039 35806 52051
rect 35965 52039 36017 52051
rect 36176 52039 36228 52051
rect 37891 52039 37943 52063
rect 38071 52039 38123 52063
rect 35332 51999 35384 52039
rect 35543 51999 35580 52039
rect 35580 51999 35595 52039
rect 35754 51999 35786 52039
rect 35786 51999 35806 52039
rect 35965 51999 35992 52039
rect 35992 51999 36017 52039
rect 36176 51999 36198 52039
rect 36198 51999 36228 52039
rect 37891 52011 37909 52039
rect 37909 52011 37943 52039
rect 38071 52011 38072 52039
rect 38072 52011 38123 52039
rect 34267 51856 34302 51891
rect 34302 51856 34319 51891
rect 34447 51856 34451 51891
rect 34451 51856 34499 51891
rect 34627 51856 34658 51891
rect 34658 51856 34679 51891
rect 34267 51839 34319 51856
rect 34447 51839 34499 51856
rect 34627 51839 34679 51856
rect 33057 51678 33109 51681
rect 33237 51678 33289 51681
rect 33057 51632 33109 51678
rect 33237 51632 33289 51678
rect 33057 51629 33109 51632
rect 33237 51629 33289 51632
rect 36678 51764 36697 51816
rect 36697 51764 36730 51816
rect 36961 51815 37013 51823
rect 37172 51815 37224 51823
rect 36961 51771 36971 51815
rect 36971 51771 37013 51815
rect 37172 51771 37206 51815
rect 37206 51771 37224 51815
rect 37384 51771 37436 51823
rect 37595 51771 37647 51823
rect 39994 52754 40046 52806
rect 39775 52574 39827 52591
rect 39775 52539 39786 52574
rect 39786 52539 39827 52574
rect 42690 52770 42742 52822
rect 41935 52539 41987 52591
rect 47486 52879 47538 52931
rect 48596 52925 48648 52977
rect 51835 53022 51887 53047
rect 52015 53022 52067 53047
rect 51835 52995 51887 53022
rect 52015 52995 52067 53022
rect 44939 52798 44991 52815
rect 45151 52798 45203 52815
rect 44939 52763 44971 52798
rect 44971 52763 44991 52798
rect 45151 52763 45197 52798
rect 45197 52763 45203 52798
rect 48596 52707 48648 52759
rect 50300 52763 50352 52815
rect 50511 52798 50563 52815
rect 50511 52763 50513 52798
rect 50513 52763 50563 52798
rect 50722 52763 50774 52815
rect 48943 52615 48984 52652
rect 48984 52615 48995 52652
rect 49154 52615 49190 52652
rect 49190 52615 49206 52652
rect 49365 52615 49396 52652
rect 49396 52615 49417 52652
rect 49576 52615 49602 52652
rect 49602 52615 49628 52652
rect 49787 52615 49839 52652
rect 48943 52600 48995 52615
rect 49154 52600 49206 52615
rect 49365 52600 49417 52615
rect 49576 52600 49628 52615
rect 49787 52600 49839 52615
rect 51073 52574 51125 52577
rect 51253 52574 51305 52577
rect 51073 52528 51086 52574
rect 51086 52528 51125 52574
rect 51253 52528 51292 52574
rect 51292 52528 51305 52574
rect 51073 52525 51125 52528
rect 51253 52525 51305 52528
rect 51835 52574 51887 52584
rect 52015 52574 52067 52584
rect 51835 52532 51887 52574
rect 52015 52532 52067 52574
rect 40253 52301 40305 52353
rect 40433 52301 40485 52353
rect 43790 52301 43842 52353
rect 44001 52301 44053 52353
rect 44213 52350 44265 52353
rect 44213 52304 44236 52350
rect 44236 52304 44265 52350
rect 44213 52301 44265 52304
rect 44424 52301 44476 52353
rect 44834 52350 44886 52353
rect 45045 52350 45097 52353
rect 45256 52350 45308 52353
rect 44834 52304 44858 52350
rect 44858 52304 44886 52350
rect 45045 52304 45084 52350
rect 45084 52304 45097 52350
rect 45256 52304 45264 52350
rect 45264 52304 45308 52350
rect 44834 52301 44886 52304
rect 45045 52301 45097 52304
rect 45256 52301 45308 52304
rect 48838 52301 48890 52353
rect 49048 52301 49100 52353
rect 49259 52301 49311 52353
rect 49471 52301 49523 52353
rect 49682 52301 49734 52353
rect 49892 52301 49944 52353
rect 50346 52301 50398 52353
rect 50557 52350 50609 52353
rect 50768 52350 50820 52353
rect 52316 52350 52368 52353
rect 52527 52350 52579 52353
rect 52738 52350 52790 52353
rect 52948 52350 53000 52353
rect 53159 52350 53211 52353
rect 53371 52350 53423 52353
rect 53582 52350 53634 52353
rect 50557 52304 50571 52350
rect 50571 52304 50609 52350
rect 50768 52304 50777 52350
rect 50777 52304 50820 52350
rect 52316 52304 52368 52350
rect 52527 52304 52579 52350
rect 52738 52304 52790 52350
rect 52948 52304 53000 52350
rect 53159 52304 53211 52350
rect 53371 52304 53423 52350
rect 53582 52304 53634 52350
rect 50557 52301 50609 52304
rect 50768 52301 50820 52304
rect 39775 52080 39786 52115
rect 39786 52080 39827 52115
rect 39775 52063 39827 52080
rect 39994 51848 40046 51900
rect 39994 51662 40046 51714
rect 52316 52301 52368 52304
rect 52527 52301 52579 52304
rect 52738 52301 52790 52304
rect 52948 52301 53000 52304
rect 53159 52301 53211 52304
rect 53371 52301 53423 52304
rect 53582 52301 53634 52304
rect 53792 52301 53844 52353
rect 54003 52301 54055 52353
rect 54214 52301 54266 52353
rect 54855 52301 54907 52353
rect 55066 52301 55118 52353
rect 55278 52350 55330 52353
rect 55278 52304 55279 52350
rect 55279 52304 55325 52350
rect 55325 52304 55330 52350
rect 55278 52301 55330 52304
rect 55489 52301 55541 52353
rect 41935 52063 41987 52115
rect 51073 52126 51125 52129
rect 51253 52126 51305 52129
rect 42690 51832 42742 51884
rect 51073 52080 51086 52126
rect 51086 52080 51125 52126
rect 51253 52080 51292 52126
rect 51292 52080 51305 52126
rect 48943 52039 48995 52054
rect 49154 52039 49206 52054
rect 49365 52039 49417 52054
rect 49576 52039 49628 52054
rect 49787 52039 49839 52054
rect 48943 52002 48984 52039
rect 48984 52002 48995 52039
rect 49154 52002 49190 52039
rect 49190 52002 49206 52039
rect 49365 52002 49396 52039
rect 49396 52002 49417 52039
rect 49576 52002 49602 52039
rect 49602 52002 49628 52039
rect 49787 52002 49839 52039
rect 51073 52077 51125 52080
rect 51253 52077 51305 52080
rect 44939 51856 44971 51891
rect 44971 51856 44991 51891
rect 45151 51856 45197 51891
rect 45197 51856 45203 51891
rect 48596 51895 48648 51947
rect 44939 51839 44991 51856
rect 45151 51839 45203 51856
rect 47864 51723 47916 51775
rect 50300 51839 50352 51891
rect 50511 51856 50513 51891
rect 50513 51856 50563 51891
rect 50511 51839 50563 51856
rect 50722 51839 50774 51891
rect 48596 51677 48648 51729
rect 51835 52080 51887 52122
rect 52015 52080 52067 52122
rect 51835 52070 51887 52080
rect 52015 52070 52067 52080
rect 35332 51545 35384 51591
rect 35543 51545 35580 51591
rect 35580 51545 35595 51591
rect 35754 51545 35786 51591
rect 35786 51545 35806 51591
rect 35965 51545 35992 51591
rect 35992 51545 36017 51591
rect 36176 51545 36198 51591
rect 36198 51545 36228 51591
rect 37891 51545 37909 51589
rect 37909 51545 37943 51589
rect 38071 51545 38072 51589
rect 38072 51545 38123 51589
rect 48943 51545 48984 51591
rect 48984 51545 48995 51591
rect 49154 51545 49190 51591
rect 49190 51545 49206 51591
rect 49365 51545 49396 51591
rect 49396 51545 49417 51591
rect 49576 51545 49602 51591
rect 49602 51545 49628 51591
rect 49787 51545 49839 51591
rect 51835 51632 51887 51659
rect 52015 51632 52067 51659
rect 51835 51607 51887 51632
rect 52015 51607 52067 51632
rect 35332 51539 35384 51545
rect 35543 51539 35595 51545
rect 35754 51539 35806 51545
rect 35965 51539 36017 51545
rect 36176 51539 36228 51545
rect 37891 51537 37943 51545
rect 38071 51537 38123 51545
rect 27790 51401 27842 51453
rect 28001 51401 28053 51453
rect 28212 51401 28264 51453
rect 28423 51401 28475 51453
rect 28634 51401 28686 51453
rect 28845 51450 28897 51453
rect 28845 51404 28856 51450
rect 28856 51404 28897 51450
rect 28845 51401 28897 51404
rect 29056 51401 29108 51453
rect 29582 51401 29634 51453
rect 29793 51450 29845 51453
rect 29793 51404 29798 51450
rect 29798 51404 29844 51450
rect 29844 51404 29845 51450
rect 29793 51401 29845 51404
rect 30005 51401 30057 51453
rect 30216 51401 30268 51453
rect 30854 51401 30906 51453
rect 31065 51401 31117 51453
rect 31276 51401 31328 51453
rect 31486 51401 31538 51453
rect 31697 51401 31749 51453
rect 31909 51401 31961 51453
rect 32120 51401 32172 51453
rect 32330 51401 32382 51453
rect 32541 51401 32593 51453
rect 32752 51401 32804 51453
rect 48943 51539 48995 51545
rect 49154 51539 49206 51545
rect 49365 51539 49417 51545
rect 49576 51539 49628 51545
rect 49787 51539 49839 51545
rect 34755 51401 34807 51453
rect 34935 51450 34987 51453
rect 34935 51404 34962 51450
rect 34962 51404 34987 51450
rect 34935 51401 34987 51404
rect 50138 51450 50190 51453
rect 50138 51404 50160 51450
rect 50160 51404 50190 51450
rect 50138 51401 50190 51404
rect 50318 51401 50370 51453
rect 35332 51309 35384 51315
rect 35543 51309 35595 51315
rect 35754 51309 35806 51315
rect 35965 51309 36017 51315
rect 36176 51309 36228 51315
rect 37891 51309 37943 51317
rect 38071 51309 38123 51317
rect 52316 51401 52368 51453
rect 52527 51401 52579 51453
rect 52738 51401 52790 51453
rect 52948 51401 53000 51453
rect 53159 51401 53211 51453
rect 53371 51401 53423 51453
rect 53582 51401 53634 51453
rect 53792 51401 53844 51453
rect 54003 51401 54055 51453
rect 54214 51401 54266 51453
rect 54855 51401 54907 51453
rect 55066 51401 55118 51453
rect 55278 51450 55330 51453
rect 55278 51404 55279 51450
rect 55279 51404 55325 51450
rect 55325 51404 55330 51450
rect 55278 51401 55330 51404
rect 55489 51401 55541 51453
rect 56015 51401 56067 51453
rect 56226 51450 56278 51453
rect 56226 51404 56267 51450
rect 56267 51404 56278 51450
rect 56226 51401 56278 51404
rect 56437 51401 56489 51453
rect 56648 51401 56700 51453
rect 56859 51401 56911 51453
rect 57070 51401 57122 51453
rect 57281 51401 57333 51453
rect 48943 51309 48995 51315
rect 49154 51309 49206 51315
rect 49365 51309 49417 51315
rect 49576 51309 49628 51315
rect 49787 51309 49839 51315
rect 33057 51222 33109 51225
rect 33237 51222 33289 51225
rect 35332 51263 35384 51309
rect 35543 51263 35580 51309
rect 35580 51263 35595 51309
rect 35754 51263 35786 51309
rect 35786 51263 35806 51309
rect 35965 51263 35992 51309
rect 35992 51263 36017 51309
rect 36176 51263 36198 51309
rect 36198 51263 36228 51309
rect 37891 51265 37909 51309
rect 37909 51265 37943 51309
rect 38071 51265 38072 51309
rect 38072 51265 38123 51309
rect 33057 51176 33109 51222
rect 33237 51176 33289 51222
rect 33057 51173 33109 51176
rect 33237 51173 33289 51176
rect 33057 50774 33109 50777
rect 33237 50774 33289 50777
rect 33057 50728 33109 50774
rect 33237 50728 33289 50774
rect 33057 50725 33109 50728
rect 33237 50725 33289 50728
rect 29582 50501 29634 50553
rect 29793 50550 29845 50553
rect 29793 50504 29798 50550
rect 29798 50504 29844 50550
rect 29844 50504 29845 50550
rect 29793 50501 29845 50504
rect 30005 50501 30057 50553
rect 30216 50501 30268 50553
rect 34267 50998 34319 51015
rect 34447 50998 34499 51015
rect 34627 50998 34679 51015
rect 34267 50963 34302 50998
rect 34302 50963 34319 50998
rect 34447 50963 34451 50998
rect 34451 50963 34499 50998
rect 34627 50963 34658 50998
rect 34658 50963 34679 50998
rect 36678 51038 36697 51090
rect 36697 51038 36730 51090
rect 48943 51263 48984 51309
rect 48984 51263 48995 51309
rect 49154 51263 49190 51309
rect 49190 51263 49206 51309
rect 49365 51263 49396 51309
rect 49396 51263 49417 51309
rect 49576 51263 49602 51309
rect 49602 51263 49628 51309
rect 49787 51263 49839 51309
rect 39994 51140 40046 51192
rect 36961 51039 36971 51083
rect 36971 51039 37013 51083
rect 37172 51039 37206 51083
rect 37206 51039 37224 51083
rect 36961 51031 37013 51039
rect 37172 51031 37224 51039
rect 37384 51031 37436 51083
rect 37595 51031 37647 51083
rect 35332 50815 35384 50855
rect 35543 50815 35580 50855
rect 35580 50815 35595 50855
rect 35754 50815 35786 50855
rect 35786 50815 35806 50855
rect 35965 50815 35992 50855
rect 35992 50815 36017 50855
rect 36176 50815 36198 50855
rect 36198 50815 36228 50855
rect 37891 50815 37909 50843
rect 37909 50815 37943 50843
rect 38071 50815 38072 50843
rect 38072 50815 38123 50843
rect 35332 50803 35384 50815
rect 35543 50803 35595 50815
rect 35754 50803 35806 50815
rect 35965 50803 36017 50815
rect 36176 50803 36228 50815
rect 33819 50728 33833 50769
rect 33833 50728 33871 50769
rect 33999 50728 34039 50769
rect 34039 50728 34051 50769
rect 37891 50791 37943 50815
rect 38071 50791 38123 50815
rect 33819 50717 33871 50728
rect 33999 50717 34051 50728
rect 30854 50501 30906 50553
rect 31065 50501 31117 50553
rect 31276 50501 31328 50553
rect 31486 50550 31538 50553
rect 31697 50550 31749 50553
rect 31909 50550 31961 50553
rect 32120 50550 32172 50553
rect 32330 50550 32382 50553
rect 32541 50550 32593 50553
rect 32752 50550 32804 50553
rect 34284 50550 34336 50553
rect 34495 50550 34547 50553
rect 31486 50504 31538 50550
rect 31697 50504 31749 50550
rect 31909 50504 31961 50550
rect 32120 50504 32172 50550
rect 32330 50504 32382 50550
rect 32541 50504 32593 50550
rect 32752 50504 32804 50550
rect 34284 50504 34302 50550
rect 34302 50504 34336 50550
rect 34495 50504 34508 50550
rect 34508 50504 34547 50550
rect 31486 50501 31538 50504
rect 31697 50501 31749 50504
rect 31909 50501 31961 50504
rect 32120 50501 32172 50504
rect 32330 50501 32382 50504
rect 32541 50501 32593 50504
rect 32752 50501 32804 50504
rect 34284 50501 34336 50504
rect 34495 50501 34547 50504
rect 34707 50501 34759 50553
rect 34918 50501 34970 50553
rect 35220 50501 35272 50553
rect 35430 50501 35482 50553
rect 35641 50501 35693 50553
rect 35853 50501 35905 50553
rect 36064 50501 36116 50553
rect 36274 50501 36326 50553
rect 38330 50550 38382 50553
rect 38330 50504 38382 50550
rect 38330 50501 38382 50504
rect 38541 50501 38593 50553
rect 38752 50501 38804 50553
rect 39052 50550 39104 50553
rect 39232 50550 39284 50553
rect 39052 50504 39062 50550
rect 39062 50504 39104 50550
rect 39232 50504 39266 50550
rect 39266 50504 39284 50550
rect 39052 50501 39104 50504
rect 39232 50501 39284 50504
rect 33057 50326 33109 50329
rect 33237 50326 33289 50329
rect 33057 50280 33109 50326
rect 33237 50280 33289 50326
rect 33057 50277 33109 50280
rect 33237 50277 33289 50280
rect 33819 50326 33871 50337
rect 33999 50326 34051 50337
rect 33819 50285 33833 50326
rect 33833 50285 33871 50326
rect 33999 50285 34039 50326
rect 34039 50285 34051 50326
rect 35332 50239 35384 50251
rect 35543 50239 35595 50251
rect 35754 50239 35806 50251
rect 35965 50239 36017 50251
rect 36176 50239 36228 50251
rect 37891 50239 37943 50263
rect 38071 50239 38123 50263
rect 35332 50199 35384 50239
rect 35543 50199 35580 50239
rect 35580 50199 35595 50239
rect 35754 50199 35786 50239
rect 35786 50199 35806 50239
rect 35965 50199 35992 50239
rect 35992 50199 36017 50239
rect 36176 50199 36198 50239
rect 36198 50199 36228 50239
rect 37891 50211 37909 50239
rect 37909 50211 37943 50239
rect 38071 50211 38072 50239
rect 38072 50211 38123 50239
rect 34267 50056 34302 50091
rect 34302 50056 34319 50091
rect 34447 50056 34451 50091
rect 34451 50056 34499 50091
rect 34627 50056 34658 50091
rect 34658 50056 34679 50091
rect 34267 50039 34319 50056
rect 34447 50039 34499 50056
rect 34627 50039 34679 50056
rect 33057 49878 33109 49881
rect 33237 49878 33289 49881
rect 33057 49832 33109 49878
rect 33237 49832 33289 49878
rect 33057 49829 33109 49832
rect 33237 49829 33289 49832
rect 36678 49964 36697 50016
rect 36697 49964 36730 50016
rect 36961 50015 37013 50023
rect 37172 50015 37224 50023
rect 36961 49971 36971 50015
rect 36971 49971 37013 50015
rect 37172 49971 37206 50015
rect 37206 49971 37224 50015
rect 37384 49971 37436 50023
rect 37595 49971 37647 50023
rect 39994 50954 40046 51006
rect 39775 50774 39827 50791
rect 39775 50739 39786 50774
rect 39786 50739 39827 50774
rect 42690 50970 42742 51022
rect 41935 50739 41987 50791
rect 48241 51079 48293 51131
rect 48596 51125 48648 51177
rect 51835 51222 51887 51247
rect 52015 51222 52067 51247
rect 51835 51195 51887 51222
rect 52015 51195 52067 51222
rect 44939 50998 44991 51015
rect 45151 50998 45203 51015
rect 44939 50963 44971 50998
rect 44971 50963 44991 50998
rect 45151 50963 45197 50998
rect 45197 50963 45203 50998
rect 48596 50907 48648 50959
rect 50300 50963 50352 51015
rect 50511 50998 50563 51015
rect 50511 50963 50513 50998
rect 50513 50963 50563 50998
rect 50722 50963 50774 51015
rect 48943 50815 48984 50852
rect 48984 50815 48995 50852
rect 49154 50815 49190 50852
rect 49190 50815 49206 50852
rect 49365 50815 49396 50852
rect 49396 50815 49417 50852
rect 49576 50815 49602 50852
rect 49602 50815 49628 50852
rect 49787 50815 49839 50852
rect 48943 50800 48995 50815
rect 49154 50800 49206 50815
rect 49365 50800 49417 50815
rect 49576 50800 49628 50815
rect 49787 50800 49839 50815
rect 51073 50774 51125 50777
rect 51253 50774 51305 50777
rect 51073 50728 51086 50774
rect 51086 50728 51125 50774
rect 51253 50728 51292 50774
rect 51292 50728 51305 50774
rect 51073 50725 51125 50728
rect 51253 50725 51305 50728
rect 51835 50774 51887 50784
rect 52015 50774 52067 50784
rect 51835 50732 51887 50774
rect 52015 50732 52067 50774
rect 40253 50501 40305 50553
rect 40433 50501 40485 50553
rect 43790 50501 43842 50553
rect 44001 50501 44053 50553
rect 44213 50550 44265 50553
rect 44213 50504 44236 50550
rect 44236 50504 44265 50550
rect 44213 50501 44265 50504
rect 44424 50501 44476 50553
rect 44834 50550 44886 50553
rect 45045 50550 45097 50553
rect 45256 50550 45308 50553
rect 44834 50504 44858 50550
rect 44858 50504 44886 50550
rect 45045 50504 45084 50550
rect 45084 50504 45097 50550
rect 45256 50504 45264 50550
rect 45264 50504 45308 50550
rect 44834 50501 44886 50504
rect 45045 50501 45097 50504
rect 45256 50501 45308 50504
rect 48838 50501 48890 50553
rect 49048 50501 49100 50553
rect 49259 50501 49311 50553
rect 49471 50501 49523 50553
rect 49682 50501 49734 50553
rect 49892 50501 49944 50553
rect 50346 50501 50398 50553
rect 50557 50550 50609 50553
rect 50768 50550 50820 50553
rect 52316 50550 52368 50553
rect 52527 50550 52579 50553
rect 52738 50550 52790 50553
rect 52948 50550 53000 50553
rect 53159 50550 53211 50553
rect 53371 50550 53423 50553
rect 53582 50550 53634 50553
rect 50557 50504 50571 50550
rect 50571 50504 50609 50550
rect 50768 50504 50777 50550
rect 50777 50504 50820 50550
rect 52316 50504 52368 50550
rect 52527 50504 52579 50550
rect 52738 50504 52790 50550
rect 52948 50504 53000 50550
rect 53159 50504 53211 50550
rect 53371 50504 53423 50550
rect 53582 50504 53634 50550
rect 50557 50501 50609 50504
rect 50768 50501 50820 50504
rect 39775 50280 39786 50315
rect 39786 50280 39827 50315
rect 39775 50263 39827 50280
rect 39994 50048 40046 50100
rect 39994 49862 40046 49914
rect 52316 50501 52368 50504
rect 52527 50501 52579 50504
rect 52738 50501 52790 50504
rect 52948 50501 53000 50504
rect 53159 50501 53211 50504
rect 53371 50501 53423 50504
rect 53582 50501 53634 50504
rect 53792 50501 53844 50553
rect 54003 50501 54055 50553
rect 54214 50501 54266 50553
rect 54855 50501 54907 50553
rect 55066 50501 55118 50553
rect 55278 50550 55330 50553
rect 55278 50504 55279 50550
rect 55279 50504 55325 50550
rect 55325 50504 55330 50550
rect 55278 50501 55330 50504
rect 55489 50501 55541 50553
rect 41935 50263 41987 50315
rect 51073 50326 51125 50329
rect 51253 50326 51305 50329
rect 43068 50032 43120 50084
rect 51073 50280 51086 50326
rect 51086 50280 51125 50326
rect 51253 50280 51292 50326
rect 51292 50280 51305 50326
rect 48943 50239 48995 50254
rect 49154 50239 49206 50254
rect 49365 50239 49417 50254
rect 49576 50239 49628 50254
rect 49787 50239 49839 50254
rect 48943 50202 48984 50239
rect 48984 50202 48995 50239
rect 49154 50202 49190 50239
rect 49190 50202 49206 50239
rect 49365 50202 49396 50239
rect 49396 50202 49417 50239
rect 49576 50202 49602 50239
rect 49602 50202 49628 50239
rect 49787 50202 49839 50239
rect 51073 50277 51125 50280
rect 51253 50277 51305 50280
rect 44939 50056 44971 50091
rect 44971 50056 44991 50091
rect 45151 50056 45197 50091
rect 45197 50056 45203 50091
rect 48596 50095 48648 50147
rect 44939 50039 44991 50056
rect 45151 50039 45203 50056
rect 45597 49937 45604 49975
rect 45604 49937 45649 49975
rect 45597 49923 45649 49937
rect 50300 50039 50352 50091
rect 50511 50056 50513 50091
rect 50513 50056 50563 50091
rect 50511 50039 50563 50056
rect 50722 50039 50774 50091
rect 48596 49877 48648 49929
rect 51835 50280 51887 50322
rect 52015 50280 52067 50322
rect 51835 50270 51887 50280
rect 52015 50270 52067 50280
rect 35332 49745 35384 49791
rect 35543 49745 35580 49791
rect 35580 49745 35595 49791
rect 35754 49745 35786 49791
rect 35786 49745 35806 49791
rect 35965 49745 35992 49791
rect 35992 49745 36017 49791
rect 36176 49745 36198 49791
rect 36198 49745 36228 49791
rect 37891 49745 37909 49789
rect 37909 49745 37943 49789
rect 38071 49745 38072 49789
rect 38072 49745 38123 49789
rect 48943 49745 48984 49791
rect 48984 49745 48995 49791
rect 49154 49745 49190 49791
rect 49190 49745 49206 49791
rect 49365 49745 49396 49791
rect 49396 49745 49417 49791
rect 49576 49745 49602 49791
rect 49602 49745 49628 49791
rect 49787 49745 49839 49791
rect 51835 49832 51887 49859
rect 52015 49832 52067 49859
rect 51835 49807 51887 49832
rect 52015 49807 52067 49832
rect 35332 49739 35384 49745
rect 35543 49739 35595 49745
rect 35754 49739 35806 49745
rect 35965 49739 36017 49745
rect 36176 49739 36228 49745
rect 37891 49737 37943 49745
rect 38071 49737 38123 49745
rect 27790 49601 27842 49653
rect 28001 49601 28053 49653
rect 28212 49601 28264 49653
rect 28423 49601 28475 49653
rect 28634 49601 28686 49653
rect 28845 49650 28897 49653
rect 28845 49604 28856 49650
rect 28856 49604 28897 49650
rect 28845 49601 28897 49604
rect 29056 49601 29108 49653
rect 29582 49601 29634 49653
rect 29793 49650 29845 49653
rect 29793 49604 29798 49650
rect 29798 49604 29844 49650
rect 29844 49604 29845 49650
rect 29793 49601 29845 49604
rect 30005 49601 30057 49653
rect 30216 49601 30268 49653
rect 30854 49601 30906 49653
rect 31065 49601 31117 49653
rect 31276 49601 31328 49653
rect 31486 49601 31538 49653
rect 31697 49601 31749 49653
rect 31909 49601 31961 49653
rect 32120 49601 32172 49653
rect 32330 49601 32382 49653
rect 32541 49601 32593 49653
rect 32752 49601 32804 49653
rect 48943 49739 48995 49745
rect 49154 49739 49206 49745
rect 49365 49739 49417 49745
rect 49576 49739 49628 49745
rect 49787 49739 49839 49745
rect 34755 49601 34807 49653
rect 34935 49650 34987 49653
rect 34935 49604 34962 49650
rect 34962 49604 34987 49650
rect 34935 49601 34987 49604
rect 50138 49650 50190 49653
rect 50138 49604 50160 49650
rect 50160 49604 50190 49650
rect 50138 49601 50190 49604
rect 50318 49601 50370 49653
rect 35332 49509 35384 49515
rect 35543 49509 35595 49515
rect 35754 49509 35806 49515
rect 35965 49509 36017 49515
rect 36176 49509 36228 49515
rect 37891 49509 37943 49517
rect 38071 49509 38123 49517
rect 52316 49601 52368 49653
rect 52527 49601 52579 49653
rect 52738 49601 52790 49653
rect 52948 49601 53000 49653
rect 53159 49601 53211 49653
rect 53371 49601 53423 49653
rect 53582 49601 53634 49653
rect 53792 49601 53844 49653
rect 54003 49601 54055 49653
rect 54214 49601 54266 49653
rect 54855 49601 54907 49653
rect 55066 49601 55118 49653
rect 55278 49650 55330 49653
rect 55278 49604 55279 49650
rect 55279 49604 55325 49650
rect 55325 49604 55330 49650
rect 55278 49601 55330 49604
rect 55489 49601 55541 49653
rect 56015 49601 56067 49653
rect 56226 49650 56278 49653
rect 56226 49604 56267 49650
rect 56267 49604 56278 49650
rect 56226 49601 56278 49604
rect 56437 49601 56489 49653
rect 56648 49601 56700 49653
rect 56859 49601 56911 49653
rect 57070 49601 57122 49653
rect 57281 49601 57333 49653
rect 48943 49509 48995 49515
rect 49154 49509 49206 49515
rect 49365 49509 49417 49515
rect 49576 49509 49628 49515
rect 49787 49509 49839 49515
rect 33057 49422 33109 49425
rect 33237 49422 33289 49425
rect 35332 49463 35384 49509
rect 35543 49463 35580 49509
rect 35580 49463 35595 49509
rect 35754 49463 35786 49509
rect 35786 49463 35806 49509
rect 35965 49463 35992 49509
rect 35992 49463 36017 49509
rect 36176 49463 36198 49509
rect 36198 49463 36228 49509
rect 37891 49465 37909 49509
rect 37909 49465 37943 49509
rect 38071 49465 38072 49509
rect 38072 49465 38123 49509
rect 33057 49376 33109 49422
rect 33237 49376 33289 49422
rect 33057 49373 33109 49376
rect 33237 49373 33289 49376
rect 33057 48974 33109 48977
rect 33237 48974 33289 48977
rect 33057 48928 33109 48974
rect 33237 48928 33289 48974
rect 33057 48925 33109 48928
rect 33237 48925 33289 48928
rect 29582 48701 29634 48753
rect 29793 48750 29845 48753
rect 29793 48704 29798 48750
rect 29798 48704 29844 48750
rect 29844 48704 29845 48750
rect 29793 48701 29845 48704
rect 30005 48701 30057 48753
rect 30216 48701 30268 48753
rect 34267 49198 34319 49215
rect 34447 49198 34499 49215
rect 34627 49198 34679 49215
rect 34267 49163 34302 49198
rect 34302 49163 34319 49198
rect 34447 49163 34451 49198
rect 34451 49163 34499 49198
rect 34627 49163 34658 49198
rect 34658 49163 34679 49198
rect 36678 49238 36697 49290
rect 36697 49238 36730 49290
rect 48943 49463 48984 49509
rect 48984 49463 48995 49509
rect 49154 49463 49190 49509
rect 49190 49463 49206 49509
rect 49365 49463 49396 49509
rect 49396 49463 49417 49509
rect 49576 49463 49602 49509
rect 49602 49463 49628 49509
rect 49787 49463 49839 49509
rect 39994 49340 40046 49392
rect 36961 49239 36971 49283
rect 36971 49239 37013 49283
rect 37172 49239 37206 49283
rect 37206 49239 37224 49283
rect 36961 49231 37013 49239
rect 37172 49231 37224 49239
rect 37384 49231 37436 49283
rect 37595 49231 37647 49283
rect 35332 49015 35384 49055
rect 35543 49015 35580 49055
rect 35580 49015 35595 49055
rect 35754 49015 35786 49055
rect 35786 49015 35806 49055
rect 35965 49015 35992 49055
rect 35992 49015 36017 49055
rect 36176 49015 36198 49055
rect 36198 49015 36228 49055
rect 37891 49015 37909 49043
rect 37909 49015 37943 49043
rect 38071 49015 38072 49043
rect 38072 49015 38123 49043
rect 35332 49003 35384 49015
rect 35543 49003 35595 49015
rect 35754 49003 35806 49015
rect 35965 49003 36017 49015
rect 36176 49003 36228 49015
rect 33819 48928 33833 48969
rect 33833 48928 33871 48969
rect 33999 48928 34039 48969
rect 34039 48928 34051 48969
rect 37891 48991 37943 49015
rect 38071 48991 38123 49015
rect 33819 48917 33871 48928
rect 33999 48917 34051 48928
rect 30854 48701 30906 48753
rect 31065 48701 31117 48753
rect 31276 48701 31328 48753
rect 31486 48750 31538 48753
rect 31697 48750 31749 48753
rect 31909 48750 31961 48753
rect 32120 48750 32172 48753
rect 32330 48750 32382 48753
rect 32541 48750 32593 48753
rect 32752 48750 32804 48753
rect 34284 48750 34336 48753
rect 34495 48750 34547 48753
rect 31486 48704 31538 48750
rect 31697 48704 31749 48750
rect 31909 48704 31961 48750
rect 32120 48704 32172 48750
rect 32330 48704 32382 48750
rect 32541 48704 32593 48750
rect 32752 48704 32804 48750
rect 34284 48704 34302 48750
rect 34302 48704 34336 48750
rect 34495 48704 34508 48750
rect 34508 48704 34547 48750
rect 31486 48701 31538 48704
rect 31697 48701 31749 48704
rect 31909 48701 31961 48704
rect 32120 48701 32172 48704
rect 32330 48701 32382 48704
rect 32541 48701 32593 48704
rect 32752 48701 32804 48704
rect 34284 48701 34336 48704
rect 34495 48701 34547 48704
rect 34707 48701 34759 48753
rect 34918 48701 34970 48753
rect 35220 48701 35272 48753
rect 35430 48701 35482 48753
rect 35641 48701 35693 48753
rect 35853 48701 35905 48753
rect 36064 48701 36116 48753
rect 36274 48701 36326 48753
rect 38330 48750 38382 48753
rect 38330 48704 38382 48750
rect 38330 48701 38382 48704
rect 38541 48701 38593 48753
rect 38752 48701 38804 48753
rect 39052 48750 39104 48753
rect 39232 48750 39284 48753
rect 39052 48704 39062 48750
rect 39062 48704 39104 48750
rect 39232 48704 39266 48750
rect 39266 48704 39284 48750
rect 39052 48701 39104 48704
rect 39232 48701 39284 48704
rect 33057 48526 33109 48529
rect 33237 48526 33289 48529
rect 33057 48480 33109 48526
rect 33237 48480 33289 48526
rect 33057 48477 33109 48480
rect 33237 48477 33289 48480
rect 33819 48526 33871 48537
rect 33999 48526 34051 48537
rect 33819 48485 33833 48526
rect 33833 48485 33871 48526
rect 33999 48485 34039 48526
rect 34039 48485 34051 48526
rect 35332 48439 35384 48451
rect 35543 48439 35595 48451
rect 35754 48439 35806 48451
rect 35965 48439 36017 48451
rect 36176 48439 36228 48451
rect 37891 48439 37943 48463
rect 38071 48439 38123 48463
rect 35332 48399 35384 48439
rect 35543 48399 35580 48439
rect 35580 48399 35595 48439
rect 35754 48399 35786 48439
rect 35786 48399 35806 48439
rect 35965 48399 35992 48439
rect 35992 48399 36017 48439
rect 36176 48399 36198 48439
rect 36198 48399 36228 48439
rect 37891 48411 37909 48439
rect 37909 48411 37943 48439
rect 38071 48411 38072 48439
rect 38072 48411 38123 48439
rect 34267 48256 34302 48291
rect 34302 48256 34319 48291
rect 34447 48256 34451 48291
rect 34451 48256 34499 48291
rect 34627 48256 34658 48291
rect 34658 48256 34679 48291
rect 34267 48239 34319 48256
rect 34447 48239 34499 48256
rect 34627 48239 34679 48256
rect 33057 48078 33109 48081
rect 33237 48078 33289 48081
rect 33057 48032 33109 48078
rect 33237 48032 33289 48078
rect 33057 48029 33109 48032
rect 33237 48029 33289 48032
rect 36678 48164 36697 48216
rect 36697 48164 36730 48216
rect 36961 48215 37013 48223
rect 37172 48215 37224 48223
rect 36961 48171 36971 48215
rect 36971 48171 37013 48215
rect 37172 48171 37206 48215
rect 37206 48171 37224 48215
rect 37384 48171 37436 48223
rect 37595 48171 37647 48223
rect 39994 49154 40046 49206
rect 39775 48974 39827 48991
rect 39775 48939 39786 48974
rect 39786 48939 39827 48974
rect 43068 49170 43120 49222
rect 41935 48939 41987 48991
rect 45975 49279 46027 49331
rect 48596 49325 48648 49377
rect 51835 49422 51887 49447
rect 52015 49422 52067 49447
rect 51835 49395 51887 49422
rect 52015 49395 52067 49422
rect 44939 49198 44991 49215
rect 45151 49198 45203 49215
rect 44939 49163 44971 49198
rect 44971 49163 44991 49198
rect 45151 49163 45197 49198
rect 45197 49163 45203 49198
rect 48596 49107 48648 49159
rect 50300 49163 50352 49215
rect 50511 49198 50563 49215
rect 50511 49163 50513 49198
rect 50513 49163 50563 49198
rect 50722 49163 50774 49215
rect 48943 49015 48984 49052
rect 48984 49015 48995 49052
rect 49154 49015 49190 49052
rect 49190 49015 49206 49052
rect 49365 49015 49396 49052
rect 49396 49015 49417 49052
rect 49576 49015 49602 49052
rect 49602 49015 49628 49052
rect 49787 49015 49839 49052
rect 48943 49000 48995 49015
rect 49154 49000 49206 49015
rect 49365 49000 49417 49015
rect 49576 49000 49628 49015
rect 49787 49000 49839 49015
rect 51073 48974 51125 48977
rect 51253 48974 51305 48977
rect 51073 48928 51086 48974
rect 51086 48928 51125 48974
rect 51253 48928 51292 48974
rect 51292 48928 51305 48974
rect 51073 48925 51125 48928
rect 51253 48925 51305 48928
rect 51835 48974 51887 48984
rect 52015 48974 52067 48984
rect 51835 48932 51887 48974
rect 52015 48932 52067 48974
rect 40253 48701 40305 48753
rect 40433 48701 40485 48753
rect 43790 48701 43842 48753
rect 44001 48701 44053 48753
rect 44213 48750 44265 48753
rect 44213 48704 44236 48750
rect 44236 48704 44265 48750
rect 44213 48701 44265 48704
rect 44424 48701 44476 48753
rect 44834 48750 44886 48753
rect 45045 48750 45097 48753
rect 45256 48750 45308 48753
rect 44834 48704 44858 48750
rect 44858 48704 44886 48750
rect 45045 48704 45084 48750
rect 45084 48704 45097 48750
rect 45256 48704 45264 48750
rect 45264 48704 45308 48750
rect 44834 48701 44886 48704
rect 45045 48701 45097 48704
rect 45256 48701 45308 48704
rect 48838 48701 48890 48753
rect 49048 48701 49100 48753
rect 49259 48701 49311 48753
rect 49471 48701 49523 48753
rect 49682 48701 49734 48753
rect 49892 48701 49944 48753
rect 50346 48701 50398 48753
rect 50557 48750 50609 48753
rect 50768 48750 50820 48753
rect 52316 48750 52368 48753
rect 52527 48750 52579 48753
rect 52738 48750 52790 48753
rect 52948 48750 53000 48753
rect 53159 48750 53211 48753
rect 53371 48750 53423 48753
rect 53582 48750 53634 48753
rect 50557 48704 50571 48750
rect 50571 48704 50609 48750
rect 50768 48704 50777 48750
rect 50777 48704 50820 48750
rect 52316 48704 52368 48750
rect 52527 48704 52579 48750
rect 52738 48704 52790 48750
rect 52948 48704 53000 48750
rect 53159 48704 53211 48750
rect 53371 48704 53423 48750
rect 53582 48704 53634 48750
rect 50557 48701 50609 48704
rect 50768 48701 50820 48704
rect 39775 48480 39786 48515
rect 39786 48480 39827 48515
rect 39775 48463 39827 48480
rect 39994 48248 40046 48300
rect 39994 48062 40046 48114
rect 52316 48701 52368 48704
rect 52527 48701 52579 48704
rect 52738 48701 52790 48704
rect 52948 48701 53000 48704
rect 53159 48701 53211 48704
rect 53371 48701 53423 48704
rect 53582 48701 53634 48704
rect 53792 48701 53844 48753
rect 54003 48701 54055 48753
rect 54214 48701 54266 48753
rect 54855 48701 54907 48753
rect 55066 48701 55118 48753
rect 55278 48750 55330 48753
rect 55278 48704 55279 48750
rect 55279 48704 55325 48750
rect 55325 48704 55330 48750
rect 55278 48701 55330 48704
rect 55489 48701 55541 48753
rect 41935 48463 41987 48515
rect 51073 48526 51125 48529
rect 51253 48526 51305 48529
rect 43068 48232 43120 48284
rect 51073 48480 51086 48526
rect 51086 48480 51125 48526
rect 51253 48480 51292 48526
rect 51292 48480 51305 48526
rect 48943 48439 48995 48454
rect 49154 48439 49206 48454
rect 49365 48439 49417 48454
rect 49576 48439 49628 48454
rect 49787 48439 49839 48454
rect 48943 48402 48984 48439
rect 48984 48402 48995 48439
rect 49154 48402 49190 48439
rect 49190 48402 49206 48439
rect 49365 48402 49396 48439
rect 49396 48402 49417 48439
rect 49576 48402 49602 48439
rect 49602 48402 49628 48439
rect 49787 48402 49839 48439
rect 51073 48477 51125 48480
rect 51253 48477 51305 48480
rect 44939 48256 44971 48291
rect 44971 48256 44991 48291
rect 45151 48256 45197 48291
rect 45197 48256 45203 48291
rect 48596 48295 48648 48347
rect 44939 48239 44991 48256
rect 45151 48239 45203 48256
rect 46353 48123 46405 48175
rect 50300 48239 50352 48291
rect 50511 48256 50513 48291
rect 50513 48256 50563 48291
rect 50511 48239 50563 48256
rect 50722 48239 50774 48291
rect 48596 48077 48648 48129
rect 51835 48480 51887 48522
rect 52015 48480 52067 48522
rect 51835 48470 51887 48480
rect 52015 48470 52067 48480
rect 35332 47945 35384 47991
rect 35543 47945 35580 47991
rect 35580 47945 35595 47991
rect 35754 47945 35786 47991
rect 35786 47945 35806 47991
rect 35965 47945 35992 47991
rect 35992 47945 36017 47991
rect 36176 47945 36198 47991
rect 36198 47945 36228 47991
rect 37891 47945 37909 47989
rect 37909 47945 37943 47989
rect 38071 47945 38072 47989
rect 38072 47945 38123 47989
rect 48943 47945 48984 47991
rect 48984 47945 48995 47991
rect 49154 47945 49190 47991
rect 49190 47945 49206 47991
rect 49365 47945 49396 47991
rect 49396 47945 49417 47991
rect 49576 47945 49602 47991
rect 49602 47945 49628 47991
rect 49787 47945 49839 47991
rect 51835 48032 51887 48059
rect 52015 48032 52067 48059
rect 51835 48007 51887 48032
rect 52015 48007 52067 48032
rect 35332 47939 35384 47945
rect 35543 47939 35595 47945
rect 35754 47939 35806 47945
rect 35965 47939 36017 47945
rect 36176 47939 36228 47945
rect 37891 47937 37943 47945
rect 38071 47937 38123 47945
rect 27790 47801 27842 47853
rect 28001 47801 28053 47853
rect 28212 47801 28264 47853
rect 28423 47801 28475 47853
rect 28634 47801 28686 47853
rect 28845 47850 28897 47853
rect 28845 47804 28856 47850
rect 28856 47804 28897 47850
rect 28845 47801 28897 47804
rect 29056 47801 29108 47853
rect 29582 47801 29634 47853
rect 29793 47850 29845 47853
rect 29793 47804 29798 47850
rect 29798 47804 29844 47850
rect 29844 47804 29845 47850
rect 29793 47801 29845 47804
rect 30005 47801 30057 47853
rect 30216 47801 30268 47853
rect 30854 47801 30906 47853
rect 31065 47801 31117 47853
rect 31276 47801 31328 47853
rect 31486 47801 31538 47853
rect 31697 47801 31749 47853
rect 31909 47801 31961 47853
rect 32120 47801 32172 47853
rect 32330 47801 32382 47853
rect 32541 47801 32593 47853
rect 32752 47801 32804 47853
rect 48943 47939 48995 47945
rect 49154 47939 49206 47945
rect 49365 47939 49417 47945
rect 49576 47939 49628 47945
rect 49787 47939 49839 47945
rect 34755 47801 34807 47853
rect 34935 47850 34987 47853
rect 34935 47804 34962 47850
rect 34962 47804 34987 47850
rect 34935 47801 34987 47804
rect 50138 47850 50190 47853
rect 50138 47804 50160 47850
rect 50160 47804 50190 47850
rect 50138 47801 50190 47804
rect 50318 47801 50370 47853
rect 35332 47709 35384 47715
rect 35543 47709 35595 47715
rect 35754 47709 35806 47715
rect 35965 47709 36017 47715
rect 36176 47709 36228 47715
rect 37891 47709 37943 47717
rect 38071 47709 38123 47717
rect 52316 47801 52368 47853
rect 52527 47801 52579 47853
rect 52738 47801 52790 47853
rect 52948 47801 53000 47853
rect 53159 47801 53211 47853
rect 53371 47801 53423 47853
rect 53582 47801 53634 47853
rect 53792 47801 53844 47853
rect 54003 47801 54055 47853
rect 54214 47801 54266 47853
rect 54855 47801 54907 47853
rect 55066 47801 55118 47853
rect 55278 47850 55330 47853
rect 55278 47804 55279 47850
rect 55279 47804 55325 47850
rect 55325 47804 55330 47850
rect 55278 47801 55330 47804
rect 55489 47801 55541 47853
rect 56015 47801 56067 47853
rect 56226 47850 56278 47853
rect 56226 47804 56267 47850
rect 56267 47804 56278 47850
rect 56226 47801 56278 47804
rect 56437 47801 56489 47853
rect 56648 47801 56700 47853
rect 56859 47801 56911 47853
rect 57070 47801 57122 47853
rect 57281 47801 57333 47853
rect 48943 47709 48995 47715
rect 49154 47709 49206 47715
rect 49365 47709 49417 47715
rect 49576 47709 49628 47715
rect 49787 47709 49839 47715
rect 33057 47622 33109 47625
rect 33237 47622 33289 47625
rect 35332 47663 35384 47709
rect 35543 47663 35580 47709
rect 35580 47663 35595 47709
rect 35754 47663 35786 47709
rect 35786 47663 35806 47709
rect 35965 47663 35992 47709
rect 35992 47663 36017 47709
rect 36176 47663 36198 47709
rect 36198 47663 36228 47709
rect 37891 47665 37909 47709
rect 37909 47665 37943 47709
rect 38071 47665 38072 47709
rect 38072 47665 38123 47709
rect 33057 47576 33109 47622
rect 33237 47576 33289 47622
rect 33057 47573 33109 47576
rect 33237 47573 33289 47576
rect 33057 47174 33109 47177
rect 33237 47174 33289 47177
rect 33057 47128 33109 47174
rect 33237 47128 33289 47174
rect 33057 47125 33109 47128
rect 33237 47125 33289 47128
rect 29582 46901 29634 46953
rect 29793 46950 29845 46953
rect 29793 46904 29798 46950
rect 29798 46904 29844 46950
rect 29844 46904 29845 46950
rect 29793 46901 29845 46904
rect 30005 46901 30057 46953
rect 30216 46901 30268 46953
rect 34267 47398 34319 47415
rect 34447 47398 34499 47415
rect 34627 47398 34679 47415
rect 34267 47363 34302 47398
rect 34302 47363 34319 47398
rect 34447 47363 34451 47398
rect 34451 47363 34499 47398
rect 34627 47363 34658 47398
rect 34658 47363 34679 47398
rect 36678 47438 36697 47490
rect 36697 47438 36730 47490
rect 48943 47663 48984 47709
rect 48984 47663 48995 47709
rect 49154 47663 49190 47709
rect 49190 47663 49206 47709
rect 49365 47663 49396 47709
rect 49396 47663 49417 47709
rect 49576 47663 49602 47709
rect 49602 47663 49628 47709
rect 49787 47663 49839 47709
rect 39994 47540 40046 47592
rect 36961 47439 36971 47483
rect 36971 47439 37013 47483
rect 37172 47439 37206 47483
rect 37206 47439 37224 47483
rect 36961 47431 37013 47439
rect 37172 47431 37224 47439
rect 37384 47431 37436 47483
rect 37595 47431 37647 47483
rect 35332 47215 35384 47255
rect 35543 47215 35580 47255
rect 35580 47215 35595 47255
rect 35754 47215 35786 47255
rect 35786 47215 35806 47255
rect 35965 47215 35992 47255
rect 35992 47215 36017 47255
rect 36176 47215 36198 47255
rect 36198 47215 36228 47255
rect 37891 47215 37909 47243
rect 37909 47215 37943 47243
rect 38071 47215 38072 47243
rect 38072 47215 38123 47243
rect 35332 47203 35384 47215
rect 35543 47203 35595 47215
rect 35754 47203 35806 47215
rect 35965 47203 36017 47215
rect 36176 47203 36228 47215
rect 33819 47128 33833 47169
rect 33833 47128 33871 47169
rect 33999 47128 34039 47169
rect 34039 47128 34051 47169
rect 37891 47191 37943 47215
rect 38071 47191 38123 47215
rect 33819 47117 33871 47128
rect 33999 47117 34051 47128
rect 30854 46901 30906 46953
rect 31065 46901 31117 46953
rect 31276 46901 31328 46953
rect 31486 46950 31538 46953
rect 31697 46950 31749 46953
rect 31909 46950 31961 46953
rect 32120 46950 32172 46953
rect 32330 46950 32382 46953
rect 32541 46950 32593 46953
rect 32752 46950 32804 46953
rect 34284 46950 34336 46953
rect 34495 46950 34547 46953
rect 31486 46904 31538 46950
rect 31697 46904 31749 46950
rect 31909 46904 31961 46950
rect 32120 46904 32172 46950
rect 32330 46904 32382 46950
rect 32541 46904 32593 46950
rect 32752 46904 32804 46950
rect 34284 46904 34302 46950
rect 34302 46904 34336 46950
rect 34495 46904 34508 46950
rect 34508 46904 34547 46950
rect 31486 46901 31538 46904
rect 31697 46901 31749 46904
rect 31909 46901 31961 46904
rect 32120 46901 32172 46904
rect 32330 46901 32382 46904
rect 32541 46901 32593 46904
rect 32752 46901 32804 46904
rect 34284 46901 34336 46904
rect 34495 46901 34547 46904
rect 34707 46901 34759 46953
rect 34918 46901 34970 46953
rect 35220 46901 35272 46953
rect 35430 46901 35482 46953
rect 35641 46901 35693 46953
rect 35853 46901 35905 46953
rect 36064 46901 36116 46953
rect 36274 46901 36326 46953
rect 38330 46950 38382 46953
rect 38330 46904 38382 46950
rect 38330 46901 38382 46904
rect 38541 46901 38593 46953
rect 38752 46901 38804 46953
rect 39052 46950 39104 46953
rect 39232 46950 39284 46953
rect 39052 46904 39062 46950
rect 39062 46904 39104 46950
rect 39232 46904 39266 46950
rect 39266 46904 39284 46950
rect 39052 46901 39104 46904
rect 39232 46901 39284 46904
rect 33057 46726 33109 46729
rect 33237 46726 33289 46729
rect 33057 46680 33109 46726
rect 33237 46680 33289 46726
rect 33057 46677 33109 46680
rect 33237 46677 33289 46680
rect 33819 46726 33871 46737
rect 33999 46726 34051 46737
rect 33819 46685 33833 46726
rect 33833 46685 33871 46726
rect 33999 46685 34039 46726
rect 34039 46685 34051 46726
rect 35332 46639 35384 46651
rect 35543 46639 35595 46651
rect 35754 46639 35806 46651
rect 35965 46639 36017 46651
rect 36176 46639 36228 46651
rect 37891 46639 37943 46663
rect 38071 46639 38123 46663
rect 35332 46599 35384 46639
rect 35543 46599 35580 46639
rect 35580 46599 35595 46639
rect 35754 46599 35786 46639
rect 35786 46599 35806 46639
rect 35965 46599 35992 46639
rect 35992 46599 36017 46639
rect 36176 46599 36198 46639
rect 36198 46599 36228 46639
rect 37891 46611 37909 46639
rect 37909 46611 37943 46639
rect 38071 46611 38072 46639
rect 38072 46611 38123 46639
rect 34267 46456 34302 46491
rect 34302 46456 34319 46491
rect 34447 46456 34451 46491
rect 34451 46456 34499 46491
rect 34627 46456 34658 46491
rect 34658 46456 34679 46491
rect 34267 46439 34319 46456
rect 34447 46439 34499 46456
rect 34627 46439 34679 46456
rect 33057 46278 33109 46281
rect 33237 46278 33289 46281
rect 33057 46232 33109 46278
rect 33237 46232 33289 46278
rect 33057 46229 33109 46232
rect 33237 46229 33289 46232
rect 36678 46364 36697 46416
rect 36697 46364 36730 46416
rect 36961 46415 37013 46423
rect 37172 46415 37224 46423
rect 36961 46371 36971 46415
rect 36971 46371 37013 46415
rect 37172 46371 37206 46415
rect 37206 46371 37224 46415
rect 37384 46371 37436 46423
rect 37595 46371 37647 46423
rect 39994 47354 40046 47406
rect 39775 47174 39827 47191
rect 39775 47139 39786 47174
rect 39786 47139 39827 47174
rect 43068 47370 43120 47422
rect 41935 47139 41987 47191
rect 46731 47479 46783 47531
rect 48596 47525 48648 47577
rect 51835 47622 51887 47647
rect 52015 47622 52067 47647
rect 51835 47595 51887 47622
rect 52015 47595 52067 47622
rect 44939 47398 44991 47415
rect 45151 47398 45203 47415
rect 44939 47363 44971 47398
rect 44971 47363 44991 47398
rect 45151 47363 45197 47398
rect 45197 47363 45203 47398
rect 48596 47307 48648 47359
rect 50300 47363 50352 47415
rect 50511 47398 50563 47415
rect 50511 47363 50513 47398
rect 50513 47363 50563 47398
rect 50722 47363 50774 47415
rect 48943 47215 48984 47252
rect 48984 47215 48995 47252
rect 49154 47215 49190 47252
rect 49190 47215 49206 47252
rect 49365 47215 49396 47252
rect 49396 47215 49417 47252
rect 49576 47215 49602 47252
rect 49602 47215 49628 47252
rect 49787 47215 49839 47252
rect 48943 47200 48995 47215
rect 49154 47200 49206 47215
rect 49365 47200 49417 47215
rect 49576 47200 49628 47215
rect 49787 47200 49839 47215
rect 51073 47174 51125 47177
rect 51253 47174 51305 47177
rect 51073 47128 51086 47174
rect 51086 47128 51125 47174
rect 51253 47128 51292 47174
rect 51292 47128 51305 47174
rect 51073 47125 51125 47128
rect 51253 47125 51305 47128
rect 51835 47174 51887 47184
rect 52015 47174 52067 47184
rect 51835 47132 51887 47174
rect 52015 47132 52067 47174
rect 40253 46901 40305 46953
rect 40433 46901 40485 46953
rect 43790 46901 43842 46953
rect 44001 46901 44053 46953
rect 44213 46950 44265 46953
rect 44213 46904 44236 46950
rect 44236 46904 44265 46950
rect 44213 46901 44265 46904
rect 44424 46901 44476 46953
rect 44834 46950 44886 46953
rect 45045 46950 45097 46953
rect 45256 46950 45308 46953
rect 44834 46904 44858 46950
rect 44858 46904 44886 46950
rect 45045 46904 45084 46950
rect 45084 46904 45097 46950
rect 45256 46904 45264 46950
rect 45264 46904 45308 46950
rect 44834 46901 44886 46904
rect 45045 46901 45097 46904
rect 45256 46901 45308 46904
rect 48838 46901 48890 46953
rect 49048 46901 49100 46953
rect 49259 46901 49311 46953
rect 49471 46901 49523 46953
rect 49682 46901 49734 46953
rect 49892 46901 49944 46953
rect 50346 46901 50398 46953
rect 50557 46950 50609 46953
rect 50768 46950 50820 46953
rect 52316 46950 52368 46953
rect 52527 46950 52579 46953
rect 52738 46950 52790 46953
rect 52948 46950 53000 46953
rect 53159 46950 53211 46953
rect 53371 46950 53423 46953
rect 53582 46950 53634 46953
rect 50557 46904 50571 46950
rect 50571 46904 50609 46950
rect 50768 46904 50777 46950
rect 50777 46904 50820 46950
rect 52316 46904 52368 46950
rect 52527 46904 52579 46950
rect 52738 46904 52790 46950
rect 52948 46904 53000 46950
rect 53159 46904 53211 46950
rect 53371 46904 53423 46950
rect 53582 46904 53634 46950
rect 50557 46901 50609 46904
rect 50768 46901 50820 46904
rect 39775 46680 39786 46715
rect 39786 46680 39827 46715
rect 39775 46663 39827 46680
rect 39994 46448 40046 46500
rect 39994 46262 40046 46314
rect 52316 46901 52368 46904
rect 52527 46901 52579 46904
rect 52738 46901 52790 46904
rect 52948 46901 53000 46904
rect 53159 46901 53211 46904
rect 53371 46901 53423 46904
rect 53582 46901 53634 46904
rect 53792 46901 53844 46953
rect 54003 46901 54055 46953
rect 54214 46901 54266 46953
rect 54855 46901 54907 46953
rect 55066 46901 55118 46953
rect 55278 46950 55330 46953
rect 55278 46904 55279 46950
rect 55279 46904 55325 46950
rect 55325 46904 55330 46950
rect 55278 46901 55330 46904
rect 55489 46901 55541 46953
rect 41935 46663 41987 46715
rect 51073 46726 51125 46729
rect 51253 46726 51305 46729
rect 43068 46432 43120 46484
rect 51073 46680 51086 46726
rect 51086 46680 51125 46726
rect 51253 46680 51292 46726
rect 51292 46680 51305 46726
rect 48943 46639 48995 46654
rect 49154 46639 49206 46654
rect 49365 46639 49417 46654
rect 49576 46639 49628 46654
rect 49787 46639 49839 46654
rect 48943 46602 48984 46639
rect 48984 46602 48995 46639
rect 49154 46602 49190 46639
rect 49190 46602 49206 46639
rect 49365 46602 49396 46639
rect 49396 46602 49417 46639
rect 49576 46602 49602 46639
rect 49602 46602 49628 46639
rect 49787 46602 49839 46639
rect 51073 46677 51125 46680
rect 51253 46677 51305 46680
rect 44939 46456 44971 46491
rect 44971 46456 44991 46491
rect 45151 46456 45197 46491
rect 45197 46456 45203 46491
rect 48596 46495 48648 46547
rect 44939 46439 44991 46456
rect 45151 46439 45203 46456
rect 47108 46323 47160 46375
rect 50300 46439 50352 46491
rect 50511 46456 50513 46491
rect 50513 46456 50563 46491
rect 50511 46439 50563 46456
rect 50722 46439 50774 46491
rect 48596 46277 48648 46329
rect 51835 46680 51887 46722
rect 52015 46680 52067 46722
rect 51835 46670 51887 46680
rect 52015 46670 52067 46680
rect 35332 46145 35384 46191
rect 35543 46145 35580 46191
rect 35580 46145 35595 46191
rect 35754 46145 35786 46191
rect 35786 46145 35806 46191
rect 35965 46145 35992 46191
rect 35992 46145 36017 46191
rect 36176 46145 36198 46191
rect 36198 46145 36228 46191
rect 37891 46145 37909 46189
rect 37909 46145 37943 46189
rect 38071 46145 38072 46189
rect 38072 46145 38123 46189
rect 48943 46145 48984 46191
rect 48984 46145 48995 46191
rect 49154 46145 49190 46191
rect 49190 46145 49206 46191
rect 49365 46145 49396 46191
rect 49396 46145 49417 46191
rect 49576 46145 49602 46191
rect 49602 46145 49628 46191
rect 49787 46145 49839 46191
rect 51835 46232 51887 46259
rect 52015 46232 52067 46259
rect 51835 46207 51887 46232
rect 52015 46207 52067 46232
rect 35332 46139 35384 46145
rect 35543 46139 35595 46145
rect 35754 46139 35806 46145
rect 35965 46139 36017 46145
rect 36176 46139 36228 46145
rect 37891 46137 37943 46145
rect 38071 46137 38123 46145
rect 27790 46001 27842 46053
rect 28001 46001 28053 46053
rect 28212 46001 28264 46053
rect 28423 46001 28475 46053
rect 28634 46001 28686 46053
rect 28845 46050 28897 46053
rect 28845 46004 28856 46050
rect 28856 46004 28897 46050
rect 28845 46001 28897 46004
rect 29056 46001 29108 46053
rect 29582 46001 29634 46053
rect 29793 46050 29845 46053
rect 29793 46004 29798 46050
rect 29798 46004 29844 46050
rect 29844 46004 29845 46050
rect 29793 46001 29845 46004
rect 30005 46001 30057 46053
rect 30216 46001 30268 46053
rect 30854 46001 30906 46053
rect 31065 46001 31117 46053
rect 31276 46001 31328 46053
rect 31486 46001 31538 46053
rect 31697 46001 31749 46053
rect 31909 46001 31961 46053
rect 32120 46001 32172 46053
rect 32330 46001 32382 46053
rect 32541 46001 32593 46053
rect 32752 46001 32804 46053
rect 48943 46139 48995 46145
rect 49154 46139 49206 46145
rect 49365 46139 49417 46145
rect 49576 46139 49628 46145
rect 49787 46139 49839 46145
rect 34755 46001 34807 46053
rect 34935 46050 34987 46053
rect 34935 46004 34962 46050
rect 34962 46004 34987 46050
rect 34935 46001 34987 46004
rect 50138 46050 50190 46053
rect 50138 46004 50160 46050
rect 50160 46004 50190 46050
rect 50138 46001 50190 46004
rect 50318 46001 50370 46053
rect 35332 45909 35384 45915
rect 35543 45909 35595 45915
rect 35754 45909 35806 45915
rect 35965 45909 36017 45915
rect 36176 45909 36228 45915
rect 37891 45909 37943 45917
rect 38071 45909 38123 45917
rect 52316 46001 52368 46053
rect 52527 46001 52579 46053
rect 52738 46001 52790 46053
rect 52948 46001 53000 46053
rect 53159 46001 53211 46053
rect 53371 46001 53423 46053
rect 53582 46001 53634 46053
rect 53792 46001 53844 46053
rect 54003 46001 54055 46053
rect 54214 46001 54266 46053
rect 54855 46001 54907 46053
rect 55066 46001 55118 46053
rect 55278 46050 55330 46053
rect 55278 46004 55279 46050
rect 55279 46004 55325 46050
rect 55325 46004 55330 46050
rect 55278 46001 55330 46004
rect 55489 46001 55541 46053
rect 56015 46001 56067 46053
rect 56226 46050 56278 46053
rect 56226 46004 56267 46050
rect 56267 46004 56278 46050
rect 56226 46001 56278 46004
rect 56437 46001 56489 46053
rect 56648 46001 56700 46053
rect 56859 46001 56911 46053
rect 57070 46001 57122 46053
rect 57281 46001 57333 46053
rect 48943 45909 48995 45915
rect 49154 45909 49206 45915
rect 49365 45909 49417 45915
rect 49576 45909 49628 45915
rect 49787 45909 49839 45915
rect 33057 45822 33109 45825
rect 33237 45822 33289 45825
rect 35332 45863 35384 45909
rect 35543 45863 35580 45909
rect 35580 45863 35595 45909
rect 35754 45863 35786 45909
rect 35786 45863 35806 45909
rect 35965 45863 35992 45909
rect 35992 45863 36017 45909
rect 36176 45863 36198 45909
rect 36198 45863 36228 45909
rect 37891 45865 37909 45909
rect 37909 45865 37943 45909
rect 38071 45865 38072 45909
rect 38072 45865 38123 45909
rect 33057 45776 33109 45822
rect 33237 45776 33289 45822
rect 33057 45773 33109 45776
rect 33237 45773 33289 45776
rect 33057 45374 33109 45377
rect 33237 45374 33289 45377
rect 33057 45328 33109 45374
rect 33237 45328 33289 45374
rect 33057 45325 33109 45328
rect 33237 45325 33289 45328
rect 29582 45101 29634 45153
rect 29793 45150 29845 45153
rect 29793 45104 29798 45150
rect 29798 45104 29844 45150
rect 29844 45104 29845 45150
rect 29793 45101 29845 45104
rect 30005 45101 30057 45153
rect 30216 45101 30268 45153
rect 34267 45598 34319 45615
rect 34447 45598 34499 45615
rect 34627 45598 34679 45615
rect 34267 45563 34302 45598
rect 34302 45563 34319 45598
rect 34447 45563 34451 45598
rect 34451 45563 34499 45598
rect 34627 45563 34658 45598
rect 34658 45563 34679 45598
rect 36678 45638 36697 45690
rect 36697 45638 36730 45690
rect 48943 45863 48984 45909
rect 48984 45863 48995 45909
rect 49154 45863 49190 45909
rect 49190 45863 49206 45909
rect 49365 45863 49396 45909
rect 49396 45863 49417 45909
rect 49576 45863 49602 45909
rect 49602 45863 49628 45909
rect 49787 45863 49839 45909
rect 39994 45740 40046 45792
rect 36961 45639 36971 45683
rect 36971 45639 37013 45683
rect 37172 45639 37206 45683
rect 37206 45639 37224 45683
rect 36961 45631 37013 45639
rect 37172 45631 37224 45639
rect 37384 45631 37436 45683
rect 37595 45631 37647 45683
rect 35332 45415 35384 45455
rect 35543 45415 35580 45455
rect 35580 45415 35595 45455
rect 35754 45415 35786 45455
rect 35786 45415 35806 45455
rect 35965 45415 35992 45455
rect 35992 45415 36017 45455
rect 36176 45415 36198 45455
rect 36198 45415 36228 45455
rect 37891 45415 37909 45443
rect 37909 45415 37943 45443
rect 38071 45415 38072 45443
rect 38072 45415 38123 45443
rect 35332 45403 35384 45415
rect 35543 45403 35595 45415
rect 35754 45403 35806 45415
rect 35965 45403 36017 45415
rect 36176 45403 36228 45415
rect 33819 45328 33833 45369
rect 33833 45328 33871 45369
rect 33999 45328 34039 45369
rect 34039 45328 34051 45369
rect 37891 45391 37943 45415
rect 38071 45391 38123 45415
rect 33819 45317 33871 45328
rect 33999 45317 34051 45328
rect 30854 45101 30906 45153
rect 31065 45101 31117 45153
rect 31276 45101 31328 45153
rect 31486 45150 31538 45153
rect 31697 45150 31749 45153
rect 31909 45150 31961 45153
rect 32120 45150 32172 45153
rect 32330 45150 32382 45153
rect 32541 45150 32593 45153
rect 32752 45150 32804 45153
rect 34284 45150 34336 45153
rect 34495 45150 34547 45153
rect 31486 45104 31538 45150
rect 31697 45104 31749 45150
rect 31909 45104 31961 45150
rect 32120 45104 32172 45150
rect 32330 45104 32382 45150
rect 32541 45104 32593 45150
rect 32752 45104 32804 45150
rect 34284 45104 34302 45150
rect 34302 45104 34336 45150
rect 34495 45104 34508 45150
rect 34508 45104 34547 45150
rect 31486 45101 31538 45104
rect 31697 45101 31749 45104
rect 31909 45101 31961 45104
rect 32120 45101 32172 45104
rect 32330 45101 32382 45104
rect 32541 45101 32593 45104
rect 32752 45101 32804 45104
rect 34284 45101 34336 45104
rect 34495 45101 34547 45104
rect 34707 45101 34759 45153
rect 34918 45101 34970 45153
rect 35220 45101 35272 45153
rect 35430 45101 35482 45153
rect 35641 45101 35693 45153
rect 35853 45101 35905 45153
rect 36064 45101 36116 45153
rect 36274 45101 36326 45153
rect 38330 45150 38382 45153
rect 38330 45104 38382 45150
rect 38330 45101 38382 45104
rect 38541 45101 38593 45153
rect 38752 45101 38804 45153
rect 39052 45150 39104 45153
rect 39232 45150 39284 45153
rect 39052 45104 39062 45150
rect 39062 45104 39104 45150
rect 39232 45104 39266 45150
rect 39266 45104 39284 45150
rect 39052 45101 39104 45104
rect 39232 45101 39284 45104
rect 33057 44926 33109 44929
rect 33237 44926 33289 44929
rect 33057 44880 33109 44926
rect 33237 44880 33289 44926
rect 33057 44877 33109 44880
rect 33237 44877 33289 44880
rect 33819 44926 33871 44937
rect 33999 44926 34051 44937
rect 33819 44885 33833 44926
rect 33833 44885 33871 44926
rect 33999 44885 34039 44926
rect 34039 44885 34051 44926
rect 35332 44839 35384 44851
rect 35543 44839 35595 44851
rect 35754 44839 35806 44851
rect 35965 44839 36017 44851
rect 36176 44839 36228 44851
rect 37891 44839 37943 44863
rect 38071 44839 38123 44863
rect 35332 44799 35384 44839
rect 35543 44799 35580 44839
rect 35580 44799 35595 44839
rect 35754 44799 35786 44839
rect 35786 44799 35806 44839
rect 35965 44799 35992 44839
rect 35992 44799 36017 44839
rect 36176 44799 36198 44839
rect 36198 44799 36228 44839
rect 37891 44811 37909 44839
rect 37909 44811 37943 44839
rect 38071 44811 38072 44839
rect 38072 44811 38123 44839
rect 34267 44656 34302 44691
rect 34302 44656 34319 44691
rect 34447 44656 34451 44691
rect 34451 44656 34499 44691
rect 34627 44656 34658 44691
rect 34658 44656 34679 44691
rect 34267 44639 34319 44656
rect 34447 44639 34499 44656
rect 34627 44639 34679 44656
rect 33057 44478 33109 44481
rect 33237 44478 33289 44481
rect 33057 44432 33109 44478
rect 33237 44432 33289 44478
rect 33057 44429 33109 44432
rect 33237 44429 33289 44432
rect 36678 44564 36697 44616
rect 36697 44564 36730 44616
rect 36961 44615 37013 44623
rect 37172 44615 37224 44623
rect 36961 44571 36971 44615
rect 36971 44571 37013 44615
rect 37172 44571 37206 44615
rect 37206 44571 37224 44615
rect 37384 44571 37436 44623
rect 37595 44571 37647 44623
rect 39994 45554 40046 45606
rect 39775 45374 39827 45391
rect 39775 45339 39786 45374
rect 39786 45339 39827 45374
rect 43068 45570 43120 45622
rect 41935 45339 41987 45391
rect 47486 45679 47538 45731
rect 48596 45725 48648 45777
rect 51835 45822 51887 45847
rect 52015 45822 52067 45847
rect 51835 45795 51887 45822
rect 52015 45795 52067 45822
rect 44939 45598 44991 45615
rect 45151 45598 45203 45615
rect 44939 45563 44971 45598
rect 44971 45563 44991 45598
rect 45151 45563 45197 45598
rect 45197 45563 45203 45598
rect 48596 45507 48648 45559
rect 50300 45563 50352 45615
rect 50511 45598 50563 45615
rect 50511 45563 50513 45598
rect 50513 45563 50563 45598
rect 50722 45563 50774 45615
rect 48943 45415 48984 45452
rect 48984 45415 48995 45452
rect 49154 45415 49190 45452
rect 49190 45415 49206 45452
rect 49365 45415 49396 45452
rect 49396 45415 49417 45452
rect 49576 45415 49602 45452
rect 49602 45415 49628 45452
rect 49787 45415 49839 45452
rect 48943 45400 48995 45415
rect 49154 45400 49206 45415
rect 49365 45400 49417 45415
rect 49576 45400 49628 45415
rect 49787 45400 49839 45415
rect 51073 45374 51125 45377
rect 51253 45374 51305 45377
rect 51073 45328 51086 45374
rect 51086 45328 51125 45374
rect 51253 45328 51292 45374
rect 51292 45328 51305 45374
rect 51073 45325 51125 45328
rect 51253 45325 51305 45328
rect 51835 45374 51887 45384
rect 52015 45374 52067 45384
rect 51835 45332 51887 45374
rect 52015 45332 52067 45374
rect 40253 45101 40305 45153
rect 40433 45101 40485 45153
rect 43790 45101 43842 45153
rect 44001 45101 44053 45153
rect 44213 45150 44265 45153
rect 44213 45104 44236 45150
rect 44236 45104 44265 45150
rect 44213 45101 44265 45104
rect 44424 45101 44476 45153
rect 44834 45150 44886 45153
rect 45045 45150 45097 45153
rect 45256 45150 45308 45153
rect 44834 45104 44858 45150
rect 44858 45104 44886 45150
rect 45045 45104 45084 45150
rect 45084 45104 45097 45150
rect 45256 45104 45264 45150
rect 45264 45104 45308 45150
rect 44834 45101 44886 45104
rect 45045 45101 45097 45104
rect 45256 45101 45308 45104
rect 48838 45101 48890 45153
rect 49048 45101 49100 45153
rect 49259 45101 49311 45153
rect 49471 45101 49523 45153
rect 49682 45101 49734 45153
rect 49892 45101 49944 45153
rect 50346 45101 50398 45153
rect 50557 45150 50609 45153
rect 50768 45150 50820 45153
rect 52316 45150 52368 45153
rect 52527 45150 52579 45153
rect 52738 45150 52790 45153
rect 52948 45150 53000 45153
rect 53159 45150 53211 45153
rect 53371 45150 53423 45153
rect 53582 45150 53634 45153
rect 50557 45104 50571 45150
rect 50571 45104 50609 45150
rect 50768 45104 50777 45150
rect 50777 45104 50820 45150
rect 52316 45104 52368 45150
rect 52527 45104 52579 45150
rect 52738 45104 52790 45150
rect 52948 45104 53000 45150
rect 53159 45104 53211 45150
rect 53371 45104 53423 45150
rect 53582 45104 53634 45150
rect 50557 45101 50609 45104
rect 50768 45101 50820 45104
rect 39775 44880 39786 44915
rect 39786 44880 39827 44915
rect 39775 44863 39827 44880
rect 39994 44648 40046 44700
rect 39994 44462 40046 44514
rect 52316 45101 52368 45104
rect 52527 45101 52579 45104
rect 52738 45101 52790 45104
rect 52948 45101 53000 45104
rect 53159 45101 53211 45104
rect 53371 45101 53423 45104
rect 53582 45101 53634 45104
rect 53792 45101 53844 45153
rect 54003 45101 54055 45153
rect 54214 45101 54266 45153
rect 54855 45101 54907 45153
rect 55066 45101 55118 45153
rect 55278 45150 55330 45153
rect 55278 45104 55279 45150
rect 55279 45104 55325 45150
rect 55325 45104 55330 45150
rect 55278 45101 55330 45104
rect 55489 45101 55541 45153
rect 41935 44863 41987 44915
rect 51073 44926 51125 44929
rect 51253 44926 51305 44929
rect 43068 44632 43120 44684
rect 51073 44880 51086 44926
rect 51086 44880 51125 44926
rect 51253 44880 51292 44926
rect 51292 44880 51305 44926
rect 48943 44839 48995 44854
rect 49154 44839 49206 44854
rect 49365 44839 49417 44854
rect 49576 44839 49628 44854
rect 49787 44839 49839 44854
rect 48943 44802 48984 44839
rect 48984 44802 48995 44839
rect 49154 44802 49190 44839
rect 49190 44802 49206 44839
rect 49365 44802 49396 44839
rect 49396 44802 49417 44839
rect 49576 44802 49602 44839
rect 49602 44802 49628 44839
rect 49787 44802 49839 44839
rect 51073 44877 51125 44880
rect 51253 44877 51305 44880
rect 44939 44656 44971 44691
rect 44971 44656 44991 44691
rect 45151 44656 45197 44691
rect 45197 44656 45203 44691
rect 48596 44695 48648 44747
rect 44939 44639 44991 44656
rect 45151 44639 45203 44656
rect 47864 44523 47916 44575
rect 50300 44639 50352 44691
rect 50511 44656 50513 44691
rect 50513 44656 50563 44691
rect 50511 44639 50563 44656
rect 50722 44639 50774 44691
rect 48596 44477 48648 44529
rect 51835 44880 51887 44922
rect 52015 44880 52067 44922
rect 51835 44870 51887 44880
rect 52015 44870 52067 44880
rect 35332 44345 35384 44391
rect 35543 44345 35580 44391
rect 35580 44345 35595 44391
rect 35754 44345 35786 44391
rect 35786 44345 35806 44391
rect 35965 44345 35992 44391
rect 35992 44345 36017 44391
rect 36176 44345 36198 44391
rect 36198 44345 36228 44391
rect 37891 44345 37909 44389
rect 37909 44345 37943 44389
rect 38071 44345 38072 44389
rect 38072 44345 38123 44389
rect 48943 44345 48984 44391
rect 48984 44345 48995 44391
rect 49154 44345 49190 44391
rect 49190 44345 49206 44391
rect 49365 44345 49396 44391
rect 49396 44345 49417 44391
rect 49576 44345 49602 44391
rect 49602 44345 49628 44391
rect 49787 44345 49839 44391
rect 51835 44432 51887 44459
rect 52015 44432 52067 44459
rect 51835 44407 51887 44432
rect 52015 44407 52067 44432
rect 35332 44339 35384 44345
rect 35543 44339 35595 44345
rect 35754 44339 35806 44345
rect 35965 44339 36017 44345
rect 36176 44339 36228 44345
rect 37891 44337 37943 44345
rect 38071 44337 38123 44345
rect 27790 44201 27842 44253
rect 28001 44201 28053 44253
rect 28212 44201 28264 44253
rect 28423 44201 28475 44253
rect 28634 44201 28686 44253
rect 28845 44250 28897 44253
rect 28845 44204 28856 44250
rect 28856 44204 28897 44250
rect 28845 44201 28897 44204
rect 29056 44201 29108 44253
rect 29582 44201 29634 44253
rect 29793 44250 29845 44253
rect 29793 44204 29798 44250
rect 29798 44204 29844 44250
rect 29844 44204 29845 44250
rect 29793 44201 29845 44204
rect 30005 44201 30057 44253
rect 30216 44201 30268 44253
rect 30854 44201 30906 44253
rect 31065 44201 31117 44253
rect 31276 44201 31328 44253
rect 31486 44201 31538 44253
rect 31697 44201 31749 44253
rect 31909 44201 31961 44253
rect 32120 44201 32172 44253
rect 32330 44201 32382 44253
rect 32541 44201 32593 44253
rect 32752 44201 32804 44253
rect 48943 44339 48995 44345
rect 49154 44339 49206 44345
rect 49365 44339 49417 44345
rect 49576 44339 49628 44345
rect 49787 44339 49839 44345
rect 34755 44201 34807 44253
rect 34935 44250 34987 44253
rect 34935 44204 34962 44250
rect 34962 44204 34987 44250
rect 34935 44201 34987 44204
rect 50138 44250 50190 44253
rect 50138 44204 50160 44250
rect 50160 44204 50190 44250
rect 50138 44201 50190 44204
rect 50318 44201 50370 44253
rect 35332 44109 35384 44115
rect 35543 44109 35595 44115
rect 35754 44109 35806 44115
rect 35965 44109 36017 44115
rect 36176 44109 36228 44115
rect 37891 44109 37943 44117
rect 38071 44109 38123 44117
rect 52316 44201 52368 44253
rect 52527 44201 52579 44253
rect 52738 44201 52790 44253
rect 52948 44201 53000 44253
rect 53159 44201 53211 44253
rect 53371 44201 53423 44253
rect 53582 44201 53634 44253
rect 53792 44201 53844 44253
rect 54003 44201 54055 44253
rect 54214 44201 54266 44253
rect 54855 44201 54907 44253
rect 55066 44201 55118 44253
rect 55278 44250 55330 44253
rect 55278 44204 55279 44250
rect 55279 44204 55325 44250
rect 55325 44204 55330 44250
rect 55278 44201 55330 44204
rect 55489 44201 55541 44253
rect 56015 44201 56067 44253
rect 56226 44250 56278 44253
rect 56226 44204 56267 44250
rect 56267 44204 56278 44250
rect 56226 44201 56278 44204
rect 56437 44201 56489 44253
rect 56648 44201 56700 44253
rect 56859 44201 56911 44253
rect 57070 44201 57122 44253
rect 57281 44201 57333 44253
rect 48943 44109 48995 44115
rect 49154 44109 49206 44115
rect 49365 44109 49417 44115
rect 49576 44109 49628 44115
rect 49787 44109 49839 44115
rect 33057 44022 33109 44025
rect 33237 44022 33289 44025
rect 35332 44063 35384 44109
rect 35543 44063 35580 44109
rect 35580 44063 35595 44109
rect 35754 44063 35786 44109
rect 35786 44063 35806 44109
rect 35965 44063 35992 44109
rect 35992 44063 36017 44109
rect 36176 44063 36198 44109
rect 36198 44063 36228 44109
rect 37891 44065 37909 44109
rect 37909 44065 37943 44109
rect 38071 44065 38072 44109
rect 38072 44065 38123 44109
rect 33057 43976 33109 44022
rect 33237 43976 33289 44022
rect 33057 43973 33109 43976
rect 33237 43973 33289 43976
rect 33057 43574 33109 43577
rect 33237 43574 33289 43577
rect 33057 43528 33109 43574
rect 33237 43528 33289 43574
rect 33057 43525 33109 43528
rect 33237 43525 33289 43528
rect 29582 43301 29634 43353
rect 29793 43350 29845 43353
rect 29793 43304 29798 43350
rect 29798 43304 29844 43350
rect 29844 43304 29845 43350
rect 29793 43301 29845 43304
rect 30005 43301 30057 43353
rect 30216 43301 30268 43353
rect 34267 43798 34319 43815
rect 34447 43798 34499 43815
rect 34627 43798 34679 43815
rect 34267 43763 34302 43798
rect 34302 43763 34319 43798
rect 34447 43763 34451 43798
rect 34451 43763 34499 43798
rect 34627 43763 34658 43798
rect 34658 43763 34679 43798
rect 36678 43838 36697 43890
rect 36697 43838 36730 43890
rect 48943 44063 48984 44109
rect 48984 44063 48995 44109
rect 49154 44063 49190 44109
rect 49190 44063 49206 44109
rect 49365 44063 49396 44109
rect 49396 44063 49417 44109
rect 49576 44063 49602 44109
rect 49602 44063 49628 44109
rect 49787 44063 49839 44109
rect 39994 43940 40046 43992
rect 36961 43839 36971 43883
rect 36971 43839 37013 43883
rect 37172 43839 37206 43883
rect 37206 43839 37224 43883
rect 36961 43831 37013 43839
rect 37172 43831 37224 43839
rect 37384 43831 37436 43883
rect 37595 43831 37647 43883
rect 35332 43615 35384 43655
rect 35543 43615 35580 43655
rect 35580 43615 35595 43655
rect 35754 43615 35786 43655
rect 35786 43615 35806 43655
rect 35965 43615 35992 43655
rect 35992 43615 36017 43655
rect 36176 43615 36198 43655
rect 36198 43615 36228 43655
rect 37891 43615 37909 43643
rect 37909 43615 37943 43643
rect 38071 43615 38072 43643
rect 38072 43615 38123 43643
rect 35332 43603 35384 43615
rect 35543 43603 35595 43615
rect 35754 43603 35806 43615
rect 35965 43603 36017 43615
rect 36176 43603 36228 43615
rect 33819 43528 33833 43569
rect 33833 43528 33871 43569
rect 33999 43528 34039 43569
rect 34039 43528 34051 43569
rect 37891 43591 37943 43615
rect 38071 43591 38123 43615
rect 33819 43517 33871 43528
rect 33999 43517 34051 43528
rect 30854 43301 30906 43353
rect 31065 43301 31117 43353
rect 31276 43301 31328 43353
rect 31486 43350 31538 43353
rect 31697 43350 31749 43353
rect 31909 43350 31961 43353
rect 32120 43350 32172 43353
rect 32330 43350 32382 43353
rect 32541 43350 32593 43353
rect 32752 43350 32804 43353
rect 34284 43350 34336 43353
rect 34495 43350 34547 43353
rect 31486 43304 31538 43350
rect 31697 43304 31749 43350
rect 31909 43304 31961 43350
rect 32120 43304 32172 43350
rect 32330 43304 32382 43350
rect 32541 43304 32593 43350
rect 32752 43304 32804 43350
rect 34284 43304 34302 43350
rect 34302 43304 34336 43350
rect 34495 43304 34508 43350
rect 34508 43304 34547 43350
rect 31486 43301 31538 43304
rect 31697 43301 31749 43304
rect 31909 43301 31961 43304
rect 32120 43301 32172 43304
rect 32330 43301 32382 43304
rect 32541 43301 32593 43304
rect 32752 43301 32804 43304
rect 34284 43301 34336 43304
rect 34495 43301 34547 43304
rect 34707 43301 34759 43353
rect 34918 43301 34970 43353
rect 35220 43301 35272 43353
rect 35430 43301 35482 43353
rect 35641 43301 35693 43353
rect 35853 43301 35905 43353
rect 36064 43301 36116 43353
rect 36274 43301 36326 43353
rect 38330 43350 38382 43353
rect 38330 43304 38382 43350
rect 38330 43301 38382 43304
rect 38541 43301 38593 43353
rect 38752 43301 38804 43353
rect 39052 43350 39104 43353
rect 39232 43350 39284 43353
rect 39052 43304 39062 43350
rect 39062 43304 39104 43350
rect 39232 43304 39266 43350
rect 39266 43304 39284 43350
rect 39052 43301 39104 43304
rect 39232 43301 39284 43304
rect 33057 43126 33109 43129
rect 33237 43126 33289 43129
rect 33057 43080 33109 43126
rect 33237 43080 33289 43126
rect 33057 43077 33109 43080
rect 33237 43077 33289 43080
rect 33819 43126 33871 43137
rect 33999 43126 34051 43137
rect 33819 43085 33833 43126
rect 33833 43085 33871 43126
rect 33999 43085 34039 43126
rect 34039 43085 34051 43126
rect 35332 43039 35384 43051
rect 35543 43039 35595 43051
rect 35754 43039 35806 43051
rect 35965 43039 36017 43051
rect 36176 43039 36228 43051
rect 37891 43039 37943 43063
rect 38071 43039 38123 43063
rect 35332 42999 35384 43039
rect 35543 42999 35580 43039
rect 35580 42999 35595 43039
rect 35754 42999 35786 43039
rect 35786 42999 35806 43039
rect 35965 42999 35992 43039
rect 35992 42999 36017 43039
rect 36176 42999 36198 43039
rect 36198 42999 36228 43039
rect 37891 43011 37909 43039
rect 37909 43011 37943 43039
rect 38071 43011 38072 43039
rect 38072 43011 38123 43039
rect 34267 42856 34302 42891
rect 34302 42856 34319 42891
rect 34447 42856 34451 42891
rect 34451 42856 34499 42891
rect 34627 42856 34658 42891
rect 34658 42856 34679 42891
rect 34267 42839 34319 42856
rect 34447 42839 34499 42856
rect 34627 42839 34679 42856
rect 33057 42678 33109 42681
rect 33237 42678 33289 42681
rect 33057 42632 33109 42678
rect 33237 42632 33289 42678
rect 33057 42629 33109 42632
rect 33237 42629 33289 42632
rect 36678 42764 36697 42816
rect 36697 42764 36730 42816
rect 36961 42815 37013 42823
rect 37172 42815 37224 42823
rect 36961 42771 36971 42815
rect 36971 42771 37013 42815
rect 37172 42771 37206 42815
rect 37206 42771 37224 42815
rect 37384 42771 37436 42823
rect 37595 42771 37647 42823
rect 39994 43754 40046 43806
rect 39775 43574 39827 43591
rect 39775 43539 39786 43574
rect 39786 43539 39827 43574
rect 43068 43770 43120 43822
rect 41935 43539 41987 43591
rect 48241 43879 48293 43931
rect 48596 43925 48648 43977
rect 51835 44022 51887 44047
rect 52015 44022 52067 44047
rect 51835 43995 51887 44022
rect 52015 43995 52067 44022
rect 44939 43798 44991 43815
rect 45151 43798 45203 43815
rect 44939 43763 44971 43798
rect 44971 43763 44991 43798
rect 45151 43763 45197 43798
rect 45197 43763 45203 43798
rect 48596 43707 48648 43759
rect 50300 43763 50352 43815
rect 50511 43798 50563 43815
rect 50511 43763 50513 43798
rect 50513 43763 50563 43798
rect 50722 43763 50774 43815
rect 48943 43615 48984 43652
rect 48984 43615 48995 43652
rect 49154 43615 49190 43652
rect 49190 43615 49206 43652
rect 49365 43615 49396 43652
rect 49396 43615 49417 43652
rect 49576 43615 49602 43652
rect 49602 43615 49628 43652
rect 49787 43615 49839 43652
rect 48943 43600 48995 43615
rect 49154 43600 49206 43615
rect 49365 43600 49417 43615
rect 49576 43600 49628 43615
rect 49787 43600 49839 43615
rect 51073 43574 51125 43577
rect 51253 43574 51305 43577
rect 51073 43528 51086 43574
rect 51086 43528 51125 43574
rect 51253 43528 51292 43574
rect 51292 43528 51305 43574
rect 51073 43525 51125 43528
rect 51253 43525 51305 43528
rect 51835 43574 51887 43584
rect 52015 43574 52067 43584
rect 51835 43532 51887 43574
rect 52015 43532 52067 43574
rect 40253 43301 40305 43353
rect 40433 43301 40485 43353
rect 43790 43301 43842 43353
rect 44001 43301 44053 43353
rect 44213 43350 44265 43353
rect 44213 43304 44236 43350
rect 44236 43304 44265 43350
rect 44213 43301 44265 43304
rect 44424 43301 44476 43353
rect 44834 43350 44886 43353
rect 45045 43350 45097 43353
rect 45256 43350 45308 43353
rect 44834 43304 44858 43350
rect 44858 43304 44886 43350
rect 45045 43304 45084 43350
rect 45084 43304 45097 43350
rect 45256 43304 45264 43350
rect 45264 43304 45308 43350
rect 44834 43301 44886 43304
rect 45045 43301 45097 43304
rect 45256 43301 45308 43304
rect 48838 43301 48890 43353
rect 49048 43301 49100 43353
rect 49259 43301 49311 43353
rect 49471 43301 49523 43353
rect 49682 43301 49734 43353
rect 49892 43301 49944 43353
rect 50346 43301 50398 43353
rect 50557 43350 50609 43353
rect 50768 43350 50820 43353
rect 52316 43350 52368 43353
rect 52527 43350 52579 43353
rect 52738 43350 52790 43353
rect 52948 43350 53000 43353
rect 53159 43350 53211 43353
rect 53371 43350 53423 43353
rect 53582 43350 53634 43353
rect 50557 43304 50571 43350
rect 50571 43304 50609 43350
rect 50768 43304 50777 43350
rect 50777 43304 50820 43350
rect 52316 43304 52368 43350
rect 52527 43304 52579 43350
rect 52738 43304 52790 43350
rect 52948 43304 53000 43350
rect 53159 43304 53211 43350
rect 53371 43304 53423 43350
rect 53582 43304 53634 43350
rect 50557 43301 50609 43304
rect 50768 43301 50820 43304
rect 39775 43080 39786 43115
rect 39786 43080 39827 43115
rect 39775 43063 39827 43080
rect 39994 42848 40046 42900
rect 39994 42662 40046 42714
rect 52316 43301 52368 43304
rect 52527 43301 52579 43304
rect 52738 43301 52790 43304
rect 52948 43301 53000 43304
rect 53159 43301 53211 43304
rect 53371 43301 53423 43304
rect 53582 43301 53634 43304
rect 53792 43301 53844 43353
rect 54003 43301 54055 43353
rect 54214 43301 54266 43353
rect 54855 43301 54907 43353
rect 55066 43301 55118 43353
rect 55278 43350 55330 43353
rect 55278 43304 55279 43350
rect 55279 43304 55325 43350
rect 55325 43304 55330 43350
rect 55278 43301 55330 43304
rect 55489 43301 55541 43353
rect 41935 43063 41987 43115
rect 51073 43126 51125 43129
rect 51253 43126 51305 43129
rect 43445 42832 43497 42884
rect 51073 43080 51086 43126
rect 51086 43080 51125 43126
rect 51253 43080 51292 43126
rect 51292 43080 51305 43126
rect 48943 43039 48995 43054
rect 49154 43039 49206 43054
rect 49365 43039 49417 43054
rect 49576 43039 49628 43054
rect 49787 43039 49839 43054
rect 48943 43002 48984 43039
rect 48984 43002 48995 43039
rect 49154 43002 49190 43039
rect 49190 43002 49206 43039
rect 49365 43002 49396 43039
rect 49396 43002 49417 43039
rect 49576 43002 49602 43039
rect 49602 43002 49628 43039
rect 49787 43002 49839 43039
rect 51073 43077 51125 43080
rect 51253 43077 51305 43080
rect 44939 42856 44971 42891
rect 44971 42856 44991 42891
rect 45151 42856 45197 42891
rect 45197 42856 45203 42891
rect 48596 42895 48648 42947
rect 44939 42839 44991 42856
rect 45151 42839 45203 42856
rect 45597 42737 45604 42775
rect 45604 42737 45649 42775
rect 45597 42723 45649 42737
rect 50300 42839 50352 42891
rect 50511 42856 50513 42891
rect 50513 42856 50563 42891
rect 50511 42839 50563 42856
rect 50722 42839 50774 42891
rect 48596 42677 48648 42729
rect 51835 43080 51887 43122
rect 52015 43080 52067 43122
rect 51835 43070 51887 43080
rect 52015 43070 52067 43080
rect 35332 42545 35384 42591
rect 35543 42545 35580 42591
rect 35580 42545 35595 42591
rect 35754 42545 35786 42591
rect 35786 42545 35806 42591
rect 35965 42545 35992 42591
rect 35992 42545 36017 42591
rect 36176 42545 36198 42591
rect 36198 42545 36228 42591
rect 37891 42545 37909 42589
rect 37909 42545 37943 42589
rect 38071 42545 38072 42589
rect 38072 42545 38123 42589
rect 48943 42545 48984 42591
rect 48984 42545 48995 42591
rect 49154 42545 49190 42591
rect 49190 42545 49206 42591
rect 49365 42545 49396 42591
rect 49396 42545 49417 42591
rect 49576 42545 49602 42591
rect 49602 42545 49628 42591
rect 49787 42545 49839 42591
rect 51835 42632 51887 42659
rect 52015 42632 52067 42659
rect 51835 42607 51887 42632
rect 52015 42607 52067 42632
rect 35332 42539 35384 42545
rect 35543 42539 35595 42545
rect 35754 42539 35806 42545
rect 35965 42539 36017 42545
rect 36176 42539 36228 42545
rect 37891 42537 37943 42545
rect 38071 42537 38123 42545
rect 27790 42401 27842 42453
rect 28001 42401 28053 42453
rect 28212 42401 28264 42453
rect 28423 42401 28475 42453
rect 28634 42401 28686 42453
rect 28845 42450 28897 42453
rect 28845 42404 28856 42450
rect 28856 42404 28897 42450
rect 28845 42401 28897 42404
rect 29056 42401 29108 42453
rect 29582 42401 29634 42453
rect 29793 42450 29845 42453
rect 29793 42404 29798 42450
rect 29798 42404 29844 42450
rect 29844 42404 29845 42450
rect 29793 42401 29845 42404
rect 30005 42401 30057 42453
rect 30216 42401 30268 42453
rect 30854 42401 30906 42453
rect 31065 42401 31117 42453
rect 31276 42401 31328 42453
rect 31486 42401 31538 42453
rect 31697 42401 31749 42453
rect 31909 42401 31961 42453
rect 32120 42401 32172 42453
rect 32330 42401 32382 42453
rect 32541 42401 32593 42453
rect 32752 42401 32804 42453
rect 48943 42539 48995 42545
rect 49154 42539 49206 42545
rect 49365 42539 49417 42545
rect 49576 42539 49628 42545
rect 49787 42539 49839 42545
rect 34755 42401 34807 42453
rect 34935 42450 34987 42453
rect 34935 42404 34962 42450
rect 34962 42404 34987 42450
rect 34935 42401 34987 42404
rect 50138 42450 50190 42453
rect 50138 42404 50160 42450
rect 50160 42404 50190 42450
rect 50138 42401 50190 42404
rect 50318 42401 50370 42453
rect 35332 42309 35384 42315
rect 35543 42309 35595 42315
rect 35754 42309 35806 42315
rect 35965 42309 36017 42315
rect 36176 42309 36228 42315
rect 37891 42309 37943 42317
rect 38071 42309 38123 42317
rect 52316 42401 52368 42453
rect 52527 42401 52579 42453
rect 52738 42401 52790 42453
rect 52948 42401 53000 42453
rect 53159 42401 53211 42453
rect 53371 42401 53423 42453
rect 53582 42401 53634 42453
rect 53792 42401 53844 42453
rect 54003 42401 54055 42453
rect 54214 42401 54266 42453
rect 54855 42401 54907 42453
rect 55066 42401 55118 42453
rect 55278 42450 55330 42453
rect 55278 42404 55279 42450
rect 55279 42404 55325 42450
rect 55325 42404 55330 42450
rect 55278 42401 55330 42404
rect 55489 42401 55541 42453
rect 56015 42401 56067 42453
rect 56226 42450 56278 42453
rect 56226 42404 56267 42450
rect 56267 42404 56278 42450
rect 56226 42401 56278 42404
rect 56437 42401 56489 42453
rect 56648 42401 56700 42453
rect 56859 42401 56911 42453
rect 57070 42401 57122 42453
rect 57281 42401 57333 42453
rect 48943 42309 48995 42315
rect 49154 42309 49206 42315
rect 49365 42309 49417 42315
rect 49576 42309 49628 42315
rect 49787 42309 49839 42315
rect 33057 42222 33109 42225
rect 33237 42222 33289 42225
rect 35332 42263 35384 42309
rect 35543 42263 35580 42309
rect 35580 42263 35595 42309
rect 35754 42263 35786 42309
rect 35786 42263 35806 42309
rect 35965 42263 35992 42309
rect 35992 42263 36017 42309
rect 36176 42263 36198 42309
rect 36198 42263 36228 42309
rect 37891 42265 37909 42309
rect 37909 42265 37943 42309
rect 38071 42265 38072 42309
rect 38072 42265 38123 42309
rect 33057 42176 33109 42222
rect 33237 42176 33289 42222
rect 33057 42173 33109 42176
rect 33237 42173 33289 42176
rect 33057 41774 33109 41777
rect 33237 41774 33289 41777
rect 33057 41728 33109 41774
rect 33237 41728 33289 41774
rect 33057 41725 33109 41728
rect 33237 41725 33289 41728
rect 29582 41501 29634 41553
rect 29793 41550 29845 41553
rect 29793 41504 29798 41550
rect 29798 41504 29844 41550
rect 29844 41504 29845 41550
rect 29793 41501 29845 41504
rect 30005 41501 30057 41553
rect 30216 41501 30268 41553
rect 34267 41998 34319 42015
rect 34447 41998 34499 42015
rect 34627 41998 34679 42015
rect 34267 41963 34302 41998
rect 34302 41963 34319 41998
rect 34447 41963 34451 41998
rect 34451 41963 34499 41998
rect 34627 41963 34658 41998
rect 34658 41963 34679 41998
rect 36678 42038 36697 42090
rect 36697 42038 36730 42090
rect 48943 42263 48984 42309
rect 48984 42263 48995 42309
rect 49154 42263 49190 42309
rect 49190 42263 49206 42309
rect 49365 42263 49396 42309
rect 49396 42263 49417 42309
rect 49576 42263 49602 42309
rect 49602 42263 49628 42309
rect 49787 42263 49839 42309
rect 39994 42140 40046 42192
rect 36961 42039 36971 42083
rect 36971 42039 37013 42083
rect 37172 42039 37206 42083
rect 37206 42039 37224 42083
rect 36961 42031 37013 42039
rect 37172 42031 37224 42039
rect 37384 42031 37436 42083
rect 37595 42031 37647 42083
rect 35332 41815 35384 41855
rect 35543 41815 35580 41855
rect 35580 41815 35595 41855
rect 35754 41815 35786 41855
rect 35786 41815 35806 41855
rect 35965 41815 35992 41855
rect 35992 41815 36017 41855
rect 36176 41815 36198 41855
rect 36198 41815 36228 41855
rect 37891 41815 37909 41843
rect 37909 41815 37943 41843
rect 38071 41815 38072 41843
rect 38072 41815 38123 41843
rect 35332 41803 35384 41815
rect 35543 41803 35595 41815
rect 35754 41803 35806 41815
rect 35965 41803 36017 41815
rect 36176 41803 36228 41815
rect 33819 41728 33833 41769
rect 33833 41728 33871 41769
rect 33999 41728 34039 41769
rect 34039 41728 34051 41769
rect 37891 41791 37943 41815
rect 38071 41791 38123 41815
rect 33819 41717 33871 41728
rect 33999 41717 34051 41728
rect 30854 41501 30906 41553
rect 31065 41501 31117 41553
rect 31276 41501 31328 41553
rect 31486 41550 31538 41553
rect 31697 41550 31749 41553
rect 31909 41550 31961 41553
rect 32120 41550 32172 41553
rect 32330 41550 32382 41553
rect 32541 41550 32593 41553
rect 32752 41550 32804 41553
rect 34284 41550 34336 41553
rect 34495 41550 34547 41553
rect 31486 41504 31538 41550
rect 31697 41504 31749 41550
rect 31909 41504 31961 41550
rect 32120 41504 32172 41550
rect 32330 41504 32382 41550
rect 32541 41504 32593 41550
rect 32752 41504 32804 41550
rect 34284 41504 34302 41550
rect 34302 41504 34336 41550
rect 34495 41504 34508 41550
rect 34508 41504 34547 41550
rect 31486 41501 31538 41504
rect 31697 41501 31749 41504
rect 31909 41501 31961 41504
rect 32120 41501 32172 41504
rect 32330 41501 32382 41504
rect 32541 41501 32593 41504
rect 32752 41501 32804 41504
rect 34284 41501 34336 41504
rect 34495 41501 34547 41504
rect 34707 41501 34759 41553
rect 34918 41501 34970 41553
rect 35220 41501 35272 41553
rect 35430 41501 35482 41553
rect 35641 41501 35693 41553
rect 35853 41501 35905 41553
rect 36064 41501 36116 41553
rect 36274 41501 36326 41553
rect 38330 41550 38382 41553
rect 38330 41504 38382 41550
rect 38330 41501 38382 41504
rect 38541 41501 38593 41553
rect 38752 41501 38804 41553
rect 39052 41550 39104 41553
rect 39232 41550 39284 41553
rect 39052 41504 39062 41550
rect 39062 41504 39104 41550
rect 39232 41504 39266 41550
rect 39266 41504 39284 41550
rect 39052 41501 39104 41504
rect 39232 41501 39284 41504
rect 33057 41326 33109 41329
rect 33237 41326 33289 41329
rect 33057 41280 33109 41326
rect 33237 41280 33289 41326
rect 33057 41277 33109 41280
rect 33237 41277 33289 41280
rect 33819 41326 33871 41337
rect 33999 41326 34051 41337
rect 33819 41285 33833 41326
rect 33833 41285 33871 41326
rect 33999 41285 34039 41326
rect 34039 41285 34051 41326
rect 35332 41239 35384 41251
rect 35543 41239 35595 41251
rect 35754 41239 35806 41251
rect 35965 41239 36017 41251
rect 36176 41239 36228 41251
rect 37891 41239 37943 41263
rect 38071 41239 38123 41263
rect 35332 41199 35384 41239
rect 35543 41199 35580 41239
rect 35580 41199 35595 41239
rect 35754 41199 35786 41239
rect 35786 41199 35806 41239
rect 35965 41199 35992 41239
rect 35992 41199 36017 41239
rect 36176 41199 36198 41239
rect 36198 41199 36228 41239
rect 37891 41211 37909 41239
rect 37909 41211 37943 41239
rect 38071 41211 38072 41239
rect 38072 41211 38123 41239
rect 34267 41056 34302 41091
rect 34302 41056 34319 41091
rect 34447 41056 34451 41091
rect 34451 41056 34499 41091
rect 34627 41056 34658 41091
rect 34658 41056 34679 41091
rect 34267 41039 34319 41056
rect 34447 41039 34499 41056
rect 34627 41039 34679 41056
rect 33057 40878 33109 40881
rect 33237 40878 33289 40881
rect 33057 40832 33109 40878
rect 33237 40832 33289 40878
rect 33057 40829 33109 40832
rect 33237 40829 33289 40832
rect 36678 40964 36697 41016
rect 36697 40964 36730 41016
rect 36961 41015 37013 41023
rect 37172 41015 37224 41023
rect 36961 40971 36971 41015
rect 36971 40971 37013 41015
rect 37172 40971 37206 41015
rect 37206 40971 37224 41015
rect 37384 40971 37436 41023
rect 37595 40971 37647 41023
rect 39994 41954 40046 42006
rect 39775 41774 39827 41791
rect 39775 41739 39786 41774
rect 39786 41739 39827 41774
rect 43445 41970 43497 42022
rect 41935 41739 41987 41791
rect 45975 42079 46027 42131
rect 48596 42125 48648 42177
rect 51835 42222 51887 42247
rect 52015 42222 52067 42247
rect 51835 42195 51887 42222
rect 52015 42195 52067 42222
rect 44939 41998 44991 42015
rect 45151 41998 45203 42015
rect 44939 41963 44971 41998
rect 44971 41963 44991 41998
rect 45151 41963 45197 41998
rect 45197 41963 45203 41998
rect 48596 41907 48648 41959
rect 50300 41963 50352 42015
rect 50511 41998 50563 42015
rect 50511 41963 50513 41998
rect 50513 41963 50563 41998
rect 50722 41963 50774 42015
rect 48943 41815 48984 41852
rect 48984 41815 48995 41852
rect 49154 41815 49190 41852
rect 49190 41815 49206 41852
rect 49365 41815 49396 41852
rect 49396 41815 49417 41852
rect 49576 41815 49602 41852
rect 49602 41815 49628 41852
rect 49787 41815 49839 41852
rect 48943 41800 48995 41815
rect 49154 41800 49206 41815
rect 49365 41800 49417 41815
rect 49576 41800 49628 41815
rect 49787 41800 49839 41815
rect 51073 41774 51125 41777
rect 51253 41774 51305 41777
rect 51073 41728 51086 41774
rect 51086 41728 51125 41774
rect 51253 41728 51292 41774
rect 51292 41728 51305 41774
rect 51073 41725 51125 41728
rect 51253 41725 51305 41728
rect 51835 41774 51887 41784
rect 52015 41774 52067 41784
rect 51835 41732 51887 41774
rect 52015 41732 52067 41774
rect 40253 41501 40305 41553
rect 40433 41501 40485 41553
rect 43790 41501 43842 41553
rect 44001 41501 44053 41553
rect 44213 41550 44265 41553
rect 44213 41504 44236 41550
rect 44236 41504 44265 41550
rect 44213 41501 44265 41504
rect 44424 41501 44476 41553
rect 44834 41550 44886 41553
rect 45045 41550 45097 41553
rect 45256 41550 45308 41553
rect 44834 41504 44858 41550
rect 44858 41504 44886 41550
rect 45045 41504 45084 41550
rect 45084 41504 45097 41550
rect 45256 41504 45264 41550
rect 45264 41504 45308 41550
rect 44834 41501 44886 41504
rect 45045 41501 45097 41504
rect 45256 41501 45308 41504
rect 48838 41501 48890 41553
rect 49048 41501 49100 41553
rect 49259 41501 49311 41553
rect 49471 41501 49523 41553
rect 49682 41501 49734 41553
rect 49892 41501 49944 41553
rect 50346 41501 50398 41553
rect 50557 41550 50609 41553
rect 50768 41550 50820 41553
rect 52316 41550 52368 41553
rect 52527 41550 52579 41553
rect 52738 41550 52790 41553
rect 52948 41550 53000 41553
rect 53159 41550 53211 41553
rect 53371 41550 53423 41553
rect 53582 41550 53634 41553
rect 50557 41504 50571 41550
rect 50571 41504 50609 41550
rect 50768 41504 50777 41550
rect 50777 41504 50820 41550
rect 52316 41504 52368 41550
rect 52527 41504 52579 41550
rect 52738 41504 52790 41550
rect 52948 41504 53000 41550
rect 53159 41504 53211 41550
rect 53371 41504 53423 41550
rect 53582 41504 53634 41550
rect 50557 41501 50609 41504
rect 50768 41501 50820 41504
rect 39775 41280 39786 41315
rect 39786 41280 39827 41315
rect 39775 41263 39827 41280
rect 39994 41048 40046 41100
rect 39994 40862 40046 40914
rect 52316 41501 52368 41504
rect 52527 41501 52579 41504
rect 52738 41501 52790 41504
rect 52948 41501 53000 41504
rect 53159 41501 53211 41504
rect 53371 41501 53423 41504
rect 53582 41501 53634 41504
rect 53792 41501 53844 41553
rect 54003 41501 54055 41553
rect 54214 41501 54266 41553
rect 54855 41501 54907 41553
rect 55066 41501 55118 41553
rect 55278 41550 55330 41553
rect 55278 41504 55279 41550
rect 55279 41504 55325 41550
rect 55325 41504 55330 41550
rect 55278 41501 55330 41504
rect 55489 41501 55541 41553
rect 41935 41263 41987 41315
rect 51073 41326 51125 41329
rect 51253 41326 51305 41329
rect 43445 41032 43497 41084
rect 51073 41280 51086 41326
rect 51086 41280 51125 41326
rect 51253 41280 51292 41326
rect 51292 41280 51305 41326
rect 48943 41239 48995 41254
rect 49154 41239 49206 41254
rect 49365 41239 49417 41254
rect 49576 41239 49628 41254
rect 49787 41239 49839 41254
rect 48943 41202 48984 41239
rect 48984 41202 48995 41239
rect 49154 41202 49190 41239
rect 49190 41202 49206 41239
rect 49365 41202 49396 41239
rect 49396 41202 49417 41239
rect 49576 41202 49602 41239
rect 49602 41202 49628 41239
rect 49787 41202 49839 41239
rect 51073 41277 51125 41280
rect 51253 41277 51305 41280
rect 44939 41056 44971 41091
rect 44971 41056 44991 41091
rect 45151 41056 45197 41091
rect 45197 41056 45203 41091
rect 48596 41095 48648 41147
rect 44939 41039 44991 41056
rect 45151 41039 45203 41056
rect 46353 40923 46405 40975
rect 50300 41039 50352 41091
rect 50511 41056 50513 41091
rect 50513 41056 50563 41091
rect 50511 41039 50563 41056
rect 50722 41039 50774 41091
rect 48596 40877 48648 40929
rect 51835 41280 51887 41322
rect 52015 41280 52067 41322
rect 51835 41270 51887 41280
rect 52015 41270 52067 41280
rect 35332 40745 35384 40791
rect 35543 40745 35580 40791
rect 35580 40745 35595 40791
rect 35754 40745 35786 40791
rect 35786 40745 35806 40791
rect 35965 40745 35992 40791
rect 35992 40745 36017 40791
rect 36176 40745 36198 40791
rect 36198 40745 36228 40791
rect 37891 40745 37909 40789
rect 37909 40745 37943 40789
rect 38071 40745 38072 40789
rect 38072 40745 38123 40789
rect 48943 40745 48984 40791
rect 48984 40745 48995 40791
rect 49154 40745 49190 40791
rect 49190 40745 49206 40791
rect 49365 40745 49396 40791
rect 49396 40745 49417 40791
rect 49576 40745 49602 40791
rect 49602 40745 49628 40791
rect 49787 40745 49839 40791
rect 51835 40832 51887 40859
rect 52015 40832 52067 40859
rect 51835 40807 51887 40832
rect 52015 40807 52067 40832
rect 35332 40739 35384 40745
rect 35543 40739 35595 40745
rect 35754 40739 35806 40745
rect 35965 40739 36017 40745
rect 36176 40739 36228 40745
rect 37891 40737 37943 40745
rect 38071 40737 38123 40745
rect 27790 40601 27842 40653
rect 28001 40601 28053 40653
rect 28212 40601 28264 40653
rect 28423 40601 28475 40653
rect 28634 40601 28686 40653
rect 28845 40650 28897 40653
rect 28845 40604 28856 40650
rect 28856 40604 28897 40650
rect 28845 40601 28897 40604
rect 29056 40601 29108 40653
rect 29582 40601 29634 40653
rect 29793 40650 29845 40653
rect 29793 40604 29798 40650
rect 29798 40604 29844 40650
rect 29844 40604 29845 40650
rect 29793 40601 29845 40604
rect 30005 40601 30057 40653
rect 30216 40601 30268 40653
rect 30854 40601 30906 40653
rect 31065 40601 31117 40653
rect 31276 40601 31328 40653
rect 31486 40601 31538 40653
rect 31697 40601 31749 40653
rect 31909 40601 31961 40653
rect 32120 40601 32172 40653
rect 32330 40601 32382 40653
rect 32541 40601 32593 40653
rect 32752 40601 32804 40653
rect 48943 40739 48995 40745
rect 49154 40739 49206 40745
rect 49365 40739 49417 40745
rect 49576 40739 49628 40745
rect 49787 40739 49839 40745
rect 34755 40601 34807 40653
rect 34935 40650 34987 40653
rect 34935 40604 34962 40650
rect 34962 40604 34987 40650
rect 34935 40601 34987 40604
rect 50138 40650 50190 40653
rect 50138 40604 50160 40650
rect 50160 40604 50190 40650
rect 50138 40601 50190 40604
rect 50318 40601 50370 40653
rect 35332 40509 35384 40515
rect 35543 40509 35595 40515
rect 35754 40509 35806 40515
rect 35965 40509 36017 40515
rect 36176 40509 36228 40515
rect 37891 40509 37943 40517
rect 38071 40509 38123 40517
rect 52316 40601 52368 40653
rect 52527 40601 52579 40653
rect 52738 40601 52790 40653
rect 52948 40601 53000 40653
rect 53159 40601 53211 40653
rect 53371 40601 53423 40653
rect 53582 40601 53634 40653
rect 53792 40601 53844 40653
rect 54003 40601 54055 40653
rect 54214 40601 54266 40653
rect 54855 40601 54907 40653
rect 55066 40601 55118 40653
rect 55278 40650 55330 40653
rect 55278 40604 55279 40650
rect 55279 40604 55325 40650
rect 55325 40604 55330 40650
rect 55278 40601 55330 40604
rect 55489 40601 55541 40653
rect 56015 40601 56067 40653
rect 56226 40650 56278 40653
rect 56226 40604 56267 40650
rect 56267 40604 56278 40650
rect 56226 40601 56278 40604
rect 56437 40601 56489 40653
rect 56648 40601 56700 40653
rect 56859 40601 56911 40653
rect 57070 40601 57122 40653
rect 57281 40601 57333 40653
rect 48943 40509 48995 40515
rect 49154 40509 49206 40515
rect 49365 40509 49417 40515
rect 49576 40509 49628 40515
rect 49787 40509 49839 40515
rect 33057 40422 33109 40425
rect 33237 40422 33289 40425
rect 35332 40463 35384 40509
rect 35543 40463 35580 40509
rect 35580 40463 35595 40509
rect 35754 40463 35786 40509
rect 35786 40463 35806 40509
rect 35965 40463 35992 40509
rect 35992 40463 36017 40509
rect 36176 40463 36198 40509
rect 36198 40463 36228 40509
rect 37891 40465 37909 40509
rect 37909 40465 37943 40509
rect 38071 40465 38072 40509
rect 38072 40465 38123 40509
rect 33057 40376 33109 40422
rect 33237 40376 33289 40422
rect 33057 40373 33109 40376
rect 33237 40373 33289 40376
rect 33057 39974 33109 39977
rect 33237 39974 33289 39977
rect 33057 39928 33109 39974
rect 33237 39928 33289 39974
rect 33057 39925 33109 39928
rect 33237 39925 33289 39928
rect 29582 39701 29634 39753
rect 29793 39750 29845 39753
rect 29793 39704 29798 39750
rect 29798 39704 29844 39750
rect 29844 39704 29845 39750
rect 29793 39701 29845 39704
rect 30005 39701 30057 39753
rect 30216 39701 30268 39753
rect 34267 40198 34319 40215
rect 34447 40198 34499 40215
rect 34627 40198 34679 40215
rect 34267 40163 34302 40198
rect 34302 40163 34319 40198
rect 34447 40163 34451 40198
rect 34451 40163 34499 40198
rect 34627 40163 34658 40198
rect 34658 40163 34679 40198
rect 36678 40238 36697 40290
rect 36697 40238 36730 40290
rect 48943 40463 48984 40509
rect 48984 40463 48995 40509
rect 49154 40463 49190 40509
rect 49190 40463 49206 40509
rect 49365 40463 49396 40509
rect 49396 40463 49417 40509
rect 49576 40463 49602 40509
rect 49602 40463 49628 40509
rect 49787 40463 49839 40509
rect 39994 40340 40046 40392
rect 36961 40239 36971 40283
rect 36971 40239 37013 40283
rect 37172 40239 37206 40283
rect 37206 40239 37224 40283
rect 36961 40231 37013 40239
rect 37172 40231 37224 40239
rect 37384 40231 37436 40283
rect 37595 40231 37647 40283
rect 35332 40015 35384 40055
rect 35543 40015 35580 40055
rect 35580 40015 35595 40055
rect 35754 40015 35786 40055
rect 35786 40015 35806 40055
rect 35965 40015 35992 40055
rect 35992 40015 36017 40055
rect 36176 40015 36198 40055
rect 36198 40015 36228 40055
rect 37891 40015 37909 40043
rect 37909 40015 37943 40043
rect 38071 40015 38072 40043
rect 38072 40015 38123 40043
rect 35332 40003 35384 40015
rect 35543 40003 35595 40015
rect 35754 40003 35806 40015
rect 35965 40003 36017 40015
rect 36176 40003 36228 40015
rect 33819 39928 33833 39969
rect 33833 39928 33871 39969
rect 33999 39928 34039 39969
rect 34039 39928 34051 39969
rect 37891 39991 37943 40015
rect 38071 39991 38123 40015
rect 33819 39917 33871 39928
rect 33999 39917 34051 39928
rect 30854 39701 30906 39753
rect 31065 39701 31117 39753
rect 31276 39701 31328 39753
rect 31486 39750 31538 39753
rect 31697 39750 31749 39753
rect 31909 39750 31961 39753
rect 32120 39750 32172 39753
rect 32330 39750 32382 39753
rect 32541 39750 32593 39753
rect 32752 39750 32804 39753
rect 34284 39750 34336 39753
rect 34495 39750 34547 39753
rect 31486 39704 31538 39750
rect 31697 39704 31749 39750
rect 31909 39704 31961 39750
rect 32120 39704 32172 39750
rect 32330 39704 32382 39750
rect 32541 39704 32593 39750
rect 32752 39704 32804 39750
rect 34284 39704 34302 39750
rect 34302 39704 34336 39750
rect 34495 39704 34508 39750
rect 34508 39704 34547 39750
rect 31486 39701 31538 39704
rect 31697 39701 31749 39704
rect 31909 39701 31961 39704
rect 32120 39701 32172 39704
rect 32330 39701 32382 39704
rect 32541 39701 32593 39704
rect 32752 39701 32804 39704
rect 34284 39701 34336 39704
rect 34495 39701 34547 39704
rect 34707 39701 34759 39753
rect 34918 39701 34970 39753
rect 35220 39701 35272 39753
rect 35430 39701 35482 39753
rect 35641 39701 35693 39753
rect 35853 39701 35905 39753
rect 36064 39701 36116 39753
rect 36274 39701 36326 39753
rect 38330 39750 38382 39753
rect 38330 39704 38382 39750
rect 38330 39701 38382 39704
rect 38541 39701 38593 39753
rect 38752 39701 38804 39753
rect 39052 39750 39104 39753
rect 39232 39750 39284 39753
rect 39052 39704 39062 39750
rect 39062 39704 39104 39750
rect 39232 39704 39266 39750
rect 39266 39704 39284 39750
rect 39052 39701 39104 39704
rect 39232 39701 39284 39704
rect 33057 39526 33109 39529
rect 33237 39526 33289 39529
rect 33057 39480 33109 39526
rect 33237 39480 33289 39526
rect 33057 39477 33109 39480
rect 33237 39477 33289 39480
rect 33819 39526 33871 39537
rect 33999 39526 34051 39537
rect 33819 39485 33833 39526
rect 33833 39485 33871 39526
rect 33999 39485 34039 39526
rect 34039 39485 34051 39526
rect 35332 39439 35384 39451
rect 35543 39439 35595 39451
rect 35754 39439 35806 39451
rect 35965 39439 36017 39451
rect 36176 39439 36228 39451
rect 37891 39439 37943 39463
rect 38071 39439 38123 39463
rect 35332 39399 35384 39439
rect 35543 39399 35580 39439
rect 35580 39399 35595 39439
rect 35754 39399 35786 39439
rect 35786 39399 35806 39439
rect 35965 39399 35992 39439
rect 35992 39399 36017 39439
rect 36176 39399 36198 39439
rect 36198 39399 36228 39439
rect 37891 39411 37909 39439
rect 37909 39411 37943 39439
rect 38071 39411 38072 39439
rect 38072 39411 38123 39439
rect 34267 39256 34302 39291
rect 34302 39256 34319 39291
rect 34447 39256 34451 39291
rect 34451 39256 34499 39291
rect 34627 39256 34658 39291
rect 34658 39256 34679 39291
rect 34267 39239 34319 39256
rect 34447 39239 34499 39256
rect 34627 39239 34679 39256
rect 33057 39078 33109 39081
rect 33237 39078 33289 39081
rect 33057 39032 33109 39078
rect 33237 39032 33289 39078
rect 33057 39029 33109 39032
rect 33237 39029 33289 39032
rect 36678 39164 36697 39216
rect 36697 39164 36730 39216
rect 36961 39215 37013 39223
rect 37172 39215 37224 39223
rect 36961 39171 36971 39215
rect 36971 39171 37013 39215
rect 37172 39171 37206 39215
rect 37206 39171 37224 39215
rect 37384 39171 37436 39223
rect 37595 39171 37647 39223
rect 39994 40154 40046 40206
rect 39775 39974 39827 39991
rect 39775 39939 39786 39974
rect 39786 39939 39827 39974
rect 43445 40170 43497 40222
rect 41935 39939 41987 39991
rect 46731 40279 46783 40331
rect 48596 40325 48648 40377
rect 51835 40422 51887 40447
rect 52015 40422 52067 40447
rect 51835 40395 51887 40422
rect 52015 40395 52067 40422
rect 44939 40198 44991 40215
rect 45151 40198 45203 40215
rect 44939 40163 44971 40198
rect 44971 40163 44991 40198
rect 45151 40163 45197 40198
rect 45197 40163 45203 40198
rect 48596 40107 48648 40159
rect 50300 40163 50352 40215
rect 50511 40198 50563 40215
rect 50511 40163 50513 40198
rect 50513 40163 50563 40198
rect 50722 40163 50774 40215
rect 48943 40015 48984 40052
rect 48984 40015 48995 40052
rect 49154 40015 49190 40052
rect 49190 40015 49206 40052
rect 49365 40015 49396 40052
rect 49396 40015 49417 40052
rect 49576 40015 49602 40052
rect 49602 40015 49628 40052
rect 49787 40015 49839 40052
rect 48943 40000 48995 40015
rect 49154 40000 49206 40015
rect 49365 40000 49417 40015
rect 49576 40000 49628 40015
rect 49787 40000 49839 40015
rect 51073 39974 51125 39977
rect 51253 39974 51305 39977
rect 51073 39928 51086 39974
rect 51086 39928 51125 39974
rect 51253 39928 51292 39974
rect 51292 39928 51305 39974
rect 51073 39925 51125 39928
rect 51253 39925 51305 39928
rect 51835 39974 51887 39984
rect 52015 39974 52067 39984
rect 51835 39932 51887 39974
rect 52015 39932 52067 39974
rect 40253 39701 40305 39753
rect 40433 39701 40485 39753
rect 43790 39701 43842 39753
rect 44001 39701 44053 39753
rect 44213 39750 44265 39753
rect 44213 39704 44236 39750
rect 44236 39704 44265 39750
rect 44213 39701 44265 39704
rect 44424 39701 44476 39753
rect 44834 39750 44886 39753
rect 45045 39750 45097 39753
rect 45256 39750 45308 39753
rect 44834 39704 44858 39750
rect 44858 39704 44886 39750
rect 45045 39704 45084 39750
rect 45084 39704 45097 39750
rect 45256 39704 45264 39750
rect 45264 39704 45308 39750
rect 44834 39701 44886 39704
rect 45045 39701 45097 39704
rect 45256 39701 45308 39704
rect 48838 39701 48890 39753
rect 49048 39701 49100 39753
rect 49259 39701 49311 39753
rect 49471 39701 49523 39753
rect 49682 39701 49734 39753
rect 49892 39701 49944 39753
rect 50346 39701 50398 39753
rect 50557 39750 50609 39753
rect 50768 39750 50820 39753
rect 52316 39750 52368 39753
rect 52527 39750 52579 39753
rect 52738 39750 52790 39753
rect 52948 39750 53000 39753
rect 53159 39750 53211 39753
rect 53371 39750 53423 39753
rect 53582 39750 53634 39753
rect 50557 39704 50571 39750
rect 50571 39704 50609 39750
rect 50768 39704 50777 39750
rect 50777 39704 50820 39750
rect 52316 39704 52368 39750
rect 52527 39704 52579 39750
rect 52738 39704 52790 39750
rect 52948 39704 53000 39750
rect 53159 39704 53211 39750
rect 53371 39704 53423 39750
rect 53582 39704 53634 39750
rect 50557 39701 50609 39704
rect 50768 39701 50820 39704
rect 39775 39480 39786 39515
rect 39786 39480 39827 39515
rect 39775 39463 39827 39480
rect 39994 39248 40046 39300
rect 39994 39062 40046 39114
rect 52316 39701 52368 39704
rect 52527 39701 52579 39704
rect 52738 39701 52790 39704
rect 52948 39701 53000 39704
rect 53159 39701 53211 39704
rect 53371 39701 53423 39704
rect 53582 39701 53634 39704
rect 53792 39701 53844 39753
rect 54003 39701 54055 39753
rect 54214 39701 54266 39753
rect 54855 39701 54907 39753
rect 55066 39701 55118 39753
rect 55278 39750 55330 39753
rect 55278 39704 55279 39750
rect 55279 39704 55325 39750
rect 55325 39704 55330 39750
rect 55278 39701 55330 39704
rect 55489 39701 55541 39753
rect 41935 39463 41987 39515
rect 51073 39526 51125 39529
rect 51253 39526 51305 39529
rect 43445 39232 43497 39284
rect 51073 39480 51086 39526
rect 51086 39480 51125 39526
rect 51253 39480 51292 39526
rect 51292 39480 51305 39526
rect 48943 39439 48995 39454
rect 49154 39439 49206 39454
rect 49365 39439 49417 39454
rect 49576 39439 49628 39454
rect 49787 39439 49839 39454
rect 48943 39402 48984 39439
rect 48984 39402 48995 39439
rect 49154 39402 49190 39439
rect 49190 39402 49206 39439
rect 49365 39402 49396 39439
rect 49396 39402 49417 39439
rect 49576 39402 49602 39439
rect 49602 39402 49628 39439
rect 49787 39402 49839 39439
rect 51073 39477 51125 39480
rect 51253 39477 51305 39480
rect 44939 39256 44971 39291
rect 44971 39256 44991 39291
rect 45151 39256 45197 39291
rect 45197 39256 45203 39291
rect 48596 39295 48648 39347
rect 44939 39239 44991 39256
rect 45151 39239 45203 39256
rect 47108 39123 47160 39175
rect 50300 39239 50352 39291
rect 50511 39256 50513 39291
rect 50513 39256 50563 39291
rect 50511 39239 50563 39256
rect 50722 39239 50774 39291
rect 48596 39077 48648 39129
rect 51835 39480 51887 39522
rect 52015 39480 52067 39522
rect 51835 39470 51887 39480
rect 52015 39470 52067 39480
rect 35332 38945 35384 38991
rect 35543 38945 35580 38991
rect 35580 38945 35595 38991
rect 35754 38945 35786 38991
rect 35786 38945 35806 38991
rect 35965 38945 35992 38991
rect 35992 38945 36017 38991
rect 36176 38945 36198 38991
rect 36198 38945 36228 38991
rect 37891 38945 37909 38989
rect 37909 38945 37943 38989
rect 38071 38945 38072 38989
rect 38072 38945 38123 38989
rect 48943 38945 48984 38991
rect 48984 38945 48995 38991
rect 49154 38945 49190 38991
rect 49190 38945 49206 38991
rect 49365 38945 49396 38991
rect 49396 38945 49417 38991
rect 49576 38945 49602 38991
rect 49602 38945 49628 38991
rect 49787 38945 49839 38991
rect 51835 39032 51887 39059
rect 52015 39032 52067 39059
rect 51835 39007 51887 39032
rect 52015 39007 52067 39032
rect 35332 38939 35384 38945
rect 35543 38939 35595 38945
rect 35754 38939 35806 38945
rect 35965 38939 36017 38945
rect 36176 38939 36228 38945
rect 37891 38937 37943 38945
rect 38071 38937 38123 38945
rect 27790 38801 27842 38853
rect 28001 38801 28053 38853
rect 28212 38801 28264 38853
rect 28423 38801 28475 38853
rect 28634 38801 28686 38853
rect 28845 38850 28897 38853
rect 28845 38804 28856 38850
rect 28856 38804 28897 38850
rect 28845 38801 28897 38804
rect 29056 38801 29108 38853
rect 29582 38801 29634 38853
rect 29793 38850 29845 38853
rect 29793 38804 29798 38850
rect 29798 38804 29844 38850
rect 29844 38804 29845 38850
rect 29793 38801 29845 38804
rect 30005 38801 30057 38853
rect 30216 38801 30268 38853
rect 30854 38801 30906 38853
rect 31065 38801 31117 38853
rect 31276 38801 31328 38853
rect 31486 38801 31538 38853
rect 31697 38801 31749 38853
rect 31909 38801 31961 38853
rect 32120 38801 32172 38853
rect 32330 38801 32382 38853
rect 32541 38801 32593 38853
rect 32752 38801 32804 38853
rect 48943 38939 48995 38945
rect 49154 38939 49206 38945
rect 49365 38939 49417 38945
rect 49576 38939 49628 38945
rect 49787 38939 49839 38945
rect 34755 38801 34807 38853
rect 34935 38850 34987 38853
rect 34935 38804 34962 38850
rect 34962 38804 34987 38850
rect 34935 38801 34987 38804
rect 50138 38850 50190 38853
rect 50138 38804 50160 38850
rect 50160 38804 50190 38850
rect 50138 38801 50190 38804
rect 50318 38801 50370 38853
rect 35332 38709 35384 38715
rect 35543 38709 35595 38715
rect 35754 38709 35806 38715
rect 35965 38709 36017 38715
rect 36176 38709 36228 38715
rect 37891 38709 37943 38717
rect 38071 38709 38123 38717
rect 52316 38801 52368 38853
rect 52527 38801 52579 38853
rect 52738 38801 52790 38853
rect 52948 38801 53000 38853
rect 53159 38801 53211 38853
rect 53371 38801 53423 38853
rect 53582 38801 53634 38853
rect 53792 38801 53844 38853
rect 54003 38801 54055 38853
rect 54214 38801 54266 38853
rect 54855 38801 54907 38853
rect 55066 38801 55118 38853
rect 55278 38850 55330 38853
rect 55278 38804 55279 38850
rect 55279 38804 55325 38850
rect 55325 38804 55330 38850
rect 55278 38801 55330 38804
rect 55489 38801 55541 38853
rect 56015 38801 56067 38853
rect 56226 38850 56278 38853
rect 56226 38804 56267 38850
rect 56267 38804 56278 38850
rect 56226 38801 56278 38804
rect 56437 38801 56489 38853
rect 56648 38801 56700 38853
rect 56859 38801 56911 38853
rect 57070 38801 57122 38853
rect 57281 38801 57333 38853
rect 48943 38709 48995 38715
rect 49154 38709 49206 38715
rect 49365 38709 49417 38715
rect 49576 38709 49628 38715
rect 49787 38709 49839 38715
rect 33057 38622 33109 38625
rect 33237 38622 33289 38625
rect 35332 38663 35384 38709
rect 35543 38663 35580 38709
rect 35580 38663 35595 38709
rect 35754 38663 35786 38709
rect 35786 38663 35806 38709
rect 35965 38663 35992 38709
rect 35992 38663 36017 38709
rect 36176 38663 36198 38709
rect 36198 38663 36228 38709
rect 37891 38665 37909 38709
rect 37909 38665 37943 38709
rect 38071 38665 38072 38709
rect 38072 38665 38123 38709
rect 33057 38576 33109 38622
rect 33237 38576 33289 38622
rect 33057 38573 33109 38576
rect 33237 38573 33289 38576
rect 33057 38174 33109 38177
rect 33237 38174 33289 38177
rect 33057 38128 33109 38174
rect 33237 38128 33289 38174
rect 33057 38125 33109 38128
rect 33237 38125 33289 38128
rect 29582 37901 29634 37953
rect 29793 37950 29845 37953
rect 29793 37904 29798 37950
rect 29798 37904 29844 37950
rect 29844 37904 29845 37950
rect 29793 37901 29845 37904
rect 30005 37901 30057 37953
rect 30216 37901 30268 37953
rect 34267 38398 34319 38415
rect 34447 38398 34499 38415
rect 34627 38398 34679 38415
rect 34267 38363 34302 38398
rect 34302 38363 34319 38398
rect 34447 38363 34451 38398
rect 34451 38363 34499 38398
rect 34627 38363 34658 38398
rect 34658 38363 34679 38398
rect 36678 38438 36697 38490
rect 36697 38438 36730 38490
rect 48943 38663 48984 38709
rect 48984 38663 48995 38709
rect 49154 38663 49190 38709
rect 49190 38663 49206 38709
rect 49365 38663 49396 38709
rect 49396 38663 49417 38709
rect 49576 38663 49602 38709
rect 49602 38663 49628 38709
rect 49787 38663 49839 38709
rect 39994 38540 40046 38592
rect 36961 38439 36971 38483
rect 36971 38439 37013 38483
rect 37172 38439 37206 38483
rect 37206 38439 37224 38483
rect 36961 38431 37013 38439
rect 37172 38431 37224 38439
rect 37384 38431 37436 38483
rect 37595 38431 37647 38483
rect 35332 38215 35384 38255
rect 35543 38215 35580 38255
rect 35580 38215 35595 38255
rect 35754 38215 35786 38255
rect 35786 38215 35806 38255
rect 35965 38215 35992 38255
rect 35992 38215 36017 38255
rect 36176 38215 36198 38255
rect 36198 38215 36228 38255
rect 37891 38215 37909 38243
rect 37909 38215 37943 38243
rect 38071 38215 38072 38243
rect 38072 38215 38123 38243
rect 35332 38203 35384 38215
rect 35543 38203 35595 38215
rect 35754 38203 35806 38215
rect 35965 38203 36017 38215
rect 36176 38203 36228 38215
rect 33819 38128 33833 38169
rect 33833 38128 33871 38169
rect 33999 38128 34039 38169
rect 34039 38128 34051 38169
rect 37891 38191 37943 38215
rect 38071 38191 38123 38215
rect 33819 38117 33871 38128
rect 33999 38117 34051 38128
rect 30854 37901 30906 37953
rect 31065 37901 31117 37953
rect 31276 37901 31328 37953
rect 31486 37950 31538 37953
rect 31697 37950 31749 37953
rect 31909 37950 31961 37953
rect 32120 37950 32172 37953
rect 32330 37950 32382 37953
rect 32541 37950 32593 37953
rect 32752 37950 32804 37953
rect 34284 37950 34336 37953
rect 34495 37950 34547 37953
rect 31486 37904 31538 37950
rect 31697 37904 31749 37950
rect 31909 37904 31961 37950
rect 32120 37904 32172 37950
rect 32330 37904 32382 37950
rect 32541 37904 32593 37950
rect 32752 37904 32804 37950
rect 34284 37904 34302 37950
rect 34302 37904 34336 37950
rect 34495 37904 34508 37950
rect 34508 37904 34547 37950
rect 31486 37901 31538 37904
rect 31697 37901 31749 37904
rect 31909 37901 31961 37904
rect 32120 37901 32172 37904
rect 32330 37901 32382 37904
rect 32541 37901 32593 37904
rect 32752 37901 32804 37904
rect 34284 37901 34336 37904
rect 34495 37901 34547 37904
rect 34707 37901 34759 37953
rect 34918 37901 34970 37953
rect 35220 37901 35272 37953
rect 35430 37901 35482 37953
rect 35641 37901 35693 37953
rect 35853 37901 35905 37953
rect 36064 37901 36116 37953
rect 36274 37901 36326 37953
rect 38330 37950 38382 37953
rect 38330 37904 38382 37950
rect 38330 37901 38382 37904
rect 38541 37901 38593 37953
rect 38752 37901 38804 37953
rect 39052 37950 39104 37953
rect 39232 37950 39284 37953
rect 39052 37904 39062 37950
rect 39062 37904 39104 37950
rect 39232 37904 39266 37950
rect 39266 37904 39284 37950
rect 39052 37901 39104 37904
rect 39232 37901 39284 37904
rect 33057 37726 33109 37729
rect 33237 37726 33289 37729
rect 33057 37680 33109 37726
rect 33237 37680 33289 37726
rect 33057 37677 33109 37680
rect 33237 37677 33289 37680
rect 33819 37726 33871 37737
rect 33999 37726 34051 37737
rect 33819 37685 33833 37726
rect 33833 37685 33871 37726
rect 33999 37685 34039 37726
rect 34039 37685 34051 37726
rect 35332 37639 35384 37651
rect 35543 37639 35595 37651
rect 35754 37639 35806 37651
rect 35965 37639 36017 37651
rect 36176 37639 36228 37651
rect 37891 37639 37943 37663
rect 38071 37639 38123 37663
rect 35332 37599 35384 37639
rect 35543 37599 35580 37639
rect 35580 37599 35595 37639
rect 35754 37599 35786 37639
rect 35786 37599 35806 37639
rect 35965 37599 35992 37639
rect 35992 37599 36017 37639
rect 36176 37599 36198 37639
rect 36198 37599 36228 37639
rect 37891 37611 37909 37639
rect 37909 37611 37943 37639
rect 38071 37611 38072 37639
rect 38072 37611 38123 37639
rect 34267 37456 34302 37491
rect 34302 37456 34319 37491
rect 34447 37456 34451 37491
rect 34451 37456 34499 37491
rect 34627 37456 34658 37491
rect 34658 37456 34679 37491
rect 34267 37439 34319 37456
rect 34447 37439 34499 37456
rect 34627 37439 34679 37456
rect 33057 37278 33109 37281
rect 33237 37278 33289 37281
rect 33057 37232 33109 37278
rect 33237 37232 33289 37278
rect 33057 37229 33109 37232
rect 33237 37229 33289 37232
rect 36678 37364 36697 37416
rect 36697 37364 36730 37416
rect 36961 37415 37013 37423
rect 37172 37415 37224 37423
rect 36961 37371 36971 37415
rect 36971 37371 37013 37415
rect 37172 37371 37206 37415
rect 37206 37371 37224 37415
rect 37384 37371 37436 37423
rect 37595 37371 37647 37423
rect 39994 38354 40046 38406
rect 39775 38174 39827 38191
rect 39775 38139 39786 38174
rect 39786 38139 39827 38174
rect 43445 38370 43497 38422
rect 41935 38139 41987 38191
rect 47486 38479 47538 38531
rect 48596 38525 48648 38577
rect 51835 38622 51887 38647
rect 52015 38622 52067 38647
rect 51835 38595 51887 38622
rect 52015 38595 52067 38622
rect 44939 38398 44991 38415
rect 45151 38398 45203 38415
rect 44939 38363 44971 38398
rect 44971 38363 44991 38398
rect 45151 38363 45197 38398
rect 45197 38363 45203 38398
rect 48596 38307 48648 38359
rect 50300 38363 50352 38415
rect 50511 38398 50563 38415
rect 50511 38363 50513 38398
rect 50513 38363 50563 38398
rect 50722 38363 50774 38415
rect 48943 38215 48984 38252
rect 48984 38215 48995 38252
rect 49154 38215 49190 38252
rect 49190 38215 49206 38252
rect 49365 38215 49396 38252
rect 49396 38215 49417 38252
rect 49576 38215 49602 38252
rect 49602 38215 49628 38252
rect 49787 38215 49839 38252
rect 48943 38200 48995 38215
rect 49154 38200 49206 38215
rect 49365 38200 49417 38215
rect 49576 38200 49628 38215
rect 49787 38200 49839 38215
rect 51073 38174 51125 38177
rect 51253 38174 51305 38177
rect 51073 38128 51086 38174
rect 51086 38128 51125 38174
rect 51253 38128 51292 38174
rect 51292 38128 51305 38174
rect 51073 38125 51125 38128
rect 51253 38125 51305 38128
rect 51835 38174 51887 38184
rect 52015 38174 52067 38184
rect 51835 38132 51887 38174
rect 52015 38132 52067 38174
rect 40253 37901 40305 37953
rect 40433 37901 40485 37953
rect 43790 37901 43842 37953
rect 44001 37901 44053 37953
rect 44213 37950 44265 37953
rect 44213 37904 44236 37950
rect 44236 37904 44265 37950
rect 44213 37901 44265 37904
rect 44424 37901 44476 37953
rect 44834 37950 44886 37953
rect 45045 37950 45097 37953
rect 45256 37950 45308 37953
rect 44834 37904 44858 37950
rect 44858 37904 44886 37950
rect 45045 37904 45084 37950
rect 45084 37904 45097 37950
rect 45256 37904 45264 37950
rect 45264 37904 45308 37950
rect 44834 37901 44886 37904
rect 45045 37901 45097 37904
rect 45256 37901 45308 37904
rect 48838 37901 48890 37953
rect 49048 37901 49100 37953
rect 49259 37901 49311 37953
rect 49471 37901 49523 37953
rect 49682 37901 49734 37953
rect 49892 37901 49944 37953
rect 50346 37901 50398 37953
rect 50557 37950 50609 37953
rect 50768 37950 50820 37953
rect 52316 37950 52368 37953
rect 52527 37950 52579 37953
rect 52738 37950 52790 37953
rect 52948 37950 53000 37953
rect 53159 37950 53211 37953
rect 53371 37950 53423 37953
rect 53582 37950 53634 37953
rect 50557 37904 50571 37950
rect 50571 37904 50609 37950
rect 50768 37904 50777 37950
rect 50777 37904 50820 37950
rect 52316 37904 52368 37950
rect 52527 37904 52579 37950
rect 52738 37904 52790 37950
rect 52948 37904 53000 37950
rect 53159 37904 53211 37950
rect 53371 37904 53423 37950
rect 53582 37904 53634 37950
rect 50557 37901 50609 37904
rect 50768 37901 50820 37904
rect 39775 37680 39786 37715
rect 39786 37680 39827 37715
rect 39775 37663 39827 37680
rect 39994 37448 40046 37500
rect 39994 37262 40046 37314
rect 52316 37901 52368 37904
rect 52527 37901 52579 37904
rect 52738 37901 52790 37904
rect 52948 37901 53000 37904
rect 53159 37901 53211 37904
rect 53371 37901 53423 37904
rect 53582 37901 53634 37904
rect 53792 37901 53844 37953
rect 54003 37901 54055 37953
rect 54214 37901 54266 37953
rect 54855 37901 54907 37953
rect 55066 37901 55118 37953
rect 55278 37950 55330 37953
rect 55278 37904 55279 37950
rect 55279 37904 55325 37950
rect 55325 37904 55330 37950
rect 55278 37901 55330 37904
rect 55489 37901 55541 37953
rect 41935 37663 41987 37715
rect 51073 37726 51125 37729
rect 51253 37726 51305 37729
rect 43445 37432 43497 37484
rect 51073 37680 51086 37726
rect 51086 37680 51125 37726
rect 51253 37680 51292 37726
rect 51292 37680 51305 37726
rect 48943 37639 48995 37654
rect 49154 37639 49206 37654
rect 49365 37639 49417 37654
rect 49576 37639 49628 37654
rect 49787 37639 49839 37654
rect 48943 37602 48984 37639
rect 48984 37602 48995 37639
rect 49154 37602 49190 37639
rect 49190 37602 49206 37639
rect 49365 37602 49396 37639
rect 49396 37602 49417 37639
rect 49576 37602 49602 37639
rect 49602 37602 49628 37639
rect 49787 37602 49839 37639
rect 51073 37677 51125 37680
rect 51253 37677 51305 37680
rect 44939 37456 44971 37491
rect 44971 37456 44991 37491
rect 45151 37456 45197 37491
rect 45197 37456 45203 37491
rect 48596 37495 48648 37547
rect 44939 37439 44991 37456
rect 45151 37439 45203 37456
rect 47864 37323 47916 37375
rect 50300 37439 50352 37491
rect 50511 37456 50513 37491
rect 50513 37456 50563 37491
rect 50511 37439 50563 37456
rect 50722 37439 50774 37491
rect 48596 37277 48648 37329
rect 51835 37680 51887 37722
rect 52015 37680 52067 37722
rect 51835 37670 51887 37680
rect 52015 37670 52067 37680
rect 35332 37145 35384 37191
rect 35543 37145 35580 37191
rect 35580 37145 35595 37191
rect 35754 37145 35786 37191
rect 35786 37145 35806 37191
rect 35965 37145 35992 37191
rect 35992 37145 36017 37191
rect 36176 37145 36198 37191
rect 36198 37145 36228 37191
rect 37891 37145 37909 37189
rect 37909 37145 37943 37189
rect 38071 37145 38072 37189
rect 38072 37145 38123 37189
rect 48943 37145 48984 37191
rect 48984 37145 48995 37191
rect 49154 37145 49190 37191
rect 49190 37145 49206 37191
rect 49365 37145 49396 37191
rect 49396 37145 49417 37191
rect 49576 37145 49602 37191
rect 49602 37145 49628 37191
rect 49787 37145 49839 37191
rect 51835 37232 51887 37259
rect 52015 37232 52067 37259
rect 51835 37207 51887 37232
rect 52015 37207 52067 37232
rect 35332 37139 35384 37145
rect 35543 37139 35595 37145
rect 35754 37139 35806 37145
rect 35965 37139 36017 37145
rect 36176 37139 36228 37145
rect 37891 37137 37943 37145
rect 38071 37137 38123 37145
rect 27790 37001 27842 37053
rect 28001 37001 28053 37053
rect 28212 37001 28264 37053
rect 28423 37001 28475 37053
rect 28634 37001 28686 37053
rect 28845 37050 28897 37053
rect 28845 37004 28856 37050
rect 28856 37004 28897 37050
rect 28845 37001 28897 37004
rect 29056 37001 29108 37053
rect 29582 37001 29634 37053
rect 29793 37050 29845 37053
rect 29793 37004 29798 37050
rect 29798 37004 29844 37050
rect 29844 37004 29845 37050
rect 29793 37001 29845 37004
rect 30005 37001 30057 37053
rect 30216 37001 30268 37053
rect 30854 37001 30906 37053
rect 31065 37001 31117 37053
rect 31276 37001 31328 37053
rect 31486 37001 31538 37053
rect 31697 37001 31749 37053
rect 31909 37001 31961 37053
rect 32120 37001 32172 37053
rect 32330 37001 32382 37053
rect 32541 37001 32593 37053
rect 32752 37001 32804 37053
rect 48943 37139 48995 37145
rect 49154 37139 49206 37145
rect 49365 37139 49417 37145
rect 49576 37139 49628 37145
rect 49787 37139 49839 37145
rect 34755 37001 34807 37053
rect 34935 37050 34987 37053
rect 34935 37004 34962 37050
rect 34962 37004 34987 37050
rect 34935 37001 34987 37004
rect 50138 37050 50190 37053
rect 50138 37004 50160 37050
rect 50160 37004 50190 37050
rect 50138 37001 50190 37004
rect 50318 37001 50370 37053
rect 35332 36909 35384 36915
rect 35543 36909 35595 36915
rect 35754 36909 35806 36915
rect 35965 36909 36017 36915
rect 36176 36909 36228 36915
rect 37891 36909 37943 36917
rect 38071 36909 38123 36917
rect 52316 37001 52368 37053
rect 52527 37001 52579 37053
rect 52738 37001 52790 37053
rect 52948 37001 53000 37053
rect 53159 37001 53211 37053
rect 53371 37001 53423 37053
rect 53582 37001 53634 37053
rect 53792 37001 53844 37053
rect 54003 37001 54055 37053
rect 54214 37001 54266 37053
rect 54855 37001 54907 37053
rect 55066 37001 55118 37053
rect 55278 37050 55330 37053
rect 55278 37004 55279 37050
rect 55279 37004 55325 37050
rect 55325 37004 55330 37050
rect 55278 37001 55330 37004
rect 55489 37001 55541 37053
rect 56015 37001 56067 37053
rect 56226 37050 56278 37053
rect 56226 37004 56267 37050
rect 56267 37004 56278 37050
rect 56226 37001 56278 37004
rect 56437 37001 56489 37053
rect 56648 37001 56700 37053
rect 56859 37001 56911 37053
rect 57070 37001 57122 37053
rect 57281 37001 57333 37053
rect 48943 36909 48995 36915
rect 49154 36909 49206 36915
rect 49365 36909 49417 36915
rect 49576 36909 49628 36915
rect 49787 36909 49839 36915
rect 33057 36822 33109 36825
rect 33237 36822 33289 36825
rect 35332 36863 35384 36909
rect 35543 36863 35580 36909
rect 35580 36863 35595 36909
rect 35754 36863 35786 36909
rect 35786 36863 35806 36909
rect 35965 36863 35992 36909
rect 35992 36863 36017 36909
rect 36176 36863 36198 36909
rect 36198 36863 36228 36909
rect 37891 36865 37909 36909
rect 37909 36865 37943 36909
rect 38071 36865 38072 36909
rect 38072 36865 38123 36909
rect 33057 36776 33109 36822
rect 33237 36776 33289 36822
rect 33057 36773 33109 36776
rect 33237 36773 33289 36776
rect 33057 36374 33109 36377
rect 33237 36374 33289 36377
rect 33057 36328 33109 36374
rect 33237 36328 33289 36374
rect 33057 36325 33109 36328
rect 33237 36325 33289 36328
rect 29582 36101 29634 36153
rect 29793 36150 29845 36153
rect 29793 36104 29798 36150
rect 29798 36104 29844 36150
rect 29844 36104 29845 36150
rect 29793 36101 29845 36104
rect 30005 36101 30057 36153
rect 30216 36101 30268 36153
rect 34267 36598 34319 36615
rect 34447 36598 34499 36615
rect 34627 36598 34679 36615
rect 34267 36563 34302 36598
rect 34302 36563 34319 36598
rect 34447 36563 34451 36598
rect 34451 36563 34499 36598
rect 34627 36563 34658 36598
rect 34658 36563 34679 36598
rect 36678 36638 36697 36690
rect 36697 36638 36730 36690
rect 48943 36863 48984 36909
rect 48984 36863 48995 36909
rect 49154 36863 49190 36909
rect 49190 36863 49206 36909
rect 49365 36863 49396 36909
rect 49396 36863 49417 36909
rect 49576 36863 49602 36909
rect 49602 36863 49628 36909
rect 49787 36863 49839 36909
rect 39994 36740 40046 36792
rect 36961 36639 36971 36683
rect 36971 36639 37013 36683
rect 37172 36639 37206 36683
rect 37206 36639 37224 36683
rect 36961 36631 37013 36639
rect 37172 36631 37224 36639
rect 37384 36631 37436 36683
rect 37595 36631 37647 36683
rect 35332 36415 35384 36455
rect 35543 36415 35580 36455
rect 35580 36415 35595 36455
rect 35754 36415 35786 36455
rect 35786 36415 35806 36455
rect 35965 36415 35992 36455
rect 35992 36415 36017 36455
rect 36176 36415 36198 36455
rect 36198 36415 36228 36455
rect 37891 36415 37909 36443
rect 37909 36415 37943 36443
rect 38071 36415 38072 36443
rect 38072 36415 38123 36443
rect 35332 36403 35384 36415
rect 35543 36403 35595 36415
rect 35754 36403 35806 36415
rect 35965 36403 36017 36415
rect 36176 36403 36228 36415
rect 33819 36328 33833 36369
rect 33833 36328 33871 36369
rect 33999 36328 34039 36369
rect 34039 36328 34051 36369
rect 37891 36391 37943 36415
rect 38071 36391 38123 36415
rect 33819 36317 33871 36328
rect 33999 36317 34051 36328
rect 30854 36101 30906 36153
rect 31065 36101 31117 36153
rect 31276 36101 31328 36153
rect 31486 36150 31538 36153
rect 31697 36150 31749 36153
rect 31909 36150 31961 36153
rect 32120 36150 32172 36153
rect 32330 36150 32382 36153
rect 32541 36150 32593 36153
rect 32752 36150 32804 36153
rect 34284 36150 34336 36153
rect 34495 36150 34547 36153
rect 31486 36104 31538 36150
rect 31697 36104 31749 36150
rect 31909 36104 31961 36150
rect 32120 36104 32172 36150
rect 32330 36104 32382 36150
rect 32541 36104 32593 36150
rect 32752 36104 32804 36150
rect 34284 36104 34302 36150
rect 34302 36104 34336 36150
rect 34495 36104 34508 36150
rect 34508 36104 34547 36150
rect 31486 36101 31538 36104
rect 31697 36101 31749 36104
rect 31909 36101 31961 36104
rect 32120 36101 32172 36104
rect 32330 36101 32382 36104
rect 32541 36101 32593 36104
rect 32752 36101 32804 36104
rect 34284 36101 34336 36104
rect 34495 36101 34547 36104
rect 34707 36101 34759 36153
rect 34918 36101 34970 36153
rect 35220 36101 35272 36153
rect 35430 36101 35482 36153
rect 35641 36101 35693 36153
rect 35853 36101 35905 36153
rect 36064 36101 36116 36153
rect 36274 36101 36326 36153
rect 38330 36150 38382 36153
rect 38330 36104 38382 36150
rect 38330 36101 38382 36104
rect 38541 36101 38593 36153
rect 38752 36101 38804 36153
rect 39052 36150 39104 36153
rect 39232 36150 39284 36153
rect 39052 36104 39062 36150
rect 39062 36104 39104 36150
rect 39232 36104 39266 36150
rect 39266 36104 39284 36150
rect 39052 36101 39104 36104
rect 39232 36101 39284 36104
rect 39994 36554 40046 36606
rect 39775 36374 39827 36391
rect 39775 36339 39786 36374
rect 39786 36339 39827 36374
rect 43445 36570 43497 36622
rect 41935 36339 41987 36391
rect 48241 36679 48293 36731
rect 48596 36725 48648 36777
rect 51835 36822 51887 36847
rect 52015 36822 52067 36847
rect 51835 36795 51887 36822
rect 52015 36795 52067 36822
rect 44939 36598 44991 36615
rect 45151 36598 45203 36615
rect 44939 36563 44971 36598
rect 44971 36563 44991 36598
rect 45151 36563 45197 36598
rect 45197 36563 45203 36598
rect 48596 36507 48648 36559
rect 50300 36563 50352 36615
rect 50511 36598 50563 36615
rect 50511 36563 50513 36598
rect 50513 36563 50563 36598
rect 50722 36563 50774 36615
rect 48943 36415 48984 36452
rect 48984 36415 48995 36452
rect 49154 36415 49190 36452
rect 49190 36415 49206 36452
rect 49365 36415 49396 36452
rect 49396 36415 49417 36452
rect 49576 36415 49602 36452
rect 49602 36415 49628 36452
rect 49787 36415 49839 36452
rect 48943 36400 48995 36415
rect 49154 36400 49206 36415
rect 49365 36400 49417 36415
rect 49576 36400 49628 36415
rect 49787 36400 49839 36415
rect 51073 36374 51125 36377
rect 51253 36374 51305 36377
rect 51073 36328 51086 36374
rect 51086 36328 51125 36374
rect 51253 36328 51292 36374
rect 51292 36328 51305 36374
rect 51073 36325 51125 36328
rect 51253 36325 51305 36328
rect 51835 36374 51887 36384
rect 52015 36374 52067 36384
rect 51835 36332 51887 36374
rect 52015 36332 52067 36374
rect 40253 36101 40305 36153
rect 40433 36101 40485 36153
rect 43790 36101 43842 36153
rect 44001 36101 44053 36153
rect 44213 36150 44265 36153
rect 44213 36104 44236 36150
rect 44236 36104 44265 36150
rect 44213 36101 44265 36104
rect 44424 36101 44476 36153
rect 44834 36150 44886 36153
rect 45045 36150 45097 36153
rect 45256 36150 45308 36153
rect 44834 36104 44858 36150
rect 44858 36104 44886 36150
rect 45045 36104 45084 36150
rect 45084 36104 45097 36150
rect 45256 36104 45264 36150
rect 45264 36104 45308 36150
rect 44834 36101 44886 36104
rect 45045 36101 45097 36104
rect 45256 36101 45308 36104
rect 48838 36101 48890 36153
rect 49048 36101 49100 36153
rect 49259 36101 49311 36153
rect 49471 36101 49523 36153
rect 49682 36101 49734 36153
rect 49892 36101 49944 36153
rect 50346 36101 50398 36153
rect 50557 36150 50609 36153
rect 50768 36150 50820 36153
rect 52316 36150 52368 36153
rect 52527 36150 52579 36153
rect 52738 36150 52790 36153
rect 52948 36150 53000 36153
rect 53159 36150 53211 36153
rect 53371 36150 53423 36153
rect 53582 36150 53634 36153
rect 50557 36104 50571 36150
rect 50571 36104 50609 36150
rect 50768 36104 50777 36150
rect 50777 36104 50820 36150
rect 52316 36104 52368 36150
rect 52527 36104 52579 36150
rect 52738 36104 52790 36150
rect 52948 36104 53000 36150
rect 53159 36104 53211 36150
rect 53371 36104 53423 36150
rect 53582 36104 53634 36150
rect 50557 36101 50609 36104
rect 50768 36101 50820 36104
rect 52316 36101 52368 36104
rect 52527 36101 52579 36104
rect 52738 36101 52790 36104
rect 52948 36101 53000 36104
rect 53159 36101 53211 36104
rect 53371 36101 53423 36104
rect 53582 36101 53634 36104
rect 53792 36101 53844 36153
rect 54003 36101 54055 36153
rect 54214 36101 54266 36153
rect 54855 36101 54907 36153
rect 55066 36101 55118 36153
rect 55278 36150 55330 36153
rect 55278 36104 55279 36150
rect 55279 36104 55325 36150
rect 55325 36104 55330 36150
rect 55278 36101 55330 36104
rect 55489 36101 55541 36153
rect 25346 34907 25398 34959
rect 25470 34907 25522 34959
rect 25594 34907 25646 34959
rect 25718 34907 25770 34959
rect 25842 34907 25894 34959
rect 25966 34907 26018 34959
rect 25346 34783 25398 34835
rect 25470 34783 25522 34835
rect 25594 34783 25646 34835
rect 25718 34783 25770 34835
rect 25842 34783 25894 34835
rect 25966 34783 26018 34835
rect 25346 34659 25398 34711
rect 25470 34659 25522 34711
rect 25594 34659 25646 34711
rect 25718 34659 25770 34711
rect 25842 34659 25894 34711
rect 25966 34659 26018 34711
rect 27469 34596 27729 34960
rect 58824 34927 58876 34979
rect 58948 34927 59000 34979
rect 59072 34927 59124 34979
rect 59196 34927 59248 34979
rect 59320 34927 59372 34979
rect 59444 34927 59496 34979
rect 58824 34803 58876 34855
rect 58948 34803 59000 34855
rect 59072 34803 59124 34855
rect 59196 34803 59248 34855
rect 59320 34803 59372 34855
rect 59444 34803 59496 34855
rect 58824 34679 58876 34731
rect 58948 34679 59000 34731
rect 59072 34679 59124 34731
rect 59196 34679 59248 34731
rect 59320 34679 59372 34731
rect 59444 34679 59496 34731
rect 26861 33380 26913 33432
rect 27073 33380 27125 33432
rect 26861 33163 26913 33215
rect 27073 33163 27125 33215
rect 26861 32945 26913 32997
rect 27073 32945 27125 32997
rect 26861 32727 26913 32779
rect 27073 32727 27125 32779
rect 26861 32510 26913 32562
rect 27073 32510 27125 32562
rect 26861 32292 26913 32344
rect 27073 32292 27125 32344
rect 26861 32075 26913 32127
rect 27073 32075 27125 32127
rect 26861 31857 26913 31909
rect 27073 31857 27125 31909
rect 26861 31639 26913 31691
rect 27073 31639 27125 31691
rect 26861 31422 26913 31474
rect 27073 31422 27125 31474
rect 26861 31204 26913 31256
rect 27073 31204 27125 31256
rect 26861 30986 26913 31038
rect 27073 30986 27125 31038
rect 26861 30769 26913 30821
rect 27073 30769 27125 30821
rect 26861 30551 26913 30603
rect 27073 30551 27125 30603
rect 26861 30334 26913 30386
rect 27073 30334 27125 30386
rect 26861 30116 26913 30168
rect 27073 30116 27125 30168
rect 26861 29898 26913 29950
rect 27073 29898 27125 29950
rect 26861 29681 26913 29733
rect 27073 29681 27125 29733
rect 26861 29463 26913 29515
rect 27073 29463 27125 29515
rect 26861 29245 26913 29297
rect 27073 29245 27125 29297
rect 26861 29028 26913 29080
rect 27073 29028 27125 29080
rect 26861 28810 26913 28862
rect 27073 28810 27125 28862
rect 26861 28592 26913 28644
rect 27073 28592 27125 28644
rect 26861 28375 26913 28427
rect 27073 28375 27125 28427
rect 26861 28157 26913 28209
rect 27073 28157 27125 28209
rect 26861 27940 26913 27992
rect 27073 27940 27125 27992
rect 26861 27722 26913 27774
rect 27073 27722 27125 27774
rect 26861 27504 26913 27556
rect 27073 27504 27125 27556
rect 26861 27287 26913 27339
rect 27073 27287 27125 27339
rect 26861 27069 26913 27121
rect 27073 27069 27125 27121
rect 26861 26851 26913 26903
rect 27073 26851 27125 26903
rect 26861 26634 26913 26686
rect 27073 26634 27125 26686
rect 26861 26416 26913 26468
rect 27073 26416 27125 26468
rect 26861 26198 26913 26250
rect 27073 26198 27125 26250
rect 26861 25981 26913 26033
rect 27073 25981 27125 26033
rect 26861 25763 26913 25815
rect 27073 25763 27125 25815
rect 26861 25546 26913 25598
rect 27073 25546 27125 25598
rect 26861 25328 26913 25380
rect 27073 25328 27125 25380
rect 26861 25110 26913 25162
rect 27073 25110 27125 25162
rect 26861 24893 26913 24945
rect 27073 24893 27125 24945
rect 26861 24675 26913 24727
rect 27073 24675 27125 24727
rect 26861 24457 26913 24509
rect 27073 24457 27125 24509
rect 26861 24240 26913 24292
rect 27073 24240 27125 24292
rect 26861 24022 26913 24074
rect 27073 24022 27125 24074
rect 26861 23805 26913 23857
rect 27073 23805 27125 23857
rect 26861 23587 26913 23639
rect 27073 23587 27125 23639
rect 26861 23369 26913 23421
rect 27073 23369 27125 23421
rect 26861 23152 26913 23204
rect 27073 23152 27125 23204
rect 26861 22934 26913 22986
rect 27073 22934 27125 22986
rect 26861 22716 26913 22768
rect 27073 22716 27125 22768
rect 26861 22499 26913 22551
rect 27073 22499 27125 22551
rect 26861 22281 26913 22333
rect 27073 22281 27125 22333
rect 26861 22063 26913 22115
rect 27073 22063 27125 22115
rect 26861 21846 26913 21898
rect 27073 21846 27125 21898
rect 26861 21628 26913 21680
rect 27073 21628 27125 21680
rect 26861 21411 26913 21463
rect 27073 21411 27125 21463
rect 26861 21193 26913 21245
rect 27073 21193 27125 21245
rect 26861 20975 26913 21027
rect 27073 20975 27125 21027
rect 26861 20758 26913 20810
rect 27073 20758 27125 20810
rect 26861 20540 26913 20592
rect 27073 20540 27125 20592
rect 26861 20322 26913 20374
rect 27073 20322 27125 20374
rect 26861 20105 26913 20157
rect 27073 20105 27125 20157
rect 26861 19887 26913 19939
rect 27073 19887 27125 19939
rect 26861 19670 26913 19722
rect 27073 19670 27125 19722
rect 26861 19452 26913 19504
rect 27073 19452 27125 19504
rect 26861 19234 26913 19286
rect 27073 19234 27125 19286
rect 26861 19016 26913 19068
rect 27073 19016 27125 19068
rect 26861 18799 26913 18851
rect 27073 18799 27125 18851
rect 26861 18581 26913 18633
rect 27073 18581 27125 18633
rect 26861 18364 26913 18416
rect 27073 18364 27125 18416
rect 26861 18146 26913 18198
rect 27073 18146 27125 18198
rect 26861 17928 26913 17980
rect 27073 17928 27125 17980
rect 26861 17711 26913 17763
rect 27073 17711 27125 17763
rect 26861 17493 26913 17545
rect 27073 17493 27125 17545
rect 26861 17275 26913 17327
rect 27073 17275 27125 17327
rect 26861 17058 26913 17110
rect 27073 17058 27125 17110
rect 26861 16840 26913 16892
rect 27073 16840 27125 16892
rect 26861 16623 26913 16675
rect 27073 16623 27125 16675
rect 26861 16405 26913 16457
rect 27073 16405 27125 16457
rect 26861 16187 26913 16239
rect 27073 16187 27125 16239
rect 26861 15970 26913 16022
rect 27073 15970 27125 16022
rect 26861 15752 26913 15804
rect 27073 15752 27125 15804
rect 26861 15534 26913 15586
rect 27073 15534 27125 15586
rect 26861 15317 26913 15369
rect 27073 15317 27125 15369
rect 26861 15099 26913 15151
rect 27073 15099 27125 15151
rect 26861 14881 26913 14933
rect 27073 14881 27125 14933
rect 26861 14664 26913 14716
rect 27073 14664 27125 14716
rect 26861 14446 26913 14498
rect 27073 14446 27125 14498
rect 26861 14229 26913 14281
rect 27073 14229 27125 14281
rect 26861 14011 26913 14063
rect 27073 14011 27125 14063
rect 26861 13793 26913 13845
rect 27073 13793 27125 13845
rect 26861 13576 26913 13628
rect 27073 13576 27125 13628
rect 26861 13358 26913 13410
rect 27073 13358 27125 13410
rect 26861 13140 26913 13192
rect 27073 13140 27125 13192
rect 26861 12923 26913 12975
rect 27073 12923 27125 12975
rect 26861 12705 26913 12757
rect 27073 12705 27125 12757
rect 26861 12488 26913 12540
rect 27073 12488 27125 12540
rect 26861 12270 26913 12322
rect 27073 12270 27125 12322
rect 26861 12052 26913 12104
rect 27073 12052 27125 12104
rect 26861 11835 26913 11887
rect 27073 11835 27125 11887
rect 26861 11617 26913 11669
rect 27073 11617 27125 11669
rect 26861 11399 26913 11451
rect 27073 11399 27125 11451
rect 26861 11182 26913 11234
rect 27073 11182 27125 11234
rect 26861 10964 26913 11016
rect 27073 10964 27125 11016
rect 26861 10746 26913 10798
rect 27073 10746 27125 10798
rect 26861 10529 26913 10581
rect 27073 10529 27125 10581
rect 26861 10311 26913 10363
rect 27073 10311 27125 10363
rect 26861 10094 26913 10146
rect 27073 10094 27125 10146
rect 26861 9876 26913 9928
rect 27073 9876 27125 9928
rect 26861 9658 26913 9710
rect 27073 9658 27125 9710
rect 26861 9441 26913 9493
rect 27073 9441 27125 9493
rect 26861 9223 26913 9275
rect 27073 9223 27125 9275
rect 26861 9005 26913 9057
rect 27073 9005 27125 9057
rect 26861 8788 26913 8840
rect 27073 8788 27125 8840
rect 26861 8570 26913 8622
rect 27073 8570 27125 8622
rect 26861 8352 26913 8404
rect 27073 8352 27125 8404
rect 26861 8135 26913 8187
rect 27073 8135 27125 8187
rect 26861 7917 26913 7969
rect 27073 7917 27125 7969
rect 26861 7700 26913 7752
rect 27073 7700 27125 7752
rect 26861 7482 26913 7534
rect 27073 7482 27125 7534
rect 26861 7264 26913 7316
rect 27073 7264 27125 7316
rect 26861 7047 26913 7099
rect 27073 7047 27125 7099
rect 26861 6829 26913 6881
rect 27073 6829 27125 6881
rect 26861 6611 26913 6663
rect 27073 6611 27125 6663
rect 26861 6394 26913 6446
rect 27073 6394 27125 6446
rect 26861 6176 26913 6228
rect 27073 6176 27125 6228
rect 26861 5959 26913 6011
rect 27073 5959 27125 6011
rect 26861 5741 26913 5793
rect 27073 5741 27125 5793
rect 26861 5523 26913 5575
rect 27073 5523 27125 5575
rect 26861 5306 26913 5358
rect 27073 5306 27125 5358
rect 26861 4535 26913 4587
rect 27073 4535 27125 4587
rect 26861 4318 26913 4370
rect 27073 4318 27125 4370
rect 26861 4100 26913 4152
rect 27073 4100 27125 4152
rect 26861 3882 26913 3934
rect 27073 3882 27125 3934
rect 26861 3665 26913 3717
rect 27073 3665 27125 3717
rect 27476 33380 27528 33432
rect 27688 33380 27740 33432
rect 27476 33163 27528 33215
rect 27688 33163 27740 33215
rect 27476 32945 27528 32997
rect 27688 32945 27740 32997
rect 27476 32727 27528 32779
rect 27688 32727 27740 32779
rect 27476 32510 27528 32562
rect 27688 32510 27740 32562
rect 27476 32292 27528 32344
rect 27688 32292 27740 32344
rect 27476 32075 27528 32127
rect 27688 32075 27740 32127
rect 27476 31857 27528 31909
rect 27688 31857 27740 31909
rect 27476 31639 27528 31691
rect 27688 31639 27740 31691
rect 27476 31422 27528 31474
rect 27688 31422 27740 31474
rect 27476 31204 27528 31256
rect 27688 31204 27740 31256
rect 27476 30986 27528 31038
rect 27688 30986 27740 31038
rect 27476 30769 27528 30821
rect 27688 30769 27740 30821
rect 27476 30551 27528 30603
rect 27688 30551 27740 30603
rect 27476 30334 27528 30386
rect 27688 30334 27740 30386
rect 27476 30116 27528 30168
rect 27688 30116 27740 30168
rect 27476 29898 27528 29950
rect 27688 29898 27740 29950
rect 27476 29681 27528 29733
rect 27688 29681 27740 29733
rect 27476 29463 27528 29515
rect 27688 29463 27740 29515
rect 27476 29245 27528 29297
rect 27688 29245 27740 29297
rect 27476 29028 27528 29080
rect 27688 29028 27740 29080
rect 27476 28810 27528 28862
rect 27688 28810 27740 28862
rect 27476 28592 27528 28644
rect 27688 28592 27740 28644
rect 27476 28375 27528 28427
rect 27688 28375 27740 28427
rect 27476 28157 27528 28209
rect 27688 28157 27740 28209
rect 27476 27940 27528 27992
rect 27688 27940 27740 27992
rect 27476 27722 27528 27774
rect 27688 27722 27740 27774
rect 27476 27504 27528 27556
rect 27688 27504 27740 27556
rect 27476 27287 27528 27339
rect 27688 27287 27740 27339
rect 27476 27069 27528 27121
rect 27688 27069 27740 27121
rect 27476 26851 27528 26903
rect 27688 26851 27740 26903
rect 27476 26634 27528 26686
rect 27688 26634 27740 26686
rect 27476 26416 27528 26468
rect 27688 26416 27740 26468
rect 27476 26198 27528 26250
rect 27688 26198 27740 26250
rect 27476 25981 27528 26033
rect 27688 25981 27740 26033
rect 27476 25763 27528 25815
rect 27688 25763 27740 25815
rect 27476 25546 27528 25598
rect 27688 25546 27740 25598
rect 27476 25328 27528 25380
rect 27688 25328 27740 25380
rect 27476 25110 27528 25162
rect 27688 25110 27740 25162
rect 27476 24893 27528 24945
rect 27688 24893 27740 24945
rect 27476 24675 27528 24727
rect 27688 24675 27740 24727
rect 27476 24457 27528 24509
rect 27688 24457 27740 24509
rect 27476 24240 27528 24292
rect 27688 24240 27740 24292
rect 27476 24022 27528 24074
rect 27688 24022 27740 24074
rect 27476 23805 27528 23857
rect 27688 23805 27740 23857
rect 27476 23587 27528 23639
rect 27688 23587 27740 23639
rect 27476 23369 27528 23421
rect 27688 23369 27740 23421
rect 27476 23152 27528 23204
rect 27688 23152 27740 23204
rect 27476 22934 27528 22986
rect 27688 22934 27740 22986
rect 27476 22716 27528 22768
rect 27688 22716 27740 22768
rect 27476 22499 27528 22551
rect 27688 22499 27740 22551
rect 27476 22281 27528 22333
rect 27688 22281 27740 22333
rect 27476 22063 27528 22115
rect 27688 22063 27740 22115
rect 27476 21846 27528 21898
rect 27688 21846 27740 21898
rect 27476 21628 27528 21680
rect 27688 21628 27740 21680
rect 27476 21411 27528 21463
rect 27688 21411 27740 21463
rect 27476 21193 27528 21245
rect 27688 21193 27740 21245
rect 27476 20975 27528 21027
rect 27688 20975 27740 21027
rect 27476 20758 27528 20810
rect 27688 20758 27740 20810
rect 27476 20540 27528 20592
rect 27688 20540 27740 20592
rect 27476 20322 27528 20374
rect 27688 20322 27740 20374
rect 27476 20105 27528 20157
rect 27688 20105 27740 20157
rect 27476 19887 27528 19939
rect 27688 19887 27740 19939
rect 27476 19670 27528 19722
rect 27688 19670 27740 19722
rect 27476 19452 27528 19504
rect 27688 19452 27740 19504
rect 27476 19234 27528 19286
rect 27688 19234 27740 19286
rect 27476 19016 27528 19068
rect 27688 19016 27740 19068
rect 27476 18799 27528 18851
rect 27688 18799 27740 18851
rect 27476 18581 27528 18633
rect 27688 18581 27740 18633
rect 27476 18364 27528 18416
rect 27688 18364 27740 18416
rect 27476 18146 27528 18198
rect 27688 18146 27740 18198
rect 27476 17928 27528 17980
rect 27688 17928 27740 17980
rect 27476 17711 27528 17763
rect 27688 17711 27740 17763
rect 27476 17493 27528 17545
rect 27688 17493 27740 17545
rect 27476 17275 27528 17327
rect 27688 17275 27740 17327
rect 27476 17058 27528 17110
rect 27688 17058 27740 17110
rect 27476 16840 27528 16892
rect 27688 16840 27740 16892
rect 27476 16623 27528 16675
rect 27688 16623 27740 16675
rect 27476 16405 27528 16457
rect 27688 16405 27740 16457
rect 27476 16187 27528 16239
rect 27688 16187 27740 16239
rect 27476 15970 27528 16022
rect 27688 15970 27740 16022
rect 27476 15752 27528 15804
rect 27688 15752 27740 15804
rect 27476 15534 27528 15586
rect 27688 15534 27740 15586
rect 27476 15317 27528 15369
rect 27688 15317 27740 15369
rect 27476 15099 27528 15151
rect 27688 15099 27740 15151
rect 27476 14881 27528 14933
rect 27688 14881 27740 14933
rect 27476 14664 27528 14716
rect 27688 14664 27740 14716
rect 27476 14446 27528 14498
rect 27688 14446 27740 14498
rect 27476 14229 27528 14281
rect 27688 14229 27740 14281
rect 27476 14011 27528 14063
rect 27688 14011 27740 14063
rect 27476 13793 27528 13845
rect 27688 13793 27740 13845
rect 27476 13576 27528 13628
rect 27688 13576 27740 13628
rect 27476 13358 27528 13410
rect 27688 13358 27740 13410
rect 27476 13140 27528 13192
rect 27688 13140 27740 13192
rect 27476 12923 27528 12975
rect 27688 12923 27740 12975
rect 27476 12705 27528 12757
rect 27688 12705 27740 12757
rect 27476 12488 27528 12540
rect 27688 12488 27740 12540
rect 27476 12270 27528 12322
rect 27688 12270 27740 12322
rect 27476 12052 27528 12104
rect 27688 12052 27740 12104
rect 27476 11835 27528 11887
rect 27688 11835 27740 11887
rect 27476 11617 27528 11669
rect 27688 11617 27740 11669
rect 27476 11399 27528 11451
rect 27688 11399 27740 11451
rect 27476 11182 27528 11234
rect 27688 11182 27740 11234
rect 27476 10964 27528 11016
rect 27688 10964 27740 11016
rect 27476 10746 27528 10798
rect 27688 10746 27740 10798
rect 27476 10529 27528 10581
rect 27688 10529 27740 10581
rect 27476 10311 27528 10363
rect 27688 10311 27740 10363
rect 27476 10094 27528 10146
rect 27688 10094 27740 10146
rect 27476 9876 27528 9928
rect 27688 9876 27740 9928
rect 27476 9658 27528 9710
rect 27688 9658 27740 9710
rect 27476 9441 27528 9493
rect 27688 9441 27740 9493
rect 27476 9223 27528 9275
rect 27688 9223 27740 9275
rect 27476 9005 27528 9057
rect 27688 9005 27740 9057
rect 27476 8788 27528 8840
rect 27688 8788 27740 8840
rect 27476 8570 27528 8622
rect 27688 8570 27740 8622
rect 27476 8352 27528 8404
rect 27688 8352 27740 8404
rect 27476 8135 27528 8187
rect 27688 8135 27740 8187
rect 27476 7917 27528 7969
rect 27688 7917 27740 7969
rect 27476 7700 27528 7752
rect 27688 7700 27740 7752
rect 27476 7482 27528 7534
rect 27688 7482 27740 7534
rect 27476 7264 27528 7316
rect 27688 7264 27740 7316
rect 27476 7047 27528 7099
rect 27688 7047 27740 7099
rect 27476 6829 27528 6881
rect 27688 6829 27740 6881
rect 27476 6611 27528 6663
rect 27688 6611 27740 6663
rect 27476 6394 27528 6446
rect 27688 6394 27740 6446
rect 57383 33380 57435 33432
rect 57595 33380 57647 33432
rect 57383 33163 57435 33215
rect 57595 33163 57647 33215
rect 57383 32945 57435 32997
rect 57595 32945 57647 32997
rect 57383 32727 57435 32779
rect 57595 32727 57647 32779
rect 57383 32510 57435 32562
rect 57595 32510 57647 32562
rect 57383 32292 57435 32344
rect 57595 32292 57647 32344
rect 57383 32075 57435 32127
rect 57595 32075 57647 32127
rect 57383 31857 57435 31909
rect 57595 31857 57647 31909
rect 57383 31639 57435 31691
rect 57595 31639 57647 31691
rect 57383 31422 57435 31474
rect 57595 31422 57647 31474
rect 57383 31204 57435 31256
rect 57595 31204 57647 31256
rect 57383 30986 57435 31038
rect 57595 30986 57647 31038
rect 57383 30769 57435 30821
rect 57595 30769 57647 30821
rect 57383 30551 57435 30603
rect 57595 30551 57647 30603
rect 57383 30334 57435 30386
rect 57595 30334 57647 30386
rect 57383 30116 57435 30168
rect 57595 30116 57647 30168
rect 57383 29898 57435 29950
rect 57595 29898 57647 29950
rect 57383 29681 57435 29733
rect 57595 29681 57647 29733
rect 57383 29463 57435 29515
rect 57595 29463 57647 29515
rect 57383 29245 57435 29297
rect 57595 29245 57647 29297
rect 57383 29028 57435 29080
rect 57595 29028 57647 29080
rect 57383 28810 57435 28862
rect 57595 28810 57647 28862
rect 57383 28592 57435 28644
rect 57595 28592 57647 28644
rect 57383 28375 57435 28427
rect 57595 28375 57647 28427
rect 57383 28157 57435 28209
rect 57595 28157 57647 28209
rect 57383 27940 57435 27992
rect 57595 27940 57647 27992
rect 57383 27722 57435 27774
rect 57595 27722 57647 27774
rect 57383 27504 57435 27556
rect 57595 27504 57647 27556
rect 57383 27287 57435 27339
rect 57595 27287 57647 27339
rect 57383 27069 57435 27121
rect 57595 27069 57647 27121
rect 57383 26851 57435 26903
rect 57595 26851 57647 26903
rect 57383 26634 57435 26686
rect 57595 26634 57647 26686
rect 57383 26416 57435 26468
rect 57595 26416 57647 26468
rect 57383 26198 57435 26250
rect 57595 26198 57647 26250
rect 57383 25981 57435 26033
rect 57595 25981 57647 26033
rect 57383 25763 57435 25815
rect 57595 25763 57647 25815
rect 57383 25546 57435 25598
rect 57595 25546 57647 25598
rect 57383 25328 57435 25380
rect 57595 25328 57647 25380
rect 57383 25110 57435 25162
rect 57595 25110 57647 25162
rect 57383 24893 57435 24945
rect 57595 24893 57647 24945
rect 57383 24675 57435 24727
rect 57595 24675 57647 24727
rect 57383 24457 57435 24509
rect 57595 24457 57647 24509
rect 57383 24240 57435 24292
rect 57595 24240 57647 24292
rect 57383 24022 57435 24074
rect 57595 24022 57647 24074
rect 57383 23805 57435 23857
rect 57595 23805 57647 23857
rect 57383 23587 57435 23639
rect 57595 23587 57647 23639
rect 57383 23369 57435 23421
rect 57595 23369 57647 23421
rect 57383 23152 57435 23204
rect 57595 23152 57647 23204
rect 57383 22934 57435 22986
rect 57595 22934 57647 22986
rect 57383 22716 57435 22768
rect 57595 22716 57647 22768
rect 57383 22499 57435 22551
rect 57595 22499 57647 22551
rect 57383 22281 57435 22333
rect 57595 22281 57647 22333
rect 57383 22063 57435 22115
rect 57595 22063 57647 22115
rect 57383 21846 57435 21898
rect 57595 21846 57647 21898
rect 57383 21628 57435 21680
rect 57595 21628 57647 21680
rect 57383 21411 57435 21463
rect 57595 21411 57647 21463
rect 57383 21193 57435 21245
rect 57595 21193 57647 21245
rect 57383 20975 57435 21027
rect 57595 20975 57647 21027
rect 57383 20758 57435 20810
rect 57595 20758 57647 20810
rect 57383 20540 57435 20592
rect 57595 20540 57647 20592
rect 57383 20322 57435 20374
rect 57595 20322 57647 20374
rect 57383 20105 57435 20157
rect 57595 20105 57647 20157
rect 57383 19887 57435 19939
rect 57595 19887 57647 19939
rect 57383 19670 57435 19722
rect 57595 19670 57647 19722
rect 57383 19452 57435 19504
rect 57595 19452 57647 19504
rect 57383 19234 57435 19286
rect 57595 19234 57647 19286
rect 57383 19016 57435 19068
rect 57595 19016 57647 19068
rect 57383 18799 57435 18851
rect 57595 18799 57647 18851
rect 57383 18581 57435 18633
rect 57595 18581 57647 18633
rect 57383 18364 57435 18416
rect 57595 18364 57647 18416
rect 57383 18146 57435 18198
rect 57595 18146 57647 18198
rect 57383 17928 57435 17980
rect 57595 17928 57647 17980
rect 57383 17711 57435 17763
rect 57595 17711 57647 17763
rect 57383 17493 57435 17545
rect 57595 17493 57647 17545
rect 57383 17275 57435 17327
rect 57595 17275 57647 17327
rect 57383 17058 57435 17110
rect 57595 17058 57647 17110
rect 57383 16840 57435 16892
rect 57595 16840 57647 16892
rect 57383 16623 57435 16675
rect 57595 16623 57647 16675
rect 57383 16405 57435 16457
rect 57595 16405 57647 16457
rect 57383 16187 57435 16239
rect 57595 16187 57647 16239
rect 57383 15970 57435 16022
rect 57595 15970 57647 16022
rect 57383 15752 57435 15804
rect 57595 15752 57647 15804
rect 57383 15534 57435 15586
rect 57595 15534 57647 15586
rect 57383 15317 57435 15369
rect 57595 15317 57647 15369
rect 57383 15099 57435 15151
rect 57595 15099 57647 15151
rect 57383 14881 57435 14933
rect 57595 14881 57647 14933
rect 57383 14664 57435 14716
rect 57595 14664 57647 14716
rect 57383 14446 57435 14498
rect 57595 14446 57647 14498
rect 57383 14229 57435 14281
rect 57595 14229 57647 14281
rect 57383 14011 57435 14063
rect 57595 14011 57647 14063
rect 57383 13793 57435 13845
rect 57595 13793 57647 13845
rect 57383 13576 57435 13628
rect 57595 13576 57647 13628
rect 57383 13358 57435 13410
rect 57595 13358 57647 13410
rect 57383 13140 57435 13192
rect 57595 13140 57647 13192
rect 57383 12923 57435 12975
rect 57595 12923 57647 12975
rect 57383 12705 57435 12757
rect 57595 12705 57647 12757
rect 57383 12488 57435 12540
rect 57595 12488 57647 12540
rect 57383 12270 57435 12322
rect 57595 12270 57647 12322
rect 57383 12052 57435 12104
rect 57595 12052 57647 12104
rect 57383 11835 57435 11887
rect 57595 11835 57647 11887
rect 57383 11617 57435 11669
rect 57595 11617 57647 11669
rect 57383 11399 57435 11451
rect 57595 11399 57647 11451
rect 57383 11182 57435 11234
rect 57595 11182 57647 11234
rect 57383 10964 57435 11016
rect 57595 10964 57647 11016
rect 57383 10746 57435 10798
rect 57595 10746 57647 10798
rect 57383 10529 57435 10581
rect 57595 10529 57647 10581
rect 57383 10311 57435 10363
rect 57595 10311 57647 10363
rect 57383 10094 57435 10146
rect 57595 10094 57647 10146
rect 57383 9876 57435 9928
rect 57595 9876 57647 9928
rect 57383 9658 57435 9710
rect 57595 9658 57647 9710
rect 57383 9441 57435 9493
rect 57595 9441 57647 9493
rect 57383 9223 57435 9275
rect 57595 9223 57647 9275
rect 57383 9005 57435 9057
rect 57595 9005 57647 9057
rect 57383 8788 57435 8840
rect 57595 8788 57647 8840
rect 57383 8570 57435 8622
rect 57595 8570 57647 8622
rect 57383 8352 57435 8404
rect 57595 8352 57647 8404
rect 57383 8135 57435 8187
rect 57595 8135 57647 8187
rect 57383 7917 57435 7969
rect 57595 7917 57647 7969
rect 57383 7700 57435 7752
rect 57595 7700 57647 7752
rect 57383 7482 57435 7534
rect 57595 7482 57647 7534
rect 57383 7264 57435 7316
rect 57595 7264 57647 7316
rect 57383 7047 57435 7099
rect 57595 7047 57647 7099
rect 57383 6829 57435 6881
rect 57595 6829 57647 6881
rect 57383 6611 57435 6663
rect 57595 6611 57647 6663
rect 57383 6394 57435 6446
rect 57595 6394 57647 6446
rect 49908 6297 50064 6349
rect 27476 6176 27528 6228
rect 27688 6176 27740 6228
rect 27476 5959 27528 6011
rect 27688 5959 27740 6011
rect 27476 5741 27528 5793
rect 27688 5741 27740 5793
rect 27476 5523 27528 5575
rect 27688 5523 27740 5575
rect 27476 5306 27528 5358
rect 27688 5306 27740 5358
rect 57383 6176 57435 6228
rect 57595 6176 57647 6228
rect 57383 5959 57435 6011
rect 57595 5959 57647 6011
rect 57383 5741 57435 5793
rect 57595 5741 57647 5793
rect 57383 5523 57435 5575
rect 57595 5523 57647 5575
rect 57383 5306 57435 5358
rect 57595 5306 57647 5358
rect 51654 5147 51810 5199
rect 27476 4535 27528 4587
rect 27688 4535 27740 4587
rect 27476 4318 27528 4370
rect 27688 4318 27740 4370
rect 27476 4100 27528 4152
rect 27688 4100 27740 4152
rect 27476 3882 27528 3934
rect 27688 3882 27740 3934
rect 57383 4535 57435 4587
rect 57595 4535 57647 4587
rect 57383 4318 57435 4370
rect 57595 4318 57647 4370
rect 57383 4100 57435 4152
rect 57595 4100 57647 4152
rect 27476 3665 27528 3717
rect 27688 3665 27740 3717
rect 40623 3230 40779 3282
rect 57383 3882 57435 3934
rect 57595 3882 57647 3934
rect 57383 3665 57435 3717
rect 57595 3665 57647 3717
rect 57998 33380 58050 33432
rect 58210 33380 58262 33432
rect 57998 33163 58050 33215
rect 58210 33163 58262 33215
rect 57998 32945 58050 32997
rect 58210 32945 58262 32997
rect 57998 32727 58050 32779
rect 58210 32727 58262 32779
rect 57998 32510 58050 32562
rect 58210 32510 58262 32562
rect 57998 32292 58050 32344
rect 58210 32292 58262 32344
rect 57998 32075 58050 32127
rect 58210 32075 58262 32127
rect 57998 31857 58050 31909
rect 58210 31857 58262 31909
rect 57998 31639 58050 31691
rect 58210 31639 58262 31691
rect 57998 31422 58050 31474
rect 58210 31422 58262 31474
rect 57998 31204 58050 31256
rect 58210 31204 58262 31256
rect 57998 30986 58050 31038
rect 58210 30986 58262 31038
rect 57998 30769 58050 30821
rect 58210 30769 58262 30821
rect 57998 30551 58050 30603
rect 58210 30551 58262 30603
rect 57998 30334 58050 30386
rect 58210 30334 58262 30386
rect 57998 30116 58050 30168
rect 58210 30116 58262 30168
rect 57998 29898 58050 29950
rect 58210 29898 58262 29950
rect 57998 29681 58050 29733
rect 58210 29681 58262 29733
rect 57998 29463 58050 29515
rect 58210 29463 58262 29515
rect 57998 29245 58050 29297
rect 58210 29245 58262 29297
rect 57998 29028 58050 29080
rect 58210 29028 58262 29080
rect 57998 28810 58050 28862
rect 58210 28810 58262 28862
rect 57998 28592 58050 28644
rect 58210 28592 58262 28644
rect 57998 28375 58050 28427
rect 58210 28375 58262 28427
rect 57998 28157 58050 28209
rect 58210 28157 58262 28209
rect 57998 27940 58050 27992
rect 58210 27940 58262 27992
rect 57998 27722 58050 27774
rect 58210 27722 58262 27774
rect 57998 27504 58050 27556
rect 58210 27504 58262 27556
rect 57998 27287 58050 27339
rect 58210 27287 58262 27339
rect 57998 27069 58050 27121
rect 58210 27069 58262 27121
rect 57998 26851 58050 26903
rect 58210 26851 58262 26903
rect 57998 26634 58050 26686
rect 58210 26634 58262 26686
rect 57998 26416 58050 26468
rect 58210 26416 58262 26468
rect 57998 26198 58050 26250
rect 58210 26198 58262 26250
rect 57998 25981 58050 26033
rect 58210 25981 58262 26033
rect 57998 25763 58050 25815
rect 58210 25763 58262 25815
rect 57998 25546 58050 25598
rect 58210 25546 58262 25598
rect 57998 25328 58050 25380
rect 58210 25328 58262 25380
rect 57998 25110 58050 25162
rect 58210 25110 58262 25162
rect 57998 24893 58050 24945
rect 58210 24893 58262 24945
rect 57998 24675 58050 24727
rect 58210 24675 58262 24727
rect 57998 24457 58050 24509
rect 58210 24457 58262 24509
rect 57998 24240 58050 24292
rect 58210 24240 58262 24292
rect 57998 24022 58050 24074
rect 58210 24022 58262 24074
rect 57998 23805 58050 23857
rect 58210 23805 58262 23857
rect 57998 23587 58050 23639
rect 58210 23587 58262 23639
rect 57998 23369 58050 23421
rect 58210 23369 58262 23421
rect 57998 23152 58050 23204
rect 58210 23152 58262 23204
rect 57998 22934 58050 22986
rect 58210 22934 58262 22986
rect 57998 22716 58050 22768
rect 58210 22716 58262 22768
rect 57998 22499 58050 22551
rect 58210 22499 58262 22551
rect 57998 22281 58050 22333
rect 58210 22281 58262 22333
rect 57998 22063 58050 22115
rect 58210 22063 58262 22115
rect 57998 21846 58050 21898
rect 58210 21846 58262 21898
rect 57998 21628 58050 21680
rect 58210 21628 58262 21680
rect 57998 21411 58050 21463
rect 58210 21411 58262 21463
rect 57998 21193 58050 21245
rect 58210 21193 58262 21245
rect 57998 20975 58050 21027
rect 58210 20975 58262 21027
rect 57998 20758 58050 20810
rect 58210 20758 58262 20810
rect 57998 20540 58050 20592
rect 58210 20540 58262 20592
rect 57998 20322 58050 20374
rect 58210 20322 58262 20374
rect 57998 20105 58050 20157
rect 58210 20105 58262 20157
rect 57998 19887 58050 19939
rect 58210 19887 58262 19939
rect 57998 19670 58050 19722
rect 58210 19670 58262 19722
rect 57998 19452 58050 19504
rect 58210 19452 58262 19504
rect 57998 19234 58050 19286
rect 58210 19234 58262 19286
rect 57998 19016 58050 19068
rect 58210 19016 58262 19068
rect 57998 18799 58050 18851
rect 58210 18799 58262 18851
rect 57998 18581 58050 18633
rect 58210 18581 58262 18633
rect 57998 18364 58050 18416
rect 58210 18364 58262 18416
rect 57998 18146 58050 18198
rect 58210 18146 58262 18198
rect 57998 17928 58050 17980
rect 58210 17928 58262 17980
rect 57998 17711 58050 17763
rect 58210 17711 58262 17763
rect 57998 17493 58050 17545
rect 58210 17493 58262 17545
rect 57998 17275 58050 17327
rect 58210 17275 58262 17327
rect 57998 17058 58050 17110
rect 58210 17058 58262 17110
rect 57998 16840 58050 16892
rect 58210 16840 58262 16892
rect 57998 16623 58050 16675
rect 58210 16623 58262 16675
rect 57998 16405 58050 16457
rect 58210 16405 58262 16457
rect 57998 16187 58050 16239
rect 58210 16187 58262 16239
rect 57998 15970 58050 16022
rect 58210 15970 58262 16022
rect 57998 15752 58050 15804
rect 58210 15752 58262 15804
rect 57998 15534 58050 15586
rect 58210 15534 58262 15586
rect 57998 15317 58050 15369
rect 58210 15317 58262 15369
rect 57998 15099 58050 15151
rect 58210 15099 58262 15151
rect 57998 14881 58050 14933
rect 58210 14881 58262 14933
rect 57998 14664 58050 14716
rect 58210 14664 58262 14716
rect 57998 14446 58050 14498
rect 58210 14446 58262 14498
rect 57998 14229 58050 14281
rect 58210 14229 58262 14281
rect 57998 14011 58050 14063
rect 58210 14011 58262 14063
rect 57998 13793 58050 13845
rect 58210 13793 58262 13845
rect 57998 13576 58050 13628
rect 58210 13576 58262 13628
rect 57998 13358 58050 13410
rect 58210 13358 58262 13410
rect 57998 13140 58050 13192
rect 58210 13140 58262 13192
rect 57998 12923 58050 12975
rect 58210 12923 58262 12975
rect 57998 12705 58050 12757
rect 58210 12705 58262 12757
rect 57998 12488 58050 12540
rect 58210 12488 58262 12540
rect 57998 12270 58050 12322
rect 58210 12270 58262 12322
rect 57998 12052 58050 12104
rect 58210 12052 58262 12104
rect 57998 11835 58050 11887
rect 58210 11835 58262 11887
rect 57998 11617 58050 11669
rect 58210 11617 58262 11669
rect 57998 11399 58050 11451
rect 58210 11399 58262 11451
rect 57998 11182 58050 11234
rect 58210 11182 58262 11234
rect 57998 10964 58050 11016
rect 58210 10964 58262 11016
rect 57998 10746 58050 10798
rect 58210 10746 58262 10798
rect 57998 10529 58050 10581
rect 58210 10529 58262 10581
rect 57998 10311 58050 10363
rect 58210 10311 58262 10363
rect 57998 10094 58050 10146
rect 58210 10094 58262 10146
rect 57998 9876 58050 9928
rect 58210 9876 58262 9928
rect 57998 9658 58050 9710
rect 58210 9658 58262 9710
rect 57998 9441 58050 9493
rect 58210 9441 58262 9493
rect 57998 9223 58050 9275
rect 58210 9223 58262 9275
rect 57998 9005 58050 9057
rect 58210 9005 58262 9057
rect 57998 8788 58050 8840
rect 58210 8788 58262 8840
rect 57998 8570 58050 8622
rect 58210 8570 58262 8622
rect 57998 8352 58050 8404
rect 58210 8352 58262 8404
rect 57998 8135 58050 8187
rect 58210 8135 58262 8187
rect 57998 7917 58050 7969
rect 58210 7917 58262 7969
rect 57998 7700 58050 7752
rect 58210 7700 58262 7752
rect 57998 7482 58050 7534
rect 58210 7482 58262 7534
rect 57998 7264 58050 7316
rect 58210 7264 58262 7316
rect 57998 7047 58050 7099
rect 58210 7047 58262 7099
rect 57998 6829 58050 6881
rect 58210 6829 58262 6881
rect 57998 6611 58050 6663
rect 58210 6611 58262 6663
rect 57998 6394 58050 6446
rect 58210 6394 58262 6446
rect 57998 6176 58050 6228
rect 58210 6176 58262 6228
rect 57998 5959 58050 6011
rect 58210 5959 58262 6011
rect 57998 5741 58050 5793
rect 58210 5741 58262 5793
rect 57998 5523 58050 5575
rect 58210 5523 58262 5575
rect 57998 5306 58050 5358
rect 58210 5306 58262 5358
rect 61289 5323 61445 5479
rect 57998 4535 58050 4587
rect 58210 4535 58262 4587
rect 57998 4318 58050 4370
rect 58210 4318 58262 4370
rect 57998 4100 58050 4152
rect 58210 4100 58262 4152
rect 57998 3882 58050 3934
rect 58210 3882 58262 3934
rect 57998 3665 58050 3717
rect 58210 3665 58262 3717
rect 2574 1637 2730 1689
rect 12639 1637 12795 1689
rect 13089 1637 13245 1689
rect 23439 1637 23595 1689
rect 62149 1637 62305 1689
rect 72215 1637 72371 1689
rect 72665 1637 72821 1689
rect 82730 1637 82886 1689
rect 29092 657 29144 917
<< metal2 >>
rect 282 67568 86090 67894
rect 706 66376 86090 67376
rect 25313 65916 26039 65976
rect 25313 65860 25378 65916
rect 25434 65860 25502 65916
rect 25558 65860 25626 65916
rect 25682 65860 25750 65916
rect 25806 65860 25874 65916
rect 25930 65860 26039 65916
rect 25313 65792 26039 65860
rect 25313 65736 25378 65792
rect 25434 65736 25502 65792
rect 25558 65736 25626 65792
rect 25682 65736 25750 65792
rect 25806 65736 25874 65792
rect 25930 65736 26039 65792
rect 25313 34961 26039 65736
rect 25313 34905 25344 34961
rect 25400 34905 25468 34961
rect 25524 34905 25592 34961
rect 25648 34905 25716 34961
rect 25772 34905 25840 34961
rect 25896 34905 25964 34961
rect 26020 34905 26039 34961
rect 25313 34837 26039 34905
rect 25313 34781 25344 34837
rect 25400 34781 25468 34837
rect 25524 34781 25592 34837
rect 25648 34781 25716 34837
rect 25772 34781 25840 34837
rect 25896 34781 25964 34837
rect 26020 34781 26039 34837
rect 25313 34713 26039 34781
rect 25313 34657 25344 34713
rect 25400 34657 25468 34713
rect 25524 34657 25592 34713
rect 25648 34657 25716 34713
rect 25772 34657 25840 34713
rect 25896 34657 25964 34713
rect 26020 34657 26039 34713
rect 25313 31248 26039 34657
rect 25313 31192 25398 31248
rect 25454 31192 25522 31248
rect 25578 31192 25646 31248
rect 25702 31192 25770 31248
rect 25826 31192 25894 31248
rect 25950 31192 26039 31248
rect 25313 31124 26039 31192
rect 25313 31068 25398 31124
rect 25454 31068 25522 31124
rect 25578 31068 25646 31124
rect 25702 31068 25770 31124
rect 25826 31068 25894 31124
rect 25950 31068 26039 31124
rect 25313 31000 26039 31068
rect 25313 30944 25398 31000
rect 25454 30944 25522 31000
rect 25578 30944 25646 31000
rect 25702 30944 25770 31000
rect 25826 30944 25894 31000
rect 25950 30944 26039 31000
rect 25313 30793 26039 30944
rect 25313 30737 25398 30793
rect 25454 30737 25522 30793
rect 25578 30737 25646 30793
rect 25702 30737 25770 30793
rect 25826 30737 25894 30793
rect 25950 30737 26039 30793
rect 25313 30669 26039 30737
rect 25313 30613 25398 30669
rect 25454 30613 25522 30669
rect 25578 30613 25646 30669
rect 25702 30613 25770 30669
rect 25826 30613 25894 30669
rect 25950 30613 26039 30669
rect 25313 30545 26039 30613
rect 25313 30489 25398 30545
rect 25454 30489 25522 30545
rect 25578 30489 25646 30545
rect 25702 30489 25770 30545
rect 25826 30489 25894 30545
rect 25950 30489 26039 30545
rect 25313 28315 26039 30489
rect 25313 28259 25404 28315
rect 25460 28259 25528 28315
rect 25584 28259 25652 28315
rect 25708 28259 25776 28315
rect 25832 28259 25900 28315
rect 25956 28259 26039 28315
rect 25313 28191 26039 28259
rect 25313 28135 25404 28191
rect 25460 28135 25528 28191
rect 25584 28135 25652 28191
rect 25708 28135 25776 28191
rect 25832 28135 25900 28191
rect 25956 28135 26039 28191
rect 25313 28067 26039 28135
rect 25313 28011 25404 28067
rect 25460 28011 25528 28067
rect 25584 28011 25652 28067
rect 25708 28011 25776 28067
rect 25832 28011 25900 28067
rect 25956 28011 26039 28067
rect 25313 27943 26039 28011
rect 25313 27887 25404 27943
rect 25460 27887 25528 27943
rect 25584 27887 25652 27943
rect 25708 27887 25776 27943
rect 25832 27887 25900 27943
rect 25956 27887 26039 27943
rect 25313 27819 26039 27887
rect 25313 27763 25404 27819
rect 25460 27763 25528 27819
rect 25584 27763 25652 27819
rect 25708 27763 25776 27819
rect 25832 27763 25900 27819
rect 25956 27763 26039 27819
rect 25313 27695 26039 27763
rect 25313 27639 25404 27695
rect 25460 27639 25528 27695
rect 25584 27639 25652 27695
rect 25708 27639 25776 27695
rect 25832 27639 25900 27695
rect 25956 27639 26039 27695
rect 25313 27571 26039 27639
rect 25313 27515 25404 27571
rect 25460 27515 25528 27571
rect 25584 27515 25652 27571
rect 25708 27515 25776 27571
rect 25832 27515 25900 27571
rect 25956 27515 26039 27571
rect 25313 27447 26039 27515
rect 25313 27391 25404 27447
rect 25460 27391 25528 27447
rect 25584 27391 25652 27447
rect 25708 27391 25776 27447
rect 25832 27391 25900 27447
rect 25956 27391 26039 27447
rect 25313 27323 26039 27391
rect 26772 34011 27214 66376
rect 29486 65928 30364 66376
rect 26772 33955 26859 34011
rect 26915 33955 27071 34011
rect 27127 33955 27214 34011
rect 26772 33793 27214 33955
rect 26772 33737 26859 33793
rect 26915 33737 27071 33793
rect 27127 33737 27214 33793
rect 26772 33576 27214 33737
rect 26772 33520 26859 33576
rect 26915 33520 27071 33576
rect 27127 33520 27214 33576
rect 26772 33432 27214 33520
rect 26772 33380 26861 33432
rect 26913 33380 27073 33432
rect 27125 33380 27214 33432
rect 26772 33358 27214 33380
rect 26772 33302 26859 33358
rect 26915 33302 27071 33358
rect 27127 33302 27214 33358
rect 26772 33215 27214 33302
rect 26772 33163 26861 33215
rect 26913 33163 27073 33215
rect 27125 33163 27214 33215
rect 26772 33140 27214 33163
rect 26772 33084 26859 33140
rect 26915 33084 27071 33140
rect 27127 33084 27214 33140
rect 26772 32997 27214 33084
rect 26772 32945 26861 32997
rect 26913 32945 27073 32997
rect 27125 32945 27214 32997
rect 26772 32922 27214 32945
rect 26772 32866 26859 32922
rect 26915 32866 27071 32922
rect 27127 32866 27214 32922
rect 26772 32779 27214 32866
rect 26772 32727 26861 32779
rect 26913 32727 27073 32779
rect 27125 32727 27214 32779
rect 26772 32705 27214 32727
rect 26772 32649 26859 32705
rect 26915 32649 27071 32705
rect 27127 32649 27214 32705
rect 26772 32562 27214 32649
rect 26772 32510 26861 32562
rect 26913 32510 27073 32562
rect 27125 32510 27214 32562
rect 26772 32487 27214 32510
rect 26772 32431 26859 32487
rect 26915 32431 27071 32487
rect 27127 32431 27214 32487
rect 26772 32344 27214 32431
rect 26772 32292 26861 32344
rect 26913 32292 27073 32344
rect 27125 32292 27214 32344
rect 26772 32127 27214 32292
rect 26772 32088 26861 32127
rect 26913 32088 27073 32127
rect 27125 32088 27214 32127
rect 26772 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 27214 32088
rect 26772 31909 27214 32032
rect 26772 31870 26861 31909
rect 26913 31870 27073 31909
rect 27125 31870 27214 31909
rect 26772 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 27214 31870
rect 26772 31691 27214 31814
rect 26772 31652 26861 31691
rect 26913 31652 27073 31691
rect 27125 31652 27214 31691
rect 26772 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 27214 31652
rect 26772 31474 27214 31596
rect 26772 31422 26861 31474
rect 26913 31422 27073 31474
rect 27125 31422 27214 31474
rect 26772 31256 27214 31422
rect 26772 31204 26861 31256
rect 26913 31204 27073 31256
rect 27125 31204 27214 31256
rect 26772 31038 27214 31204
rect 26772 30986 26861 31038
rect 26913 30986 27073 31038
rect 27125 30986 27214 31038
rect 26772 30821 27214 30986
rect 26772 30769 26861 30821
rect 26913 30769 27073 30821
rect 27125 30769 27214 30821
rect 26772 30603 27214 30769
rect 26772 30551 26861 30603
rect 26913 30551 27073 30603
rect 27125 30551 27214 30603
rect 26772 30386 27214 30551
rect 26772 30334 26861 30386
rect 26913 30334 27073 30386
rect 27125 30334 27214 30386
rect 26772 30168 27214 30334
rect 26772 30116 26861 30168
rect 26913 30116 27073 30168
rect 27125 30116 27214 30168
rect 26772 29968 27214 30116
rect 26772 29912 26859 29968
rect 26915 29912 27071 29968
rect 27127 29912 27214 29968
rect 26772 29898 26861 29912
rect 26913 29898 27073 29912
rect 27125 29898 27214 29912
rect 26772 29750 27214 29898
rect 26772 29694 26859 29750
rect 26915 29694 27071 29750
rect 27127 29694 27214 29750
rect 26772 29681 26861 29694
rect 26913 29681 27073 29694
rect 27125 29681 27214 29694
rect 26772 29533 27214 29681
rect 26772 29477 26859 29533
rect 26915 29477 27071 29533
rect 27127 29477 27214 29533
rect 26772 29463 26861 29477
rect 26913 29463 27073 29477
rect 27125 29463 27214 29477
rect 26772 29315 27214 29463
rect 26772 29259 26859 29315
rect 26915 29259 27071 29315
rect 27127 29259 27214 29315
rect 26772 29245 26861 29259
rect 26913 29245 27073 29259
rect 27125 29245 27214 29259
rect 26772 29098 27214 29245
rect 26772 29042 26859 29098
rect 26915 29042 27071 29098
rect 27127 29042 27214 29098
rect 26772 29028 26861 29042
rect 26913 29028 27073 29042
rect 27125 29028 27214 29042
rect 26772 28880 27214 29028
rect 26772 28824 26859 28880
rect 26915 28824 27071 28880
rect 27127 28824 27214 28880
rect 26772 28810 26861 28824
rect 26913 28810 27073 28824
rect 27125 28810 27214 28824
rect 26772 28662 27214 28810
rect 26772 28606 26859 28662
rect 26915 28606 27071 28662
rect 27127 28606 27214 28662
rect 26772 28592 26861 28606
rect 26913 28592 27073 28606
rect 27125 28592 27214 28606
rect 26772 28444 27214 28592
rect 26772 28388 26859 28444
rect 26915 28388 27071 28444
rect 27127 28388 27214 28444
rect 26772 28375 26861 28388
rect 26913 28375 27073 28388
rect 27125 28375 27214 28388
rect 26772 28227 27214 28375
rect 26772 28171 26859 28227
rect 26915 28171 27071 28227
rect 27127 28171 27214 28227
rect 26772 28157 26861 28171
rect 26913 28157 27073 28171
rect 27125 28157 27214 28171
rect 26772 28009 27214 28157
rect 26772 27953 26859 28009
rect 26915 27953 27071 28009
rect 27127 27953 27214 28009
rect 26772 27940 26861 27953
rect 26913 27940 27073 27953
rect 27125 27940 27214 27953
rect 26772 27792 27214 27940
rect 26772 27736 26859 27792
rect 26915 27736 27071 27792
rect 27127 27736 27214 27792
rect 26772 27722 26861 27736
rect 26913 27722 27073 27736
rect 27125 27722 27214 27736
rect 26772 27574 27214 27722
rect 26772 27518 26859 27574
rect 26915 27518 27071 27574
rect 27127 27518 27214 27574
rect 26772 27504 26861 27518
rect 26913 27504 27073 27518
rect 27125 27504 27214 27518
rect 26772 27382 27214 27504
rect 27387 65855 29146 65894
rect 27387 65799 27788 65855
rect 27844 65799 27999 65855
rect 28055 65799 28210 65855
rect 28266 65799 28421 65855
rect 28477 65799 28632 65855
rect 28688 65799 28843 65855
rect 28899 65799 29054 65855
rect 29110 65799 29146 65855
rect 27387 65760 29146 65799
rect 29485 65853 30365 65928
rect 29485 65801 29582 65853
rect 29634 65801 29793 65853
rect 29845 65801 30005 65853
rect 30057 65801 30216 65853
rect 30268 65801 30365 65853
rect 27387 64094 27828 65760
rect 29485 64955 30365 65801
rect 29485 64899 29580 64955
rect 29636 64899 29791 64955
rect 29847 64899 30003 64955
rect 30059 64899 30214 64955
rect 30270 64899 30365 64955
rect 30769 65853 32888 66376
rect 30769 65801 30807 65853
rect 30859 65801 31018 65853
rect 31070 65801 31229 65853
rect 31281 65801 31440 65853
rect 31492 65801 31651 65853
rect 31703 65801 31861 65853
rect 31913 65801 32072 65853
rect 32124 65801 32283 65853
rect 32335 65801 32494 65853
rect 32546 65801 32888 65853
rect 30769 65635 32888 65801
rect 30769 65583 30807 65635
rect 30859 65583 31018 65635
rect 31070 65583 31229 65635
rect 31281 65583 31440 65635
rect 31492 65583 31651 65635
rect 31703 65583 31861 65635
rect 31913 65583 32072 65635
rect 32124 65583 32283 65635
rect 32335 65583 32494 65635
rect 32546 65583 32888 65635
rect 30769 65418 32888 65583
rect 30769 65366 30807 65418
rect 30859 65366 31018 65418
rect 31070 65366 31229 65418
rect 31281 65366 31440 65418
rect 31492 65366 31651 65418
rect 31703 65366 31861 65418
rect 31913 65366 32072 65418
rect 32124 65366 32283 65418
rect 32335 65366 32494 65418
rect 32546 65366 32888 65418
rect 34227 65855 35024 65928
rect 34227 65799 34288 65855
rect 34344 65799 34499 65855
rect 34555 65799 34710 65855
rect 34766 65799 34921 65855
rect 34977 65799 35024 65855
rect 34227 65635 35024 65799
rect 34227 65583 34290 65635
rect 34342 65583 34501 65635
rect 34553 65583 34712 65635
rect 34764 65583 34923 65635
rect 34975 65583 35024 65635
rect 30769 65078 32888 65366
rect 33011 65374 33984 65413
rect 33011 65318 33048 65374
rect 33104 65318 33259 65374
rect 33315 65318 33470 65374
rect 33526 65318 33681 65374
rect 33737 65318 33892 65374
rect 33948 65318 33984 65374
rect 33011 65280 33984 65318
rect 34227 65078 35024 65583
rect 35128 65833 36415 66376
rect 35128 65781 35443 65833
rect 35495 65781 35654 65833
rect 35706 65781 35865 65833
rect 35917 65781 36076 65833
rect 36128 65781 36287 65833
rect 36339 65781 36415 65833
rect 35128 65370 36415 65781
rect 35128 65318 35443 65370
rect 35495 65318 35654 65370
rect 35706 65318 35865 65370
rect 35917 65318 36076 65370
rect 36128 65318 36287 65370
rect 36339 65318 36415 65370
rect 30769 64955 32889 65078
rect 30769 64940 30852 64955
rect 27387 64055 29146 64094
rect 27387 63999 27788 64055
rect 27844 63999 27999 64055
rect 28055 63999 28210 64055
rect 28266 63999 28421 64055
rect 28477 63999 28632 64055
rect 28688 63999 28843 64055
rect 28899 63999 29054 64055
rect 29110 63999 29146 64055
rect 27387 63960 29146 63999
rect 29485 64053 30365 64899
rect 29485 64001 29582 64053
rect 29634 64001 29793 64053
rect 29845 64001 30005 64053
rect 30057 64001 30216 64053
rect 30268 64001 30365 64053
rect 27387 62294 27828 63960
rect 29485 63155 30365 64001
rect 29485 63099 29580 63155
rect 29636 63099 29791 63155
rect 29847 63099 30003 63155
rect 30059 63099 30214 63155
rect 30270 63099 30365 63155
rect 27387 62255 29146 62294
rect 27387 62199 27788 62255
rect 27844 62199 27999 62255
rect 28055 62199 28210 62255
rect 28266 62199 28421 62255
rect 28477 62199 28632 62255
rect 28688 62199 28843 62255
rect 28899 62199 29054 62255
rect 29110 62199 29146 62255
rect 27387 62160 29146 62199
rect 29485 62253 30365 63099
rect 29485 62201 29582 62253
rect 29634 62201 29793 62253
rect 29845 62201 30005 62253
rect 30057 62201 30216 62253
rect 30268 62201 30365 62253
rect 27387 60494 27828 62160
rect 29485 61355 30365 62201
rect 29485 61299 29580 61355
rect 29636 61299 29791 61355
rect 29847 61299 30003 61355
rect 30059 61299 30214 61355
rect 30270 61299 30365 61355
rect 27387 60455 29146 60494
rect 27387 60399 27788 60455
rect 27844 60399 27999 60455
rect 28055 60399 28210 60455
rect 28266 60399 28421 60455
rect 28477 60399 28632 60455
rect 28688 60399 28843 60455
rect 28899 60399 29054 60455
rect 29110 60399 29146 60455
rect 27387 60360 29146 60399
rect 29485 60453 30365 61299
rect 29485 60401 29582 60453
rect 29634 60401 29793 60453
rect 29845 60401 30005 60453
rect 30057 60401 30216 60453
rect 30268 60401 30365 60453
rect 27387 58694 27828 60360
rect 29485 59555 30365 60401
rect 29485 59499 29580 59555
rect 29636 59499 29791 59555
rect 29847 59499 30003 59555
rect 30059 59499 30214 59555
rect 30270 59499 30365 59555
rect 27387 58655 29146 58694
rect 27387 58599 27788 58655
rect 27844 58599 27999 58655
rect 28055 58599 28210 58655
rect 28266 58599 28421 58655
rect 28477 58599 28632 58655
rect 28688 58599 28843 58655
rect 28899 58599 29054 58655
rect 29110 58599 29146 58655
rect 27387 58560 29146 58599
rect 29485 58653 30365 59499
rect 29485 58601 29582 58653
rect 29634 58601 29793 58653
rect 29845 58601 30005 58653
rect 30057 58601 30216 58653
rect 30268 58601 30365 58653
rect 27387 56894 27828 58560
rect 29485 57755 30365 58601
rect 29485 57699 29580 57755
rect 29636 57699 29791 57755
rect 29847 57699 30003 57755
rect 30059 57699 30214 57755
rect 30270 57699 30365 57755
rect 27387 56855 29146 56894
rect 27387 56799 27788 56855
rect 27844 56799 27999 56855
rect 28055 56799 28210 56855
rect 28266 56799 28421 56855
rect 28477 56799 28632 56855
rect 28688 56799 28843 56855
rect 28899 56799 29054 56855
rect 29110 56799 29146 56855
rect 27387 56760 29146 56799
rect 29485 56853 30365 57699
rect 29485 56801 29582 56853
rect 29634 56801 29793 56853
rect 29845 56801 30005 56853
rect 30057 56801 30216 56853
rect 30268 56801 30365 56853
rect 27387 55094 27828 56760
rect 29485 55955 30365 56801
rect 29485 55899 29580 55955
rect 29636 55899 29791 55955
rect 29847 55899 30003 55955
rect 30059 55899 30214 55955
rect 30270 55899 30365 55955
rect 27387 55055 29146 55094
rect 27387 54999 27788 55055
rect 27844 54999 27999 55055
rect 28055 54999 28210 55055
rect 28266 54999 28421 55055
rect 28477 54999 28632 55055
rect 28688 54999 28843 55055
rect 28899 54999 29054 55055
rect 29110 54999 29146 55055
rect 27387 54960 29146 54999
rect 29485 55053 30365 55899
rect 29485 55001 29582 55053
rect 29634 55001 29793 55053
rect 29845 55001 30005 55053
rect 30057 55001 30216 55053
rect 30268 55001 30365 55053
rect 27387 53294 27828 54960
rect 29485 54155 30365 55001
rect 29485 54099 29580 54155
rect 29636 54099 29791 54155
rect 29847 54099 30003 54155
rect 30059 54099 30214 54155
rect 30270 54099 30365 54155
rect 27387 53255 29146 53294
rect 27387 53199 27788 53255
rect 27844 53199 27999 53255
rect 28055 53199 28210 53255
rect 28266 53199 28421 53255
rect 28477 53199 28632 53255
rect 28688 53199 28843 53255
rect 28899 53199 29054 53255
rect 29110 53199 29146 53255
rect 27387 53160 29146 53199
rect 29485 53253 30365 54099
rect 29485 53201 29582 53253
rect 29634 53201 29793 53253
rect 29845 53201 30005 53253
rect 30057 53201 30216 53253
rect 30268 53201 30365 53253
rect 27387 51494 27828 53160
rect 29485 52355 30365 53201
rect 29485 52299 29580 52355
rect 29636 52299 29791 52355
rect 29847 52299 30003 52355
rect 30059 52299 30214 52355
rect 30270 52299 30365 52355
rect 27387 51455 29146 51494
rect 27387 51399 27788 51455
rect 27844 51399 27999 51455
rect 28055 51399 28210 51455
rect 28266 51399 28421 51455
rect 28477 51399 28632 51455
rect 28688 51399 28843 51455
rect 28899 51399 29054 51455
rect 29110 51399 29146 51455
rect 27387 51360 29146 51399
rect 29485 51453 30365 52299
rect 29485 51401 29582 51453
rect 29634 51401 29793 51453
rect 29845 51401 30005 51453
rect 30057 51401 30216 51453
rect 30268 51401 30365 51453
rect 27387 49694 27828 51360
rect 29485 50555 30365 51401
rect 29485 50499 29580 50555
rect 29636 50499 29791 50555
rect 29847 50499 30003 50555
rect 30059 50499 30214 50555
rect 30270 50499 30365 50555
rect 27387 49655 29146 49694
rect 27387 49599 27788 49655
rect 27844 49599 27999 49655
rect 28055 49599 28210 49655
rect 28266 49599 28421 49655
rect 28477 49599 28632 49655
rect 28688 49599 28843 49655
rect 28899 49599 29054 49655
rect 29110 49599 29146 49655
rect 27387 49560 29146 49599
rect 29485 49653 30365 50499
rect 29485 49601 29582 49653
rect 29634 49601 29793 49653
rect 29845 49601 30005 49653
rect 30057 49601 30216 49653
rect 30268 49601 30365 49653
rect 27387 47894 27828 49560
rect 29485 48755 30365 49601
rect 29485 48699 29580 48755
rect 29636 48699 29791 48755
rect 29847 48699 30003 48755
rect 30059 48699 30214 48755
rect 30270 48699 30365 48755
rect 27387 47855 29146 47894
rect 27387 47799 27788 47855
rect 27844 47799 27999 47855
rect 28055 47799 28210 47855
rect 28266 47799 28421 47855
rect 28477 47799 28632 47855
rect 28688 47799 28843 47855
rect 28899 47799 29054 47855
rect 29110 47799 29146 47855
rect 27387 47760 29146 47799
rect 29485 47853 30365 48699
rect 29485 47801 29582 47853
rect 29634 47801 29793 47853
rect 29845 47801 30005 47853
rect 30057 47801 30216 47853
rect 30268 47801 30365 47853
rect 27387 46094 27828 47760
rect 29485 46955 30365 47801
rect 29485 46899 29580 46955
rect 29636 46899 29791 46955
rect 29847 46899 30003 46955
rect 30059 46899 30214 46955
rect 30270 46899 30365 46955
rect 27387 46055 29146 46094
rect 27387 45999 27788 46055
rect 27844 45999 27999 46055
rect 28055 45999 28210 46055
rect 28266 45999 28421 46055
rect 28477 45999 28632 46055
rect 28688 45999 28843 46055
rect 28899 45999 29054 46055
rect 29110 45999 29146 46055
rect 27387 45960 29146 45999
rect 29485 46053 30365 46899
rect 29485 46001 29582 46053
rect 29634 46001 29793 46053
rect 29845 46001 30005 46053
rect 30057 46001 30216 46053
rect 30268 46001 30365 46053
rect 27387 44294 27828 45960
rect 29485 45155 30365 46001
rect 29485 45099 29580 45155
rect 29636 45099 29791 45155
rect 29847 45099 30003 45155
rect 30059 45099 30214 45155
rect 30270 45099 30365 45155
rect 27387 44255 29146 44294
rect 27387 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 29146 44255
rect 27387 44160 29146 44199
rect 29485 44253 30365 45099
rect 29485 44201 29582 44253
rect 29634 44201 29793 44253
rect 29845 44201 30005 44253
rect 30057 44201 30216 44253
rect 30268 44201 30365 44253
rect 27387 42494 27828 44160
rect 29485 43355 30365 44201
rect 29485 43299 29580 43355
rect 29636 43299 29791 43355
rect 29847 43299 30003 43355
rect 30059 43299 30214 43355
rect 30270 43299 30365 43355
rect 27387 42455 29146 42494
rect 27387 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 29146 42455
rect 27387 42360 29146 42399
rect 29485 42453 30365 43299
rect 29485 42401 29582 42453
rect 29634 42401 29793 42453
rect 29845 42401 30005 42453
rect 30057 42401 30216 42453
rect 30268 42401 30365 42453
rect 27387 40694 27828 42360
rect 29485 41555 30365 42401
rect 29485 41499 29580 41555
rect 29636 41499 29791 41555
rect 29847 41499 30003 41555
rect 30059 41499 30214 41555
rect 30270 41499 30365 41555
rect 27387 40655 29146 40694
rect 27387 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 29146 40655
rect 27387 40560 29146 40599
rect 29485 40653 30365 41499
rect 29485 40601 29582 40653
rect 29634 40601 29793 40653
rect 29845 40601 30005 40653
rect 30057 40601 30216 40653
rect 30268 40601 30365 40653
rect 27387 38894 27828 40560
rect 29485 39755 30365 40601
rect 29485 39699 29580 39755
rect 29636 39699 29791 39755
rect 29847 39699 30003 39755
rect 30059 39699 30214 39755
rect 30270 39699 30365 39755
rect 27387 38855 29146 38894
rect 27387 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 29146 38855
rect 27387 38760 29146 38799
rect 29485 38853 30365 39699
rect 29485 38801 29582 38853
rect 29634 38801 29793 38853
rect 29845 38801 30005 38853
rect 30057 38801 30216 38853
rect 30268 38801 30365 38853
rect 27387 37094 27828 38760
rect 29485 37955 30365 38801
rect 29485 37899 29580 37955
rect 29636 37899 29791 37955
rect 29847 37899 30003 37955
rect 30059 37899 30214 37955
rect 30270 37899 30365 37955
rect 27387 37055 29146 37094
rect 27387 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 29146 37055
rect 27387 36960 29146 36999
rect 29485 37053 30365 37899
rect 29485 37001 29582 37053
rect 29634 37001 29793 37053
rect 29845 37001 30005 37053
rect 30057 37001 30216 37053
rect 30268 37001 30365 37053
rect 27387 35024 27828 36960
rect 29485 36155 30365 37001
rect 29485 36099 29580 36155
rect 29636 36099 29791 36155
rect 29847 36099 30003 36155
rect 30059 36099 30214 36155
rect 30270 36099 30365 36155
rect 29485 36027 30365 36099
rect 30770 64899 30852 64940
rect 30908 64899 31063 64955
rect 31119 64899 31274 64955
rect 31330 64899 31484 64955
rect 31540 64899 31695 64955
rect 31751 64899 31907 64955
rect 31963 64899 32118 64955
rect 32174 64899 32328 64955
rect 32384 64899 32539 64955
rect 32595 64899 32750 64955
rect 32806 64899 32889 64955
rect 34227 64953 35025 65078
rect 34227 64940 34284 64953
rect 30770 64053 32889 64899
rect 34228 64901 34284 64940
rect 34336 64901 34495 64953
rect 34547 64901 34707 64953
rect 34759 64901 34918 64953
rect 34970 64901 35025 64953
rect 35128 64955 36415 65318
rect 35128 64940 35218 64955
rect 33019 64729 33327 64770
rect 33019 64677 33057 64729
rect 33109 64677 33237 64729
rect 33289 64677 33327 64729
rect 33019 64522 33327 64677
rect 33019 64466 33055 64522
rect 33111 64466 33235 64522
rect 33291 64466 33327 64522
rect 33019 64281 33327 64466
rect 33731 64737 34090 64778
rect 33731 64685 33819 64737
rect 33871 64685 33999 64737
rect 34051 64685 34090 64737
rect 33731 64515 34090 64685
rect 33731 64459 33817 64515
rect 33873 64459 33997 64515
rect 34053 64459 34090 64515
rect 33731 64386 34090 64459
rect 34228 64491 35025 64901
rect 34228 64439 34267 64491
rect 34319 64439 34447 64491
rect 34499 64439 34627 64491
rect 34679 64439 35025 64491
rect 33019 64229 33057 64281
rect 33109 64229 33237 64281
rect 33289 64229 33327 64281
rect 33019 64189 33327 64229
rect 30770 64001 30854 64053
rect 30906 64001 31065 64053
rect 31117 64001 31276 64053
rect 31328 64001 31486 64053
rect 31538 64001 31697 64053
rect 31749 64001 31909 64053
rect 31961 64001 32120 64053
rect 32172 64001 32330 64053
rect 32382 64001 32541 64053
rect 32593 64001 32752 64053
rect 32804 64001 32889 64053
rect 30770 63155 32889 64001
rect 34228 64055 35025 64439
rect 34228 63999 34282 64055
rect 34338 63999 34493 64055
rect 34549 63999 34705 64055
rect 34761 64053 34916 64055
rect 34972 64053 35025 64055
rect 34807 64001 34916 64053
rect 34987 64001 35025 64053
rect 34761 63999 34916 64001
rect 34972 63999 35025 64001
rect 33019 63825 33327 63865
rect 33019 63773 33057 63825
rect 33109 63773 33237 63825
rect 33289 63773 33327 63825
rect 33019 63588 33327 63773
rect 33019 63532 33055 63588
rect 33111 63532 33235 63588
rect 33291 63532 33327 63588
rect 33019 63377 33327 63532
rect 33019 63325 33057 63377
rect 33109 63325 33237 63377
rect 33289 63325 33327 63377
rect 33019 63284 33327 63325
rect 33731 63595 34090 63668
rect 33731 63539 33817 63595
rect 33873 63539 33997 63595
rect 34053 63539 34090 63595
rect 33731 63369 34090 63539
rect 33731 63317 33819 63369
rect 33871 63317 33999 63369
rect 34051 63317 34090 63369
rect 33731 63276 34090 63317
rect 34228 63615 35025 63999
rect 34228 63563 34267 63615
rect 34319 63563 34447 63615
rect 34499 63563 34627 63615
rect 34679 63563 35025 63615
rect 30770 63099 30852 63155
rect 30908 63099 31063 63155
rect 31119 63099 31274 63155
rect 31330 63099 31484 63155
rect 31540 63099 31695 63155
rect 31751 63099 31907 63155
rect 31963 63099 32118 63155
rect 32174 63099 32328 63155
rect 32384 63099 32539 63155
rect 32595 63099 32750 63155
rect 32806 63099 32889 63155
rect 30770 62253 32889 63099
rect 34228 63153 35025 63563
rect 34228 63101 34284 63153
rect 34336 63101 34495 63153
rect 34547 63101 34707 63153
rect 34759 63101 34918 63153
rect 34970 63101 35025 63153
rect 33019 62929 33327 62970
rect 33019 62877 33057 62929
rect 33109 62877 33237 62929
rect 33289 62877 33327 62929
rect 33019 62722 33327 62877
rect 33019 62666 33055 62722
rect 33111 62666 33235 62722
rect 33291 62666 33327 62722
rect 33019 62481 33327 62666
rect 33731 62937 34090 62978
rect 33731 62885 33819 62937
rect 33871 62885 33999 62937
rect 34051 62885 34090 62937
rect 33731 62715 34090 62885
rect 33731 62659 33817 62715
rect 33873 62659 33997 62715
rect 34053 62659 34090 62715
rect 33731 62586 34090 62659
rect 34228 62691 35025 63101
rect 34228 62639 34267 62691
rect 34319 62639 34447 62691
rect 34499 62639 34627 62691
rect 34679 62639 35025 62691
rect 33019 62429 33057 62481
rect 33109 62429 33237 62481
rect 33289 62429 33327 62481
rect 33019 62389 33327 62429
rect 30770 62201 30854 62253
rect 30906 62201 31065 62253
rect 31117 62201 31276 62253
rect 31328 62201 31486 62253
rect 31538 62201 31697 62253
rect 31749 62201 31909 62253
rect 31961 62201 32120 62253
rect 32172 62201 32330 62253
rect 32382 62201 32541 62253
rect 32593 62201 32752 62253
rect 32804 62201 32889 62253
rect 30770 61355 32889 62201
rect 34228 62255 35025 62639
rect 34228 62199 34282 62255
rect 34338 62199 34493 62255
rect 34549 62199 34705 62255
rect 34761 62253 34916 62255
rect 34972 62253 35025 62255
rect 34807 62201 34916 62253
rect 34987 62201 35025 62253
rect 34761 62199 34916 62201
rect 34972 62199 35025 62201
rect 33019 62025 33327 62065
rect 33019 61973 33057 62025
rect 33109 61973 33237 62025
rect 33289 61973 33327 62025
rect 33019 61788 33327 61973
rect 33019 61732 33055 61788
rect 33111 61732 33235 61788
rect 33291 61732 33327 61788
rect 33019 61577 33327 61732
rect 33019 61525 33057 61577
rect 33109 61525 33237 61577
rect 33289 61525 33327 61577
rect 33019 61484 33327 61525
rect 33731 61795 34090 61868
rect 33731 61739 33817 61795
rect 33873 61739 33997 61795
rect 34053 61739 34090 61795
rect 33731 61569 34090 61739
rect 33731 61517 33819 61569
rect 33871 61517 33999 61569
rect 34051 61517 34090 61569
rect 33731 61476 34090 61517
rect 34228 61815 35025 62199
rect 34228 61763 34267 61815
rect 34319 61763 34447 61815
rect 34499 61763 34627 61815
rect 34679 61763 35025 61815
rect 30770 61299 30852 61355
rect 30908 61299 31063 61355
rect 31119 61299 31274 61355
rect 31330 61299 31484 61355
rect 31540 61299 31695 61355
rect 31751 61299 31907 61355
rect 31963 61299 32118 61355
rect 32174 61299 32328 61355
rect 32384 61299 32539 61355
rect 32595 61299 32750 61355
rect 32806 61299 32889 61355
rect 30770 60453 32889 61299
rect 34228 61353 35025 61763
rect 34228 61301 34284 61353
rect 34336 61301 34495 61353
rect 34547 61301 34707 61353
rect 34759 61301 34918 61353
rect 34970 61301 35025 61353
rect 33019 61129 33327 61170
rect 33019 61077 33057 61129
rect 33109 61077 33237 61129
rect 33289 61077 33327 61129
rect 33019 60922 33327 61077
rect 33019 60866 33055 60922
rect 33111 60866 33235 60922
rect 33291 60866 33327 60922
rect 33019 60681 33327 60866
rect 33731 61137 34090 61178
rect 33731 61085 33819 61137
rect 33871 61085 33999 61137
rect 34051 61085 34090 61137
rect 33731 60915 34090 61085
rect 33731 60859 33817 60915
rect 33873 60859 33997 60915
rect 34053 60859 34090 60915
rect 33731 60786 34090 60859
rect 34228 60891 35025 61301
rect 34228 60839 34267 60891
rect 34319 60839 34447 60891
rect 34499 60839 34627 60891
rect 34679 60839 35025 60891
rect 33019 60629 33057 60681
rect 33109 60629 33237 60681
rect 33289 60629 33327 60681
rect 33019 60589 33327 60629
rect 30770 60401 30854 60453
rect 30906 60401 31065 60453
rect 31117 60401 31276 60453
rect 31328 60401 31486 60453
rect 31538 60401 31697 60453
rect 31749 60401 31909 60453
rect 31961 60401 32120 60453
rect 32172 60401 32330 60453
rect 32382 60401 32541 60453
rect 32593 60401 32752 60453
rect 32804 60401 32889 60453
rect 30770 59555 32889 60401
rect 34228 60455 35025 60839
rect 34228 60399 34282 60455
rect 34338 60399 34493 60455
rect 34549 60399 34705 60455
rect 34761 60453 34916 60455
rect 34972 60453 35025 60455
rect 34807 60401 34916 60453
rect 34987 60401 35025 60453
rect 34761 60399 34916 60401
rect 34972 60399 35025 60401
rect 33019 60225 33327 60265
rect 33019 60173 33057 60225
rect 33109 60173 33237 60225
rect 33289 60173 33327 60225
rect 33019 59988 33327 60173
rect 33019 59932 33055 59988
rect 33111 59932 33235 59988
rect 33291 59932 33327 59988
rect 33019 59777 33327 59932
rect 33019 59725 33057 59777
rect 33109 59725 33237 59777
rect 33289 59725 33327 59777
rect 33019 59684 33327 59725
rect 33731 59995 34090 60068
rect 33731 59939 33817 59995
rect 33873 59939 33997 59995
rect 34053 59939 34090 59995
rect 33731 59769 34090 59939
rect 33731 59717 33819 59769
rect 33871 59717 33999 59769
rect 34051 59717 34090 59769
rect 33731 59676 34090 59717
rect 34228 60015 35025 60399
rect 34228 59963 34267 60015
rect 34319 59963 34447 60015
rect 34499 59963 34627 60015
rect 34679 59963 35025 60015
rect 30770 59499 30852 59555
rect 30908 59499 31063 59555
rect 31119 59499 31274 59555
rect 31330 59499 31484 59555
rect 31540 59499 31695 59555
rect 31751 59499 31907 59555
rect 31963 59499 32118 59555
rect 32174 59499 32328 59555
rect 32384 59499 32539 59555
rect 32595 59499 32750 59555
rect 32806 59499 32889 59555
rect 30770 58653 32889 59499
rect 34228 59553 35025 59963
rect 34228 59501 34284 59553
rect 34336 59501 34495 59553
rect 34547 59501 34707 59553
rect 34759 59501 34918 59553
rect 34970 59501 35025 59553
rect 33019 59329 33327 59370
rect 33019 59277 33057 59329
rect 33109 59277 33237 59329
rect 33289 59277 33327 59329
rect 33019 59122 33327 59277
rect 33019 59066 33055 59122
rect 33111 59066 33235 59122
rect 33291 59066 33327 59122
rect 33019 58881 33327 59066
rect 33731 59337 34090 59378
rect 33731 59285 33819 59337
rect 33871 59285 33999 59337
rect 34051 59285 34090 59337
rect 33731 59115 34090 59285
rect 33731 59059 33817 59115
rect 33873 59059 33997 59115
rect 34053 59059 34090 59115
rect 33731 58986 34090 59059
rect 34228 59091 35025 59501
rect 34228 59039 34267 59091
rect 34319 59039 34447 59091
rect 34499 59039 34627 59091
rect 34679 59039 35025 59091
rect 33019 58829 33057 58881
rect 33109 58829 33237 58881
rect 33289 58829 33327 58881
rect 33019 58789 33327 58829
rect 30770 58601 30854 58653
rect 30906 58601 31065 58653
rect 31117 58601 31276 58653
rect 31328 58601 31486 58653
rect 31538 58601 31697 58653
rect 31749 58601 31909 58653
rect 31961 58601 32120 58653
rect 32172 58601 32330 58653
rect 32382 58601 32541 58653
rect 32593 58601 32752 58653
rect 32804 58601 32889 58653
rect 30770 57755 32889 58601
rect 34228 58655 35025 59039
rect 34228 58599 34282 58655
rect 34338 58599 34493 58655
rect 34549 58599 34705 58655
rect 34761 58653 34916 58655
rect 34972 58653 35025 58655
rect 34807 58601 34916 58653
rect 34987 58601 35025 58653
rect 34761 58599 34916 58601
rect 34972 58599 35025 58601
rect 33019 58425 33327 58465
rect 33019 58373 33057 58425
rect 33109 58373 33237 58425
rect 33289 58373 33327 58425
rect 33019 58188 33327 58373
rect 33019 58132 33055 58188
rect 33111 58132 33235 58188
rect 33291 58132 33327 58188
rect 33019 57977 33327 58132
rect 33019 57925 33057 57977
rect 33109 57925 33237 57977
rect 33289 57925 33327 57977
rect 33019 57884 33327 57925
rect 33731 58195 34090 58268
rect 33731 58139 33817 58195
rect 33873 58139 33997 58195
rect 34053 58139 34090 58195
rect 33731 57969 34090 58139
rect 33731 57917 33819 57969
rect 33871 57917 33999 57969
rect 34051 57917 34090 57969
rect 33731 57876 34090 57917
rect 34228 58215 35025 58599
rect 34228 58163 34267 58215
rect 34319 58163 34447 58215
rect 34499 58163 34627 58215
rect 34679 58163 35025 58215
rect 30770 57699 30852 57755
rect 30908 57699 31063 57755
rect 31119 57699 31274 57755
rect 31330 57699 31484 57755
rect 31540 57699 31695 57755
rect 31751 57699 31907 57755
rect 31963 57699 32118 57755
rect 32174 57699 32328 57755
rect 32384 57699 32539 57755
rect 32595 57699 32750 57755
rect 32806 57699 32889 57755
rect 30770 56853 32889 57699
rect 34228 57753 35025 58163
rect 34228 57701 34284 57753
rect 34336 57701 34495 57753
rect 34547 57701 34707 57753
rect 34759 57701 34918 57753
rect 34970 57701 35025 57753
rect 33019 57529 33327 57570
rect 33019 57477 33057 57529
rect 33109 57477 33237 57529
rect 33289 57477 33327 57529
rect 33019 57322 33327 57477
rect 33019 57266 33055 57322
rect 33111 57266 33235 57322
rect 33291 57266 33327 57322
rect 33019 57081 33327 57266
rect 33731 57537 34090 57578
rect 33731 57485 33819 57537
rect 33871 57485 33999 57537
rect 34051 57485 34090 57537
rect 33731 57315 34090 57485
rect 33731 57259 33817 57315
rect 33873 57259 33997 57315
rect 34053 57259 34090 57315
rect 33731 57186 34090 57259
rect 34228 57291 35025 57701
rect 34228 57239 34267 57291
rect 34319 57239 34447 57291
rect 34499 57239 34627 57291
rect 34679 57239 35025 57291
rect 33019 57029 33057 57081
rect 33109 57029 33237 57081
rect 33289 57029 33327 57081
rect 33019 56989 33327 57029
rect 30770 56801 30854 56853
rect 30906 56801 31065 56853
rect 31117 56801 31276 56853
rect 31328 56801 31486 56853
rect 31538 56801 31697 56853
rect 31749 56801 31909 56853
rect 31961 56801 32120 56853
rect 32172 56801 32330 56853
rect 32382 56801 32541 56853
rect 32593 56801 32752 56853
rect 32804 56801 32889 56853
rect 30770 55955 32889 56801
rect 34228 56855 35025 57239
rect 34228 56799 34282 56855
rect 34338 56799 34493 56855
rect 34549 56799 34705 56855
rect 34761 56853 34916 56855
rect 34972 56853 35025 56855
rect 34807 56801 34916 56853
rect 34987 56801 35025 56853
rect 34761 56799 34916 56801
rect 34972 56799 35025 56801
rect 33019 56625 33327 56665
rect 33019 56573 33057 56625
rect 33109 56573 33237 56625
rect 33289 56573 33327 56625
rect 33019 56388 33327 56573
rect 33019 56332 33055 56388
rect 33111 56332 33235 56388
rect 33291 56332 33327 56388
rect 33019 56177 33327 56332
rect 33019 56125 33057 56177
rect 33109 56125 33237 56177
rect 33289 56125 33327 56177
rect 33019 56084 33327 56125
rect 33731 56395 34090 56468
rect 33731 56339 33817 56395
rect 33873 56339 33997 56395
rect 34053 56339 34090 56395
rect 33731 56169 34090 56339
rect 33731 56117 33819 56169
rect 33871 56117 33999 56169
rect 34051 56117 34090 56169
rect 33731 56076 34090 56117
rect 34228 56415 35025 56799
rect 34228 56363 34267 56415
rect 34319 56363 34447 56415
rect 34499 56363 34627 56415
rect 34679 56363 35025 56415
rect 30770 55899 30852 55955
rect 30908 55899 31063 55955
rect 31119 55899 31274 55955
rect 31330 55899 31484 55955
rect 31540 55899 31695 55955
rect 31751 55899 31907 55955
rect 31963 55899 32118 55955
rect 32174 55899 32328 55955
rect 32384 55899 32539 55955
rect 32595 55899 32750 55955
rect 32806 55899 32889 55955
rect 30770 55053 32889 55899
rect 34228 55953 35025 56363
rect 34228 55901 34284 55953
rect 34336 55901 34495 55953
rect 34547 55901 34707 55953
rect 34759 55901 34918 55953
rect 34970 55901 35025 55953
rect 33019 55729 33327 55770
rect 33019 55677 33057 55729
rect 33109 55677 33237 55729
rect 33289 55677 33327 55729
rect 33019 55522 33327 55677
rect 33019 55466 33055 55522
rect 33111 55466 33235 55522
rect 33291 55466 33327 55522
rect 33019 55281 33327 55466
rect 33731 55737 34090 55778
rect 33731 55685 33819 55737
rect 33871 55685 33999 55737
rect 34051 55685 34090 55737
rect 33731 55515 34090 55685
rect 33731 55459 33817 55515
rect 33873 55459 33997 55515
rect 34053 55459 34090 55515
rect 33731 55386 34090 55459
rect 34228 55491 35025 55901
rect 34228 55439 34267 55491
rect 34319 55439 34447 55491
rect 34499 55439 34627 55491
rect 34679 55439 35025 55491
rect 33019 55229 33057 55281
rect 33109 55229 33237 55281
rect 33289 55229 33327 55281
rect 33019 55189 33327 55229
rect 30770 55001 30854 55053
rect 30906 55001 31065 55053
rect 31117 55001 31276 55053
rect 31328 55001 31486 55053
rect 31538 55001 31697 55053
rect 31749 55001 31909 55053
rect 31961 55001 32120 55053
rect 32172 55001 32330 55053
rect 32382 55001 32541 55053
rect 32593 55001 32752 55053
rect 32804 55001 32889 55053
rect 30770 54155 32889 55001
rect 34228 55055 35025 55439
rect 34228 54999 34282 55055
rect 34338 54999 34493 55055
rect 34549 54999 34705 55055
rect 34761 55053 34916 55055
rect 34972 55053 35025 55055
rect 34807 55001 34916 55053
rect 34987 55001 35025 55053
rect 34761 54999 34916 55001
rect 34972 54999 35025 55001
rect 33019 54825 33327 54865
rect 33019 54773 33057 54825
rect 33109 54773 33237 54825
rect 33289 54773 33327 54825
rect 33019 54588 33327 54773
rect 33019 54532 33055 54588
rect 33111 54532 33235 54588
rect 33291 54532 33327 54588
rect 33019 54377 33327 54532
rect 33019 54325 33057 54377
rect 33109 54325 33237 54377
rect 33289 54325 33327 54377
rect 33019 54284 33327 54325
rect 33731 54595 34090 54668
rect 33731 54539 33817 54595
rect 33873 54539 33997 54595
rect 34053 54539 34090 54595
rect 33731 54369 34090 54539
rect 33731 54317 33819 54369
rect 33871 54317 33999 54369
rect 34051 54317 34090 54369
rect 33731 54276 34090 54317
rect 34228 54615 35025 54999
rect 34228 54563 34267 54615
rect 34319 54563 34447 54615
rect 34499 54563 34627 54615
rect 34679 54563 35025 54615
rect 30770 54099 30852 54155
rect 30908 54099 31063 54155
rect 31119 54099 31274 54155
rect 31330 54099 31484 54155
rect 31540 54099 31695 54155
rect 31751 54099 31907 54155
rect 31963 54099 32118 54155
rect 32174 54099 32328 54155
rect 32384 54099 32539 54155
rect 32595 54099 32750 54155
rect 32806 54099 32889 54155
rect 30770 53253 32889 54099
rect 34228 54153 35025 54563
rect 34228 54101 34284 54153
rect 34336 54101 34495 54153
rect 34547 54101 34707 54153
rect 34759 54101 34918 54153
rect 34970 54101 35025 54153
rect 33019 53929 33327 53970
rect 33019 53877 33057 53929
rect 33109 53877 33237 53929
rect 33289 53877 33327 53929
rect 33019 53722 33327 53877
rect 33019 53666 33055 53722
rect 33111 53666 33235 53722
rect 33291 53666 33327 53722
rect 33019 53481 33327 53666
rect 33731 53937 34090 53978
rect 33731 53885 33819 53937
rect 33871 53885 33999 53937
rect 34051 53885 34090 53937
rect 33731 53715 34090 53885
rect 33731 53659 33817 53715
rect 33873 53659 33997 53715
rect 34053 53659 34090 53715
rect 33731 53586 34090 53659
rect 34228 53691 35025 54101
rect 34228 53639 34267 53691
rect 34319 53639 34447 53691
rect 34499 53639 34627 53691
rect 34679 53639 35025 53691
rect 33019 53429 33057 53481
rect 33109 53429 33237 53481
rect 33289 53429 33327 53481
rect 33019 53389 33327 53429
rect 30770 53201 30854 53253
rect 30906 53201 31065 53253
rect 31117 53201 31276 53253
rect 31328 53201 31486 53253
rect 31538 53201 31697 53253
rect 31749 53201 31909 53253
rect 31961 53201 32120 53253
rect 32172 53201 32330 53253
rect 32382 53201 32541 53253
rect 32593 53201 32752 53253
rect 32804 53201 32889 53253
rect 30770 52355 32889 53201
rect 34228 53255 35025 53639
rect 34228 53199 34282 53255
rect 34338 53199 34493 53255
rect 34549 53199 34705 53255
rect 34761 53253 34916 53255
rect 34972 53253 35025 53255
rect 34807 53201 34916 53253
rect 34987 53201 35025 53253
rect 34761 53199 34916 53201
rect 34972 53199 35025 53201
rect 33019 53025 33327 53065
rect 33019 52973 33057 53025
rect 33109 52973 33237 53025
rect 33289 52973 33327 53025
rect 33019 52788 33327 52973
rect 33019 52732 33055 52788
rect 33111 52732 33235 52788
rect 33291 52732 33327 52788
rect 33019 52577 33327 52732
rect 33019 52525 33057 52577
rect 33109 52525 33237 52577
rect 33289 52525 33327 52577
rect 33019 52484 33327 52525
rect 33731 52795 34090 52868
rect 33731 52739 33817 52795
rect 33873 52739 33997 52795
rect 34053 52739 34090 52795
rect 33731 52569 34090 52739
rect 33731 52517 33819 52569
rect 33871 52517 33999 52569
rect 34051 52517 34090 52569
rect 33731 52476 34090 52517
rect 34228 52815 35025 53199
rect 34228 52763 34267 52815
rect 34319 52763 34447 52815
rect 34499 52763 34627 52815
rect 34679 52763 35025 52815
rect 30770 52299 30852 52355
rect 30908 52299 31063 52355
rect 31119 52299 31274 52355
rect 31330 52299 31484 52355
rect 31540 52299 31695 52355
rect 31751 52299 31907 52355
rect 31963 52299 32118 52355
rect 32174 52299 32328 52355
rect 32384 52299 32539 52355
rect 32595 52299 32750 52355
rect 32806 52299 32889 52355
rect 30770 51453 32889 52299
rect 34228 52353 35025 52763
rect 34228 52301 34284 52353
rect 34336 52301 34495 52353
rect 34547 52301 34707 52353
rect 34759 52301 34918 52353
rect 34970 52301 35025 52353
rect 33019 52129 33327 52170
rect 33019 52077 33057 52129
rect 33109 52077 33237 52129
rect 33289 52077 33327 52129
rect 33019 51922 33327 52077
rect 33019 51866 33055 51922
rect 33111 51866 33235 51922
rect 33291 51866 33327 51922
rect 33019 51681 33327 51866
rect 33731 52137 34090 52178
rect 33731 52085 33819 52137
rect 33871 52085 33999 52137
rect 34051 52085 34090 52137
rect 33731 51915 34090 52085
rect 33731 51859 33817 51915
rect 33873 51859 33997 51915
rect 34053 51859 34090 51915
rect 33731 51786 34090 51859
rect 34228 51891 35025 52301
rect 34228 51839 34267 51891
rect 34319 51839 34447 51891
rect 34499 51839 34627 51891
rect 34679 51839 35025 51891
rect 33019 51629 33057 51681
rect 33109 51629 33237 51681
rect 33289 51629 33327 51681
rect 33019 51589 33327 51629
rect 30770 51401 30854 51453
rect 30906 51401 31065 51453
rect 31117 51401 31276 51453
rect 31328 51401 31486 51453
rect 31538 51401 31697 51453
rect 31749 51401 31909 51453
rect 31961 51401 32120 51453
rect 32172 51401 32330 51453
rect 32382 51401 32541 51453
rect 32593 51401 32752 51453
rect 32804 51401 32889 51453
rect 30770 50555 32889 51401
rect 34228 51455 35025 51839
rect 34228 51399 34282 51455
rect 34338 51399 34493 51455
rect 34549 51399 34705 51455
rect 34761 51453 34916 51455
rect 34972 51453 35025 51455
rect 34807 51401 34916 51453
rect 34987 51401 35025 51453
rect 34761 51399 34916 51401
rect 34972 51399 35025 51401
rect 33019 51225 33327 51265
rect 33019 51173 33057 51225
rect 33109 51173 33237 51225
rect 33289 51173 33327 51225
rect 33019 50988 33327 51173
rect 33019 50932 33055 50988
rect 33111 50932 33235 50988
rect 33291 50932 33327 50988
rect 33019 50777 33327 50932
rect 33019 50725 33057 50777
rect 33109 50725 33237 50777
rect 33289 50725 33327 50777
rect 33019 50684 33327 50725
rect 33731 50995 34090 51068
rect 33731 50939 33817 50995
rect 33873 50939 33997 50995
rect 34053 50939 34090 50995
rect 33731 50769 34090 50939
rect 33731 50717 33819 50769
rect 33871 50717 33999 50769
rect 34051 50717 34090 50769
rect 33731 50676 34090 50717
rect 34228 51015 35025 51399
rect 34228 50963 34267 51015
rect 34319 50963 34447 51015
rect 34499 50963 34627 51015
rect 34679 50963 35025 51015
rect 30770 50499 30852 50555
rect 30908 50499 31063 50555
rect 31119 50499 31274 50555
rect 31330 50499 31484 50555
rect 31540 50499 31695 50555
rect 31751 50499 31907 50555
rect 31963 50499 32118 50555
rect 32174 50499 32328 50555
rect 32384 50499 32539 50555
rect 32595 50499 32750 50555
rect 32806 50499 32889 50555
rect 30770 49653 32889 50499
rect 34228 50553 35025 50963
rect 34228 50501 34284 50553
rect 34336 50501 34495 50553
rect 34547 50501 34707 50553
rect 34759 50501 34918 50553
rect 34970 50501 35025 50553
rect 33019 50329 33327 50370
rect 33019 50277 33057 50329
rect 33109 50277 33237 50329
rect 33289 50277 33327 50329
rect 33019 50122 33327 50277
rect 33019 50066 33055 50122
rect 33111 50066 33235 50122
rect 33291 50066 33327 50122
rect 33019 49881 33327 50066
rect 33731 50337 34090 50378
rect 33731 50285 33819 50337
rect 33871 50285 33999 50337
rect 34051 50285 34090 50337
rect 33731 50115 34090 50285
rect 33731 50059 33817 50115
rect 33873 50059 33997 50115
rect 34053 50059 34090 50115
rect 33731 49986 34090 50059
rect 34228 50091 35025 50501
rect 34228 50039 34267 50091
rect 34319 50039 34447 50091
rect 34499 50039 34627 50091
rect 34679 50039 35025 50091
rect 33019 49829 33057 49881
rect 33109 49829 33237 49881
rect 33289 49829 33327 49881
rect 33019 49789 33327 49829
rect 30770 49601 30854 49653
rect 30906 49601 31065 49653
rect 31117 49601 31276 49653
rect 31328 49601 31486 49653
rect 31538 49601 31697 49653
rect 31749 49601 31909 49653
rect 31961 49601 32120 49653
rect 32172 49601 32330 49653
rect 32382 49601 32541 49653
rect 32593 49601 32752 49653
rect 32804 49601 32889 49653
rect 30770 48755 32889 49601
rect 34228 49655 35025 50039
rect 34228 49599 34282 49655
rect 34338 49599 34493 49655
rect 34549 49599 34705 49655
rect 34761 49653 34916 49655
rect 34972 49653 35025 49655
rect 34807 49601 34916 49653
rect 34987 49601 35025 49653
rect 34761 49599 34916 49601
rect 34972 49599 35025 49601
rect 33019 49425 33327 49465
rect 33019 49373 33057 49425
rect 33109 49373 33237 49425
rect 33289 49373 33327 49425
rect 33019 49188 33327 49373
rect 33019 49132 33055 49188
rect 33111 49132 33235 49188
rect 33291 49132 33327 49188
rect 33019 48977 33327 49132
rect 33019 48925 33057 48977
rect 33109 48925 33237 48977
rect 33289 48925 33327 48977
rect 33019 48884 33327 48925
rect 33731 49195 34090 49268
rect 33731 49139 33817 49195
rect 33873 49139 33997 49195
rect 34053 49139 34090 49195
rect 33731 48969 34090 49139
rect 33731 48917 33819 48969
rect 33871 48917 33999 48969
rect 34051 48917 34090 48969
rect 33731 48876 34090 48917
rect 34228 49215 35025 49599
rect 34228 49163 34267 49215
rect 34319 49163 34447 49215
rect 34499 49163 34627 49215
rect 34679 49163 35025 49215
rect 30770 48699 30852 48755
rect 30908 48699 31063 48755
rect 31119 48699 31274 48755
rect 31330 48699 31484 48755
rect 31540 48699 31695 48755
rect 31751 48699 31907 48755
rect 31963 48699 32118 48755
rect 32174 48699 32328 48755
rect 32384 48699 32539 48755
rect 32595 48699 32750 48755
rect 32806 48699 32889 48755
rect 30770 47853 32889 48699
rect 34228 48753 35025 49163
rect 34228 48701 34284 48753
rect 34336 48701 34495 48753
rect 34547 48701 34707 48753
rect 34759 48701 34918 48753
rect 34970 48701 35025 48753
rect 33019 48529 33327 48570
rect 33019 48477 33057 48529
rect 33109 48477 33237 48529
rect 33289 48477 33327 48529
rect 33019 48322 33327 48477
rect 33019 48266 33055 48322
rect 33111 48266 33235 48322
rect 33291 48266 33327 48322
rect 33019 48081 33327 48266
rect 33731 48537 34090 48578
rect 33731 48485 33819 48537
rect 33871 48485 33999 48537
rect 34051 48485 34090 48537
rect 33731 48315 34090 48485
rect 33731 48259 33817 48315
rect 33873 48259 33997 48315
rect 34053 48259 34090 48315
rect 33731 48186 34090 48259
rect 34228 48291 35025 48701
rect 34228 48239 34267 48291
rect 34319 48239 34447 48291
rect 34499 48239 34627 48291
rect 34679 48239 35025 48291
rect 33019 48029 33057 48081
rect 33109 48029 33237 48081
rect 33289 48029 33327 48081
rect 33019 47989 33327 48029
rect 30770 47801 30854 47853
rect 30906 47801 31065 47853
rect 31117 47801 31276 47853
rect 31328 47801 31486 47853
rect 31538 47801 31697 47853
rect 31749 47801 31909 47853
rect 31961 47801 32120 47853
rect 32172 47801 32330 47853
rect 32382 47801 32541 47853
rect 32593 47801 32752 47853
rect 32804 47801 32889 47853
rect 30770 46955 32889 47801
rect 34228 47855 35025 48239
rect 34228 47799 34282 47855
rect 34338 47799 34493 47855
rect 34549 47799 34705 47855
rect 34761 47853 34916 47855
rect 34972 47853 35025 47855
rect 34807 47801 34916 47853
rect 34987 47801 35025 47853
rect 34761 47799 34916 47801
rect 34972 47799 35025 47801
rect 33019 47625 33327 47665
rect 33019 47573 33057 47625
rect 33109 47573 33237 47625
rect 33289 47573 33327 47625
rect 33019 47388 33327 47573
rect 33019 47332 33055 47388
rect 33111 47332 33235 47388
rect 33291 47332 33327 47388
rect 33019 47177 33327 47332
rect 33019 47125 33057 47177
rect 33109 47125 33237 47177
rect 33289 47125 33327 47177
rect 33019 47084 33327 47125
rect 33731 47395 34090 47468
rect 33731 47339 33817 47395
rect 33873 47339 33997 47395
rect 34053 47339 34090 47395
rect 33731 47169 34090 47339
rect 33731 47117 33819 47169
rect 33871 47117 33999 47169
rect 34051 47117 34090 47169
rect 33731 47076 34090 47117
rect 34228 47415 35025 47799
rect 34228 47363 34267 47415
rect 34319 47363 34447 47415
rect 34499 47363 34627 47415
rect 34679 47363 35025 47415
rect 30770 46899 30852 46955
rect 30908 46899 31063 46955
rect 31119 46899 31274 46955
rect 31330 46899 31484 46955
rect 31540 46899 31695 46955
rect 31751 46899 31907 46955
rect 31963 46899 32118 46955
rect 32174 46899 32328 46955
rect 32384 46899 32539 46955
rect 32595 46899 32750 46955
rect 32806 46899 32889 46955
rect 30770 46053 32889 46899
rect 34228 46953 35025 47363
rect 34228 46901 34284 46953
rect 34336 46901 34495 46953
rect 34547 46901 34707 46953
rect 34759 46901 34918 46953
rect 34970 46901 35025 46953
rect 33019 46729 33327 46770
rect 33019 46677 33057 46729
rect 33109 46677 33237 46729
rect 33289 46677 33327 46729
rect 33019 46522 33327 46677
rect 33019 46466 33055 46522
rect 33111 46466 33235 46522
rect 33291 46466 33327 46522
rect 33019 46281 33327 46466
rect 33731 46737 34090 46778
rect 33731 46685 33819 46737
rect 33871 46685 33999 46737
rect 34051 46685 34090 46737
rect 33731 46515 34090 46685
rect 33731 46459 33817 46515
rect 33873 46459 33997 46515
rect 34053 46459 34090 46515
rect 33731 46386 34090 46459
rect 34228 46491 35025 46901
rect 34228 46439 34267 46491
rect 34319 46439 34447 46491
rect 34499 46439 34627 46491
rect 34679 46439 35025 46491
rect 33019 46229 33057 46281
rect 33109 46229 33237 46281
rect 33289 46229 33327 46281
rect 33019 46189 33327 46229
rect 30770 46001 30854 46053
rect 30906 46001 31065 46053
rect 31117 46001 31276 46053
rect 31328 46001 31486 46053
rect 31538 46001 31697 46053
rect 31749 46001 31909 46053
rect 31961 46001 32120 46053
rect 32172 46001 32330 46053
rect 32382 46001 32541 46053
rect 32593 46001 32752 46053
rect 32804 46001 32889 46053
rect 30770 45155 32889 46001
rect 34228 46055 35025 46439
rect 34228 45999 34282 46055
rect 34338 45999 34493 46055
rect 34549 45999 34705 46055
rect 34761 46053 34916 46055
rect 34972 46053 35025 46055
rect 34807 46001 34916 46053
rect 34987 46001 35025 46053
rect 34761 45999 34916 46001
rect 34972 45999 35025 46001
rect 33019 45825 33327 45865
rect 33019 45773 33057 45825
rect 33109 45773 33237 45825
rect 33289 45773 33327 45825
rect 33019 45588 33327 45773
rect 33019 45532 33055 45588
rect 33111 45532 33235 45588
rect 33291 45532 33327 45588
rect 33019 45377 33327 45532
rect 33019 45325 33057 45377
rect 33109 45325 33237 45377
rect 33289 45325 33327 45377
rect 33019 45284 33327 45325
rect 33731 45595 34090 45668
rect 33731 45539 33817 45595
rect 33873 45539 33997 45595
rect 34053 45539 34090 45595
rect 33731 45369 34090 45539
rect 33731 45317 33819 45369
rect 33871 45317 33999 45369
rect 34051 45317 34090 45369
rect 33731 45276 34090 45317
rect 34228 45615 35025 45999
rect 34228 45563 34267 45615
rect 34319 45563 34447 45615
rect 34499 45563 34627 45615
rect 34679 45563 35025 45615
rect 30770 45099 30852 45155
rect 30908 45099 31063 45155
rect 31119 45099 31274 45155
rect 31330 45099 31484 45155
rect 31540 45099 31695 45155
rect 31751 45099 31907 45155
rect 31963 45099 32118 45155
rect 32174 45099 32328 45155
rect 32384 45099 32539 45155
rect 32595 45099 32750 45155
rect 32806 45099 32889 45155
rect 30770 44253 32889 45099
rect 34228 45153 35025 45563
rect 34228 45101 34284 45153
rect 34336 45101 34495 45153
rect 34547 45101 34707 45153
rect 34759 45101 34918 45153
rect 34970 45101 35025 45153
rect 33019 44929 33327 44970
rect 33019 44877 33057 44929
rect 33109 44877 33237 44929
rect 33289 44877 33327 44929
rect 33019 44722 33327 44877
rect 33019 44666 33055 44722
rect 33111 44666 33235 44722
rect 33291 44666 33327 44722
rect 33019 44481 33327 44666
rect 33731 44937 34090 44978
rect 33731 44885 33819 44937
rect 33871 44885 33999 44937
rect 34051 44885 34090 44937
rect 33731 44715 34090 44885
rect 33731 44659 33817 44715
rect 33873 44659 33997 44715
rect 34053 44659 34090 44715
rect 33731 44586 34090 44659
rect 34228 44691 35025 45101
rect 34228 44639 34267 44691
rect 34319 44639 34447 44691
rect 34499 44639 34627 44691
rect 34679 44639 35025 44691
rect 33019 44429 33057 44481
rect 33109 44429 33237 44481
rect 33289 44429 33327 44481
rect 33019 44389 33327 44429
rect 30770 44201 30854 44253
rect 30906 44201 31065 44253
rect 31117 44201 31276 44253
rect 31328 44201 31486 44253
rect 31538 44201 31697 44253
rect 31749 44201 31909 44253
rect 31961 44201 32120 44253
rect 32172 44201 32330 44253
rect 32382 44201 32541 44253
rect 32593 44201 32752 44253
rect 32804 44201 32889 44253
rect 30770 43355 32889 44201
rect 34228 44255 35025 44639
rect 34228 44199 34282 44255
rect 34338 44199 34493 44255
rect 34549 44199 34705 44255
rect 34761 44253 34916 44255
rect 34972 44253 35025 44255
rect 34807 44201 34916 44253
rect 34987 44201 35025 44253
rect 34761 44199 34916 44201
rect 34972 44199 35025 44201
rect 33019 44025 33327 44065
rect 33019 43973 33057 44025
rect 33109 43973 33237 44025
rect 33289 43973 33327 44025
rect 33019 43788 33327 43973
rect 33019 43732 33055 43788
rect 33111 43732 33235 43788
rect 33291 43732 33327 43788
rect 33019 43577 33327 43732
rect 33019 43525 33057 43577
rect 33109 43525 33237 43577
rect 33289 43525 33327 43577
rect 33019 43484 33327 43525
rect 33731 43795 34090 43868
rect 33731 43739 33817 43795
rect 33873 43739 33997 43795
rect 34053 43739 34090 43795
rect 33731 43569 34090 43739
rect 33731 43517 33819 43569
rect 33871 43517 33999 43569
rect 34051 43517 34090 43569
rect 33731 43476 34090 43517
rect 34228 43815 35025 44199
rect 34228 43763 34267 43815
rect 34319 43763 34447 43815
rect 34499 43763 34627 43815
rect 34679 43763 35025 43815
rect 30770 43299 30852 43355
rect 30908 43299 31063 43355
rect 31119 43299 31274 43355
rect 31330 43299 31484 43355
rect 31540 43299 31695 43355
rect 31751 43299 31907 43355
rect 31963 43299 32118 43355
rect 32174 43299 32328 43355
rect 32384 43299 32539 43355
rect 32595 43299 32750 43355
rect 32806 43299 32889 43355
rect 30770 42453 32889 43299
rect 34228 43353 35025 43763
rect 34228 43301 34284 43353
rect 34336 43301 34495 43353
rect 34547 43301 34707 43353
rect 34759 43301 34918 43353
rect 34970 43301 35025 43353
rect 33019 43129 33327 43170
rect 33019 43077 33057 43129
rect 33109 43077 33237 43129
rect 33289 43077 33327 43129
rect 33019 42922 33327 43077
rect 33019 42866 33055 42922
rect 33111 42866 33235 42922
rect 33291 42866 33327 42922
rect 33019 42681 33327 42866
rect 33731 43137 34090 43178
rect 33731 43085 33819 43137
rect 33871 43085 33999 43137
rect 34051 43085 34090 43137
rect 33731 42915 34090 43085
rect 33731 42859 33817 42915
rect 33873 42859 33997 42915
rect 34053 42859 34090 42915
rect 33731 42786 34090 42859
rect 34228 42891 35025 43301
rect 34228 42839 34267 42891
rect 34319 42839 34447 42891
rect 34499 42839 34627 42891
rect 34679 42839 35025 42891
rect 33019 42629 33057 42681
rect 33109 42629 33237 42681
rect 33289 42629 33327 42681
rect 33019 42589 33327 42629
rect 30770 42401 30854 42453
rect 30906 42401 31065 42453
rect 31117 42401 31276 42453
rect 31328 42401 31486 42453
rect 31538 42401 31697 42453
rect 31749 42401 31909 42453
rect 31961 42401 32120 42453
rect 32172 42401 32330 42453
rect 32382 42401 32541 42453
rect 32593 42401 32752 42453
rect 32804 42401 32889 42453
rect 30770 41555 32889 42401
rect 34228 42455 35025 42839
rect 34228 42399 34282 42455
rect 34338 42399 34493 42455
rect 34549 42399 34705 42455
rect 34761 42453 34916 42455
rect 34972 42453 35025 42455
rect 34807 42401 34916 42453
rect 34987 42401 35025 42453
rect 34761 42399 34916 42401
rect 34972 42399 35025 42401
rect 33019 42225 33327 42265
rect 33019 42173 33057 42225
rect 33109 42173 33237 42225
rect 33289 42173 33327 42225
rect 33019 41988 33327 42173
rect 33019 41932 33055 41988
rect 33111 41932 33235 41988
rect 33291 41932 33327 41988
rect 33019 41777 33327 41932
rect 33019 41725 33057 41777
rect 33109 41725 33237 41777
rect 33289 41725 33327 41777
rect 33019 41684 33327 41725
rect 33731 41995 34090 42068
rect 33731 41939 33817 41995
rect 33873 41939 33997 41995
rect 34053 41939 34090 41995
rect 33731 41769 34090 41939
rect 33731 41717 33819 41769
rect 33871 41717 33999 41769
rect 34051 41717 34090 41769
rect 33731 41676 34090 41717
rect 34228 42015 35025 42399
rect 34228 41963 34267 42015
rect 34319 41963 34447 42015
rect 34499 41963 34627 42015
rect 34679 41963 35025 42015
rect 30770 41499 30852 41555
rect 30908 41499 31063 41555
rect 31119 41499 31274 41555
rect 31330 41499 31484 41555
rect 31540 41499 31695 41555
rect 31751 41499 31907 41555
rect 31963 41499 32118 41555
rect 32174 41499 32328 41555
rect 32384 41499 32539 41555
rect 32595 41499 32750 41555
rect 32806 41499 32889 41555
rect 30770 40653 32889 41499
rect 34228 41553 35025 41963
rect 34228 41501 34284 41553
rect 34336 41501 34495 41553
rect 34547 41501 34707 41553
rect 34759 41501 34918 41553
rect 34970 41501 35025 41553
rect 33019 41329 33327 41370
rect 33019 41277 33057 41329
rect 33109 41277 33237 41329
rect 33289 41277 33327 41329
rect 33019 41122 33327 41277
rect 33019 41066 33055 41122
rect 33111 41066 33235 41122
rect 33291 41066 33327 41122
rect 33019 40881 33327 41066
rect 33731 41337 34090 41378
rect 33731 41285 33819 41337
rect 33871 41285 33999 41337
rect 34051 41285 34090 41337
rect 33731 41115 34090 41285
rect 33731 41059 33817 41115
rect 33873 41059 33997 41115
rect 34053 41059 34090 41115
rect 33731 40986 34090 41059
rect 34228 41091 35025 41501
rect 34228 41039 34267 41091
rect 34319 41039 34447 41091
rect 34499 41039 34627 41091
rect 34679 41039 35025 41091
rect 33019 40829 33057 40881
rect 33109 40829 33237 40881
rect 33289 40829 33327 40881
rect 33019 40789 33327 40829
rect 30770 40601 30854 40653
rect 30906 40601 31065 40653
rect 31117 40601 31276 40653
rect 31328 40601 31486 40653
rect 31538 40601 31697 40653
rect 31749 40601 31909 40653
rect 31961 40601 32120 40653
rect 32172 40601 32330 40653
rect 32382 40601 32541 40653
rect 32593 40601 32752 40653
rect 32804 40601 32889 40653
rect 30770 39755 32889 40601
rect 34228 40655 35025 41039
rect 34228 40599 34282 40655
rect 34338 40599 34493 40655
rect 34549 40599 34705 40655
rect 34761 40653 34916 40655
rect 34972 40653 35025 40655
rect 34807 40601 34916 40653
rect 34987 40601 35025 40653
rect 34761 40599 34916 40601
rect 34972 40599 35025 40601
rect 33019 40425 33327 40465
rect 33019 40373 33057 40425
rect 33109 40373 33237 40425
rect 33289 40373 33327 40425
rect 33019 40188 33327 40373
rect 33019 40132 33055 40188
rect 33111 40132 33235 40188
rect 33291 40132 33327 40188
rect 33019 39977 33327 40132
rect 33019 39925 33057 39977
rect 33109 39925 33237 39977
rect 33289 39925 33327 39977
rect 33019 39884 33327 39925
rect 33731 40195 34090 40268
rect 33731 40139 33817 40195
rect 33873 40139 33997 40195
rect 34053 40139 34090 40195
rect 33731 39969 34090 40139
rect 33731 39917 33819 39969
rect 33871 39917 33999 39969
rect 34051 39917 34090 39969
rect 33731 39876 34090 39917
rect 34228 40215 35025 40599
rect 34228 40163 34267 40215
rect 34319 40163 34447 40215
rect 34499 40163 34627 40215
rect 34679 40163 35025 40215
rect 30770 39699 30852 39755
rect 30908 39699 31063 39755
rect 31119 39699 31274 39755
rect 31330 39699 31484 39755
rect 31540 39699 31695 39755
rect 31751 39699 31907 39755
rect 31963 39699 32118 39755
rect 32174 39699 32328 39755
rect 32384 39699 32539 39755
rect 32595 39699 32750 39755
rect 32806 39699 32889 39755
rect 30770 38853 32889 39699
rect 34228 39753 35025 40163
rect 34228 39701 34284 39753
rect 34336 39701 34495 39753
rect 34547 39701 34707 39753
rect 34759 39701 34918 39753
rect 34970 39701 35025 39753
rect 33019 39529 33327 39570
rect 33019 39477 33057 39529
rect 33109 39477 33237 39529
rect 33289 39477 33327 39529
rect 33019 39322 33327 39477
rect 33019 39266 33055 39322
rect 33111 39266 33235 39322
rect 33291 39266 33327 39322
rect 33019 39081 33327 39266
rect 33731 39537 34090 39578
rect 33731 39485 33819 39537
rect 33871 39485 33999 39537
rect 34051 39485 34090 39537
rect 33731 39315 34090 39485
rect 33731 39259 33817 39315
rect 33873 39259 33997 39315
rect 34053 39259 34090 39315
rect 33731 39186 34090 39259
rect 34228 39291 35025 39701
rect 34228 39239 34267 39291
rect 34319 39239 34447 39291
rect 34499 39239 34627 39291
rect 34679 39239 35025 39291
rect 33019 39029 33057 39081
rect 33109 39029 33237 39081
rect 33289 39029 33327 39081
rect 33019 38989 33327 39029
rect 30770 38801 30854 38853
rect 30906 38801 31065 38853
rect 31117 38801 31276 38853
rect 31328 38801 31486 38853
rect 31538 38801 31697 38853
rect 31749 38801 31909 38853
rect 31961 38801 32120 38853
rect 32172 38801 32330 38853
rect 32382 38801 32541 38853
rect 32593 38801 32752 38853
rect 32804 38801 32889 38853
rect 30770 37955 32889 38801
rect 34228 38855 35025 39239
rect 34228 38799 34282 38855
rect 34338 38799 34493 38855
rect 34549 38799 34705 38855
rect 34761 38853 34916 38855
rect 34972 38853 35025 38855
rect 34807 38801 34916 38853
rect 34987 38801 35025 38853
rect 34761 38799 34916 38801
rect 34972 38799 35025 38801
rect 33019 38625 33327 38665
rect 33019 38573 33057 38625
rect 33109 38573 33237 38625
rect 33289 38573 33327 38625
rect 33019 38388 33327 38573
rect 33019 38332 33055 38388
rect 33111 38332 33235 38388
rect 33291 38332 33327 38388
rect 33019 38177 33327 38332
rect 33019 38125 33057 38177
rect 33109 38125 33237 38177
rect 33289 38125 33327 38177
rect 33019 38084 33327 38125
rect 33731 38395 34090 38468
rect 33731 38339 33817 38395
rect 33873 38339 33997 38395
rect 34053 38339 34090 38395
rect 33731 38169 34090 38339
rect 33731 38117 33819 38169
rect 33871 38117 33999 38169
rect 34051 38117 34090 38169
rect 33731 38076 34090 38117
rect 34228 38415 35025 38799
rect 34228 38363 34267 38415
rect 34319 38363 34447 38415
rect 34499 38363 34627 38415
rect 34679 38363 35025 38415
rect 30770 37899 30852 37955
rect 30908 37899 31063 37955
rect 31119 37899 31274 37955
rect 31330 37899 31484 37955
rect 31540 37899 31695 37955
rect 31751 37899 31907 37955
rect 31963 37899 32118 37955
rect 32174 37899 32328 37955
rect 32384 37899 32539 37955
rect 32595 37899 32750 37955
rect 32806 37899 32889 37955
rect 30770 37053 32889 37899
rect 34228 37953 35025 38363
rect 34228 37901 34284 37953
rect 34336 37901 34495 37953
rect 34547 37901 34707 37953
rect 34759 37901 34918 37953
rect 34970 37901 35025 37953
rect 33019 37729 33327 37770
rect 33019 37677 33057 37729
rect 33109 37677 33237 37729
rect 33289 37677 33327 37729
rect 33019 37522 33327 37677
rect 33019 37466 33055 37522
rect 33111 37466 33235 37522
rect 33291 37466 33327 37522
rect 33019 37281 33327 37466
rect 33731 37737 34090 37778
rect 33731 37685 33819 37737
rect 33871 37685 33999 37737
rect 34051 37685 34090 37737
rect 33731 37515 34090 37685
rect 33731 37459 33817 37515
rect 33873 37459 33997 37515
rect 34053 37459 34090 37515
rect 33731 37386 34090 37459
rect 34228 37491 35025 37901
rect 34228 37439 34267 37491
rect 34319 37439 34447 37491
rect 34499 37439 34627 37491
rect 34679 37439 35025 37491
rect 33019 37229 33057 37281
rect 33109 37229 33237 37281
rect 33289 37229 33327 37281
rect 33019 37189 33327 37229
rect 30770 37001 30854 37053
rect 30906 37001 31065 37053
rect 31117 37001 31276 37053
rect 31328 37001 31486 37053
rect 31538 37001 31697 37053
rect 31749 37001 31909 37053
rect 31961 37001 32120 37053
rect 32172 37001 32330 37053
rect 32382 37001 32541 37053
rect 32593 37001 32752 37053
rect 32804 37001 32889 37053
rect 30770 36155 32889 37001
rect 34228 37055 35025 37439
rect 34228 36999 34282 37055
rect 34338 36999 34493 37055
rect 34549 36999 34705 37055
rect 34761 37053 34916 37055
rect 34972 37053 35025 37055
rect 34807 37001 34916 37053
rect 34987 37001 35025 37053
rect 34761 36999 34916 37001
rect 34972 36999 35025 37001
rect 33019 36825 33327 36865
rect 33019 36773 33057 36825
rect 33109 36773 33237 36825
rect 33289 36773 33327 36825
rect 33019 36588 33327 36773
rect 33019 36532 33055 36588
rect 33111 36532 33235 36588
rect 33291 36532 33327 36588
rect 33019 36377 33327 36532
rect 33019 36325 33057 36377
rect 33109 36325 33237 36377
rect 33289 36325 33327 36377
rect 33019 36284 33327 36325
rect 33731 36595 34090 36668
rect 33731 36539 33817 36595
rect 33873 36539 33997 36595
rect 34053 36539 34090 36595
rect 33731 36369 34090 36539
rect 33731 36317 33819 36369
rect 33871 36317 33999 36369
rect 34051 36317 34090 36369
rect 33731 36276 34090 36317
rect 34228 36615 35025 36999
rect 34228 36563 34267 36615
rect 34319 36563 34447 36615
rect 34499 36563 34627 36615
rect 34679 36563 35025 36615
rect 30770 36099 30852 36155
rect 30908 36099 31063 36155
rect 31119 36099 31274 36155
rect 31330 36099 31484 36155
rect 31540 36099 31695 36155
rect 31751 36099 31907 36155
rect 31963 36099 32118 36155
rect 32174 36099 32328 36155
rect 32384 36099 32539 36155
rect 32595 36099 32750 36155
rect 32806 36099 32889 36155
rect 30770 35976 32889 36099
rect 34228 36153 35025 36563
rect 34228 36101 34284 36153
rect 34336 36101 34495 36153
rect 34547 36101 34707 36153
rect 34759 36101 34918 36153
rect 34970 36101 35025 36153
rect 34228 35976 35025 36101
rect 35131 64899 35218 64940
rect 35274 64899 35428 64955
rect 35484 64899 35639 64955
rect 35695 64899 35851 64955
rect 35907 64899 36062 64955
rect 36118 64899 36272 64955
rect 36328 64899 36415 64955
rect 36863 65372 37743 65411
rect 36863 65316 36899 65372
rect 36955 65316 37110 65372
rect 37166 65316 37321 65372
rect 37377 65316 37532 65372
rect 37588 65316 37743 65372
rect 36863 65078 37743 65316
rect 38268 65078 38863 65928
rect 38953 65601 39618 66376
rect 38953 65549 39053 65601
rect 39105 65549 39264 65601
rect 39316 65549 39475 65601
rect 39527 65549 39618 65601
rect 38953 65078 39618 65549
rect 40214 65858 40523 65928
rect 42671 65905 43222 65946
rect 40214 65855 40252 65858
rect 40304 65855 40432 65858
rect 40484 65855 40523 65858
rect 40214 65799 40250 65855
rect 40306 65799 40430 65855
rect 40486 65799 40523 65855
rect 40214 65640 40523 65799
rect 42208 65844 42548 65885
rect 42208 65792 42246 65844
rect 42298 65792 42458 65844
rect 42510 65792 42548 65844
rect 42208 65751 42548 65792
rect 42671 65853 42710 65905
rect 42762 65853 42921 65905
rect 42973 65853 43132 65905
rect 43184 65853 43222 65905
rect 40214 65588 40252 65640
rect 40304 65588 40432 65640
rect 40484 65588 40523 65640
rect 40214 65078 40523 65588
rect 40971 65372 42155 65411
rect 40971 65316 41008 65372
rect 41064 65316 41219 65372
rect 41275 65316 41430 65372
rect 41486 65316 41641 65372
rect 41697 65316 41852 65372
rect 41908 65316 42062 65372
rect 42118 65316 42155 65372
rect 40971 65277 42155 65316
rect 42671 65365 43222 65853
rect 42671 65309 42708 65365
rect 42764 65309 42919 65365
rect 42975 65309 43130 65365
rect 43186 65309 43222 65365
rect 42671 65271 43222 65309
rect 43703 65905 44564 65946
rect 43703 65853 43777 65905
rect 43829 65853 43988 65905
rect 44040 65853 44199 65905
rect 44251 65853 44410 65905
rect 44462 65853 44564 65905
rect 40717 65078 41316 65091
rect 36863 64940 37744 65078
rect 38268 64953 38864 65078
rect 38268 64940 38330 64953
rect 35131 64651 36415 64899
rect 35131 64599 35332 64651
rect 35384 64599 35543 64651
rect 35595 64599 35754 64651
rect 35806 64599 35965 64651
rect 36017 64599 36176 64651
rect 36228 64599 36415 64651
rect 35131 64191 36415 64599
rect 36640 64563 36768 64602
rect 36640 64507 36676 64563
rect 36732 64540 36768 64563
rect 36732 64507 36769 64540
rect 36640 64416 36769 64507
rect 36640 64364 36678 64416
rect 36730 64364 36769 64416
rect 36640 64323 36769 64364
rect 36864 64423 37744 64940
rect 38269 64901 38330 64940
rect 38382 64901 38541 64953
rect 38593 64901 38752 64953
rect 38804 64901 38864 64953
rect 38953 64955 39619 65078
rect 38953 64940 39050 64955
rect 36864 64371 36961 64423
rect 37013 64371 37172 64423
rect 37224 64371 37384 64423
rect 37436 64371 37595 64423
rect 37647 64371 37744 64423
rect 35131 64139 35332 64191
rect 35384 64139 35543 64191
rect 35595 64139 35754 64191
rect 35806 64139 35965 64191
rect 36017 64139 36176 64191
rect 36228 64139 36415 64191
rect 35131 63915 36415 64139
rect 35131 63863 35332 63915
rect 35384 63863 35543 63915
rect 35595 63863 35754 63915
rect 35806 63863 35965 63915
rect 36017 63863 36176 63915
rect 36228 63863 36415 63915
rect 35131 63455 36415 63863
rect 35131 63403 35332 63455
rect 35384 63403 35543 63455
rect 35595 63403 35754 63455
rect 35806 63403 35965 63455
rect 36017 63403 36176 63455
rect 36228 63403 36415 63455
rect 36640 63690 36769 63731
rect 36640 63638 36678 63690
rect 36730 63638 36769 63690
rect 36640 63547 36769 63638
rect 36640 63491 36676 63547
rect 36732 63514 36769 63547
rect 36864 63683 37744 64371
rect 37852 64663 38161 64704
rect 37852 64611 37891 64663
rect 37943 64611 38071 64663
rect 38123 64611 38161 64663
rect 37852 64332 38161 64611
rect 37852 64276 37889 64332
rect 37945 64276 38069 64332
rect 38125 64276 38161 64332
rect 37852 64189 38161 64276
rect 37852 64137 37891 64189
rect 37943 64137 38071 64189
rect 38123 64137 38161 64189
rect 37852 64096 38161 64137
rect 38269 64055 38864 64901
rect 38269 63999 38328 64055
rect 38384 63999 38539 64055
rect 38595 63999 38750 64055
rect 38806 63999 38864 64055
rect 36864 63631 36961 63683
rect 37013 63631 37172 63683
rect 37224 63631 37384 63683
rect 37436 63631 37595 63683
rect 37647 63631 37744 63683
rect 36732 63491 36768 63514
rect 36640 63452 36768 63491
rect 35131 63155 36415 63403
rect 35131 63099 35218 63155
rect 35274 63099 35428 63155
rect 35484 63099 35639 63155
rect 35695 63099 35851 63155
rect 35907 63099 36062 63155
rect 36118 63099 36272 63155
rect 36328 63099 36415 63155
rect 35131 62851 36415 63099
rect 35131 62799 35332 62851
rect 35384 62799 35543 62851
rect 35595 62799 35754 62851
rect 35806 62799 35965 62851
rect 36017 62799 36176 62851
rect 36228 62799 36415 62851
rect 35131 62391 36415 62799
rect 36640 62763 36768 62802
rect 36640 62707 36676 62763
rect 36732 62740 36768 62763
rect 36732 62707 36769 62740
rect 36640 62616 36769 62707
rect 36640 62564 36678 62616
rect 36730 62564 36769 62616
rect 36640 62523 36769 62564
rect 36864 62623 37744 63631
rect 37852 63917 38161 63958
rect 37852 63865 37891 63917
rect 37943 63865 38071 63917
rect 38123 63865 38161 63917
rect 37852 63778 38161 63865
rect 37852 63722 37889 63778
rect 37945 63722 38069 63778
rect 38125 63722 38161 63778
rect 37852 63443 38161 63722
rect 37852 63391 37891 63443
rect 37943 63391 38071 63443
rect 38123 63391 38161 63443
rect 37852 63350 38161 63391
rect 38269 63153 38864 63999
rect 38269 63101 38330 63153
rect 38382 63101 38541 63153
rect 38593 63101 38752 63153
rect 38804 63101 38864 63153
rect 36864 62571 36961 62623
rect 37013 62571 37172 62623
rect 37224 62571 37384 62623
rect 37436 62571 37595 62623
rect 37647 62571 37744 62623
rect 35131 62339 35332 62391
rect 35384 62339 35543 62391
rect 35595 62339 35754 62391
rect 35806 62339 35965 62391
rect 36017 62339 36176 62391
rect 36228 62339 36415 62391
rect 35131 62115 36415 62339
rect 35131 62063 35332 62115
rect 35384 62063 35543 62115
rect 35595 62063 35754 62115
rect 35806 62063 35965 62115
rect 36017 62063 36176 62115
rect 36228 62063 36415 62115
rect 35131 61655 36415 62063
rect 35131 61603 35332 61655
rect 35384 61603 35543 61655
rect 35595 61603 35754 61655
rect 35806 61603 35965 61655
rect 36017 61603 36176 61655
rect 36228 61603 36415 61655
rect 36640 61890 36769 61931
rect 36640 61838 36678 61890
rect 36730 61838 36769 61890
rect 36640 61747 36769 61838
rect 36640 61691 36676 61747
rect 36732 61714 36769 61747
rect 36864 61883 37744 62571
rect 37852 62863 38161 62904
rect 37852 62811 37891 62863
rect 37943 62811 38071 62863
rect 38123 62811 38161 62863
rect 37852 62532 38161 62811
rect 37852 62476 37889 62532
rect 37945 62476 38069 62532
rect 38125 62476 38161 62532
rect 37852 62389 38161 62476
rect 37852 62337 37891 62389
rect 37943 62337 38071 62389
rect 38123 62337 38161 62389
rect 37852 62296 38161 62337
rect 38269 62255 38864 63101
rect 38269 62199 38328 62255
rect 38384 62199 38539 62255
rect 38595 62199 38750 62255
rect 38806 62199 38864 62255
rect 36864 61831 36961 61883
rect 37013 61831 37172 61883
rect 37224 61831 37384 61883
rect 37436 61831 37595 61883
rect 37647 61831 37744 61883
rect 36732 61691 36768 61714
rect 36640 61652 36768 61691
rect 35131 61355 36415 61603
rect 35131 61299 35218 61355
rect 35274 61299 35428 61355
rect 35484 61299 35639 61355
rect 35695 61299 35851 61355
rect 35907 61299 36062 61355
rect 36118 61299 36272 61355
rect 36328 61299 36415 61355
rect 35131 61051 36415 61299
rect 35131 60999 35332 61051
rect 35384 60999 35543 61051
rect 35595 60999 35754 61051
rect 35806 60999 35965 61051
rect 36017 60999 36176 61051
rect 36228 60999 36415 61051
rect 35131 60591 36415 60999
rect 36640 60963 36768 61002
rect 36640 60907 36676 60963
rect 36732 60940 36768 60963
rect 36732 60907 36769 60940
rect 36640 60816 36769 60907
rect 36640 60764 36678 60816
rect 36730 60764 36769 60816
rect 36640 60723 36769 60764
rect 36864 60823 37744 61831
rect 37852 62117 38161 62158
rect 37852 62065 37891 62117
rect 37943 62065 38071 62117
rect 38123 62065 38161 62117
rect 37852 61978 38161 62065
rect 37852 61922 37889 61978
rect 37945 61922 38069 61978
rect 38125 61922 38161 61978
rect 37852 61643 38161 61922
rect 37852 61591 37891 61643
rect 37943 61591 38071 61643
rect 38123 61591 38161 61643
rect 37852 61550 38161 61591
rect 38269 61353 38864 62199
rect 38269 61301 38330 61353
rect 38382 61301 38541 61353
rect 38593 61301 38752 61353
rect 38804 61301 38864 61353
rect 36864 60771 36961 60823
rect 37013 60771 37172 60823
rect 37224 60771 37384 60823
rect 37436 60771 37595 60823
rect 37647 60771 37744 60823
rect 35131 60539 35332 60591
rect 35384 60539 35543 60591
rect 35595 60539 35754 60591
rect 35806 60539 35965 60591
rect 36017 60539 36176 60591
rect 36228 60539 36415 60591
rect 35131 60315 36415 60539
rect 35131 60263 35332 60315
rect 35384 60263 35543 60315
rect 35595 60263 35754 60315
rect 35806 60263 35965 60315
rect 36017 60263 36176 60315
rect 36228 60263 36415 60315
rect 35131 59855 36415 60263
rect 35131 59803 35332 59855
rect 35384 59803 35543 59855
rect 35595 59803 35754 59855
rect 35806 59803 35965 59855
rect 36017 59803 36176 59855
rect 36228 59803 36415 59855
rect 36640 60090 36769 60131
rect 36640 60038 36678 60090
rect 36730 60038 36769 60090
rect 36640 59947 36769 60038
rect 36640 59891 36676 59947
rect 36732 59914 36769 59947
rect 36864 60083 37744 60771
rect 37852 61063 38161 61104
rect 37852 61011 37891 61063
rect 37943 61011 38071 61063
rect 38123 61011 38161 61063
rect 37852 60732 38161 61011
rect 37852 60676 37889 60732
rect 37945 60676 38069 60732
rect 38125 60676 38161 60732
rect 37852 60589 38161 60676
rect 37852 60537 37891 60589
rect 37943 60537 38071 60589
rect 38123 60537 38161 60589
rect 37852 60496 38161 60537
rect 38269 60455 38864 61301
rect 38269 60399 38328 60455
rect 38384 60399 38539 60455
rect 38595 60399 38750 60455
rect 38806 60399 38864 60455
rect 36864 60031 36961 60083
rect 37013 60031 37172 60083
rect 37224 60031 37384 60083
rect 37436 60031 37595 60083
rect 37647 60031 37744 60083
rect 36732 59891 36768 59914
rect 36640 59852 36768 59891
rect 35131 59555 36415 59803
rect 35131 59499 35218 59555
rect 35274 59499 35428 59555
rect 35484 59499 35639 59555
rect 35695 59499 35851 59555
rect 35907 59499 36062 59555
rect 36118 59499 36272 59555
rect 36328 59499 36415 59555
rect 35131 59251 36415 59499
rect 35131 59199 35332 59251
rect 35384 59199 35543 59251
rect 35595 59199 35754 59251
rect 35806 59199 35965 59251
rect 36017 59199 36176 59251
rect 36228 59199 36415 59251
rect 35131 58791 36415 59199
rect 36640 59163 36768 59202
rect 36640 59107 36676 59163
rect 36732 59140 36768 59163
rect 36732 59107 36769 59140
rect 36640 59016 36769 59107
rect 36640 58964 36678 59016
rect 36730 58964 36769 59016
rect 36640 58923 36769 58964
rect 36864 59023 37744 60031
rect 37852 60317 38161 60358
rect 37852 60265 37891 60317
rect 37943 60265 38071 60317
rect 38123 60265 38161 60317
rect 37852 60178 38161 60265
rect 37852 60122 37889 60178
rect 37945 60122 38069 60178
rect 38125 60122 38161 60178
rect 37852 59843 38161 60122
rect 37852 59791 37891 59843
rect 37943 59791 38071 59843
rect 38123 59791 38161 59843
rect 37852 59750 38161 59791
rect 38269 59553 38864 60399
rect 38269 59501 38330 59553
rect 38382 59501 38541 59553
rect 38593 59501 38752 59553
rect 38804 59501 38864 59553
rect 36864 58971 36961 59023
rect 37013 58971 37172 59023
rect 37224 58971 37384 59023
rect 37436 58971 37595 59023
rect 37647 58971 37744 59023
rect 35131 58739 35332 58791
rect 35384 58739 35543 58791
rect 35595 58739 35754 58791
rect 35806 58739 35965 58791
rect 36017 58739 36176 58791
rect 36228 58739 36415 58791
rect 35131 58515 36415 58739
rect 35131 58463 35332 58515
rect 35384 58463 35543 58515
rect 35595 58463 35754 58515
rect 35806 58463 35965 58515
rect 36017 58463 36176 58515
rect 36228 58463 36415 58515
rect 35131 58055 36415 58463
rect 35131 58003 35332 58055
rect 35384 58003 35543 58055
rect 35595 58003 35754 58055
rect 35806 58003 35965 58055
rect 36017 58003 36176 58055
rect 36228 58003 36415 58055
rect 36640 58290 36769 58331
rect 36640 58238 36678 58290
rect 36730 58238 36769 58290
rect 36640 58147 36769 58238
rect 36640 58091 36676 58147
rect 36732 58114 36769 58147
rect 36864 58283 37744 58971
rect 37852 59263 38161 59304
rect 37852 59211 37891 59263
rect 37943 59211 38071 59263
rect 38123 59211 38161 59263
rect 37852 58932 38161 59211
rect 37852 58876 37889 58932
rect 37945 58876 38069 58932
rect 38125 58876 38161 58932
rect 37852 58789 38161 58876
rect 37852 58737 37891 58789
rect 37943 58737 38071 58789
rect 38123 58737 38161 58789
rect 37852 58696 38161 58737
rect 38269 58655 38864 59501
rect 38269 58599 38328 58655
rect 38384 58599 38539 58655
rect 38595 58599 38750 58655
rect 38806 58599 38864 58655
rect 36864 58231 36961 58283
rect 37013 58231 37172 58283
rect 37224 58231 37384 58283
rect 37436 58231 37595 58283
rect 37647 58231 37744 58283
rect 36732 58091 36768 58114
rect 36640 58052 36768 58091
rect 35131 57755 36415 58003
rect 35131 57699 35218 57755
rect 35274 57699 35428 57755
rect 35484 57699 35639 57755
rect 35695 57699 35851 57755
rect 35907 57699 36062 57755
rect 36118 57699 36272 57755
rect 36328 57699 36415 57755
rect 35131 57451 36415 57699
rect 35131 57399 35332 57451
rect 35384 57399 35543 57451
rect 35595 57399 35754 57451
rect 35806 57399 35965 57451
rect 36017 57399 36176 57451
rect 36228 57399 36415 57451
rect 35131 56991 36415 57399
rect 36640 57363 36768 57402
rect 36640 57307 36676 57363
rect 36732 57340 36768 57363
rect 36732 57307 36769 57340
rect 36640 57216 36769 57307
rect 36640 57164 36678 57216
rect 36730 57164 36769 57216
rect 36640 57123 36769 57164
rect 36864 57223 37744 58231
rect 37852 58517 38161 58558
rect 37852 58465 37891 58517
rect 37943 58465 38071 58517
rect 38123 58465 38161 58517
rect 37852 58378 38161 58465
rect 37852 58322 37889 58378
rect 37945 58322 38069 58378
rect 38125 58322 38161 58378
rect 37852 58043 38161 58322
rect 37852 57991 37891 58043
rect 37943 57991 38071 58043
rect 38123 57991 38161 58043
rect 37852 57950 38161 57991
rect 38269 57753 38864 58599
rect 38269 57701 38330 57753
rect 38382 57701 38541 57753
rect 38593 57701 38752 57753
rect 38804 57701 38864 57753
rect 36864 57171 36961 57223
rect 37013 57171 37172 57223
rect 37224 57171 37384 57223
rect 37436 57171 37595 57223
rect 37647 57171 37744 57223
rect 35131 56939 35332 56991
rect 35384 56939 35543 56991
rect 35595 56939 35754 56991
rect 35806 56939 35965 56991
rect 36017 56939 36176 56991
rect 36228 56939 36415 56991
rect 35131 56715 36415 56939
rect 35131 56663 35332 56715
rect 35384 56663 35543 56715
rect 35595 56663 35754 56715
rect 35806 56663 35965 56715
rect 36017 56663 36176 56715
rect 36228 56663 36415 56715
rect 35131 56255 36415 56663
rect 35131 56203 35332 56255
rect 35384 56203 35543 56255
rect 35595 56203 35754 56255
rect 35806 56203 35965 56255
rect 36017 56203 36176 56255
rect 36228 56203 36415 56255
rect 36640 56490 36769 56531
rect 36640 56438 36678 56490
rect 36730 56438 36769 56490
rect 36640 56347 36769 56438
rect 36640 56291 36676 56347
rect 36732 56314 36769 56347
rect 36864 56483 37744 57171
rect 37852 57463 38161 57504
rect 37852 57411 37891 57463
rect 37943 57411 38071 57463
rect 38123 57411 38161 57463
rect 37852 57132 38161 57411
rect 37852 57076 37889 57132
rect 37945 57076 38069 57132
rect 38125 57076 38161 57132
rect 37852 56989 38161 57076
rect 37852 56937 37891 56989
rect 37943 56937 38071 56989
rect 38123 56937 38161 56989
rect 37852 56896 38161 56937
rect 38269 56855 38864 57701
rect 38269 56799 38328 56855
rect 38384 56799 38539 56855
rect 38595 56799 38750 56855
rect 38806 56799 38864 56855
rect 36864 56431 36961 56483
rect 37013 56431 37172 56483
rect 37224 56431 37384 56483
rect 37436 56431 37595 56483
rect 37647 56431 37744 56483
rect 36732 56291 36768 56314
rect 36640 56252 36768 56291
rect 35131 55955 36415 56203
rect 35131 55899 35218 55955
rect 35274 55899 35428 55955
rect 35484 55899 35639 55955
rect 35695 55899 35851 55955
rect 35907 55899 36062 55955
rect 36118 55899 36272 55955
rect 36328 55899 36415 55955
rect 35131 55651 36415 55899
rect 35131 55599 35332 55651
rect 35384 55599 35543 55651
rect 35595 55599 35754 55651
rect 35806 55599 35965 55651
rect 36017 55599 36176 55651
rect 36228 55599 36415 55651
rect 35131 55191 36415 55599
rect 36640 55563 36768 55602
rect 36640 55507 36676 55563
rect 36732 55540 36768 55563
rect 36732 55507 36769 55540
rect 36640 55416 36769 55507
rect 36640 55364 36678 55416
rect 36730 55364 36769 55416
rect 36640 55323 36769 55364
rect 36864 55423 37744 56431
rect 37852 56717 38161 56758
rect 37852 56665 37891 56717
rect 37943 56665 38071 56717
rect 38123 56665 38161 56717
rect 37852 56578 38161 56665
rect 37852 56522 37889 56578
rect 37945 56522 38069 56578
rect 38125 56522 38161 56578
rect 37852 56243 38161 56522
rect 37852 56191 37891 56243
rect 37943 56191 38071 56243
rect 38123 56191 38161 56243
rect 37852 56150 38161 56191
rect 38269 55953 38864 56799
rect 38269 55901 38330 55953
rect 38382 55901 38541 55953
rect 38593 55901 38752 55953
rect 38804 55901 38864 55953
rect 36864 55371 36961 55423
rect 37013 55371 37172 55423
rect 37224 55371 37384 55423
rect 37436 55371 37595 55423
rect 37647 55371 37744 55423
rect 35131 55139 35332 55191
rect 35384 55139 35543 55191
rect 35595 55139 35754 55191
rect 35806 55139 35965 55191
rect 36017 55139 36176 55191
rect 36228 55139 36415 55191
rect 35131 54915 36415 55139
rect 35131 54863 35332 54915
rect 35384 54863 35543 54915
rect 35595 54863 35754 54915
rect 35806 54863 35965 54915
rect 36017 54863 36176 54915
rect 36228 54863 36415 54915
rect 35131 54455 36415 54863
rect 35131 54403 35332 54455
rect 35384 54403 35543 54455
rect 35595 54403 35754 54455
rect 35806 54403 35965 54455
rect 36017 54403 36176 54455
rect 36228 54403 36415 54455
rect 36640 54690 36769 54731
rect 36640 54638 36678 54690
rect 36730 54638 36769 54690
rect 36640 54547 36769 54638
rect 36640 54491 36676 54547
rect 36732 54514 36769 54547
rect 36864 54683 37744 55371
rect 37852 55663 38161 55704
rect 37852 55611 37891 55663
rect 37943 55611 38071 55663
rect 38123 55611 38161 55663
rect 37852 55332 38161 55611
rect 37852 55276 37889 55332
rect 37945 55276 38069 55332
rect 38125 55276 38161 55332
rect 37852 55189 38161 55276
rect 37852 55137 37891 55189
rect 37943 55137 38071 55189
rect 38123 55137 38161 55189
rect 37852 55096 38161 55137
rect 38269 55055 38864 55901
rect 38269 54999 38328 55055
rect 38384 54999 38539 55055
rect 38595 54999 38750 55055
rect 38806 54999 38864 55055
rect 36864 54631 36961 54683
rect 37013 54631 37172 54683
rect 37224 54631 37384 54683
rect 37436 54631 37595 54683
rect 37647 54631 37744 54683
rect 36732 54491 36768 54514
rect 36640 54452 36768 54491
rect 35131 54155 36415 54403
rect 35131 54099 35218 54155
rect 35274 54099 35428 54155
rect 35484 54099 35639 54155
rect 35695 54099 35851 54155
rect 35907 54099 36062 54155
rect 36118 54099 36272 54155
rect 36328 54099 36415 54155
rect 35131 53851 36415 54099
rect 35131 53799 35332 53851
rect 35384 53799 35543 53851
rect 35595 53799 35754 53851
rect 35806 53799 35965 53851
rect 36017 53799 36176 53851
rect 36228 53799 36415 53851
rect 35131 53391 36415 53799
rect 36640 53763 36768 53802
rect 36640 53707 36676 53763
rect 36732 53740 36768 53763
rect 36732 53707 36769 53740
rect 36640 53616 36769 53707
rect 36640 53564 36678 53616
rect 36730 53564 36769 53616
rect 36640 53523 36769 53564
rect 36864 53623 37744 54631
rect 37852 54917 38161 54958
rect 37852 54865 37891 54917
rect 37943 54865 38071 54917
rect 38123 54865 38161 54917
rect 37852 54778 38161 54865
rect 37852 54722 37889 54778
rect 37945 54722 38069 54778
rect 38125 54722 38161 54778
rect 37852 54443 38161 54722
rect 37852 54391 37891 54443
rect 37943 54391 38071 54443
rect 38123 54391 38161 54443
rect 37852 54350 38161 54391
rect 38269 54153 38864 54999
rect 38269 54101 38330 54153
rect 38382 54101 38541 54153
rect 38593 54101 38752 54153
rect 38804 54101 38864 54153
rect 36864 53571 36961 53623
rect 37013 53571 37172 53623
rect 37224 53571 37384 53623
rect 37436 53571 37595 53623
rect 37647 53571 37744 53623
rect 35131 53339 35332 53391
rect 35384 53339 35543 53391
rect 35595 53339 35754 53391
rect 35806 53339 35965 53391
rect 36017 53339 36176 53391
rect 36228 53339 36415 53391
rect 35131 53115 36415 53339
rect 35131 53063 35332 53115
rect 35384 53063 35543 53115
rect 35595 53063 35754 53115
rect 35806 53063 35965 53115
rect 36017 53063 36176 53115
rect 36228 53063 36415 53115
rect 35131 52655 36415 53063
rect 35131 52603 35332 52655
rect 35384 52603 35543 52655
rect 35595 52603 35754 52655
rect 35806 52603 35965 52655
rect 36017 52603 36176 52655
rect 36228 52603 36415 52655
rect 36640 52890 36769 52931
rect 36640 52838 36678 52890
rect 36730 52838 36769 52890
rect 36640 52747 36769 52838
rect 36640 52691 36676 52747
rect 36732 52714 36769 52747
rect 36864 52883 37744 53571
rect 37852 53863 38161 53904
rect 37852 53811 37891 53863
rect 37943 53811 38071 53863
rect 38123 53811 38161 53863
rect 37852 53532 38161 53811
rect 37852 53476 37889 53532
rect 37945 53476 38069 53532
rect 38125 53476 38161 53532
rect 37852 53389 38161 53476
rect 37852 53337 37891 53389
rect 37943 53337 38071 53389
rect 38123 53337 38161 53389
rect 37852 53296 38161 53337
rect 38269 53255 38864 54101
rect 38269 53199 38328 53255
rect 38384 53199 38539 53255
rect 38595 53199 38750 53255
rect 38806 53199 38864 53255
rect 36864 52831 36961 52883
rect 37013 52831 37172 52883
rect 37224 52831 37384 52883
rect 37436 52831 37595 52883
rect 37647 52831 37744 52883
rect 36732 52691 36768 52714
rect 36640 52652 36768 52691
rect 35131 52355 36415 52603
rect 35131 52299 35218 52355
rect 35274 52299 35428 52355
rect 35484 52299 35639 52355
rect 35695 52299 35851 52355
rect 35907 52299 36062 52355
rect 36118 52299 36272 52355
rect 36328 52299 36415 52355
rect 35131 52051 36415 52299
rect 35131 51999 35332 52051
rect 35384 51999 35543 52051
rect 35595 51999 35754 52051
rect 35806 51999 35965 52051
rect 36017 51999 36176 52051
rect 36228 51999 36415 52051
rect 35131 51591 36415 51999
rect 36640 51963 36768 52002
rect 36640 51907 36676 51963
rect 36732 51940 36768 51963
rect 36732 51907 36769 51940
rect 36640 51816 36769 51907
rect 36640 51764 36678 51816
rect 36730 51764 36769 51816
rect 36640 51723 36769 51764
rect 36864 51823 37744 52831
rect 37852 53117 38161 53158
rect 37852 53065 37891 53117
rect 37943 53065 38071 53117
rect 38123 53065 38161 53117
rect 37852 52978 38161 53065
rect 37852 52922 37889 52978
rect 37945 52922 38069 52978
rect 38125 52922 38161 52978
rect 37852 52643 38161 52922
rect 37852 52591 37891 52643
rect 37943 52591 38071 52643
rect 38123 52591 38161 52643
rect 37852 52550 38161 52591
rect 38269 52353 38864 53199
rect 38269 52301 38330 52353
rect 38382 52301 38541 52353
rect 38593 52301 38752 52353
rect 38804 52301 38864 52353
rect 36864 51771 36961 51823
rect 37013 51771 37172 51823
rect 37224 51771 37384 51823
rect 37436 51771 37595 51823
rect 37647 51771 37744 51823
rect 35131 51539 35332 51591
rect 35384 51539 35543 51591
rect 35595 51539 35754 51591
rect 35806 51539 35965 51591
rect 36017 51539 36176 51591
rect 36228 51539 36415 51591
rect 35131 51315 36415 51539
rect 35131 51263 35332 51315
rect 35384 51263 35543 51315
rect 35595 51263 35754 51315
rect 35806 51263 35965 51315
rect 36017 51263 36176 51315
rect 36228 51263 36415 51315
rect 35131 50855 36415 51263
rect 35131 50803 35332 50855
rect 35384 50803 35543 50855
rect 35595 50803 35754 50855
rect 35806 50803 35965 50855
rect 36017 50803 36176 50855
rect 36228 50803 36415 50855
rect 36640 51090 36769 51131
rect 36640 51038 36678 51090
rect 36730 51038 36769 51090
rect 36640 50947 36769 51038
rect 36640 50891 36676 50947
rect 36732 50914 36769 50947
rect 36864 51083 37744 51771
rect 37852 52063 38161 52104
rect 37852 52011 37891 52063
rect 37943 52011 38071 52063
rect 38123 52011 38161 52063
rect 37852 51732 38161 52011
rect 37852 51676 37889 51732
rect 37945 51676 38069 51732
rect 38125 51676 38161 51732
rect 37852 51589 38161 51676
rect 37852 51537 37891 51589
rect 37943 51537 38071 51589
rect 38123 51537 38161 51589
rect 37852 51496 38161 51537
rect 38269 51455 38864 52301
rect 38269 51399 38328 51455
rect 38384 51399 38539 51455
rect 38595 51399 38750 51455
rect 38806 51399 38864 51455
rect 36864 51031 36961 51083
rect 37013 51031 37172 51083
rect 37224 51031 37384 51083
rect 37436 51031 37595 51083
rect 37647 51031 37744 51083
rect 36732 50891 36768 50914
rect 36640 50852 36768 50891
rect 35131 50555 36415 50803
rect 35131 50499 35218 50555
rect 35274 50499 35428 50555
rect 35484 50499 35639 50555
rect 35695 50499 35851 50555
rect 35907 50499 36062 50555
rect 36118 50499 36272 50555
rect 36328 50499 36415 50555
rect 35131 50251 36415 50499
rect 35131 50199 35332 50251
rect 35384 50199 35543 50251
rect 35595 50199 35754 50251
rect 35806 50199 35965 50251
rect 36017 50199 36176 50251
rect 36228 50199 36415 50251
rect 35131 49791 36415 50199
rect 36640 50163 36768 50202
rect 36640 50107 36676 50163
rect 36732 50140 36768 50163
rect 36732 50107 36769 50140
rect 36640 50016 36769 50107
rect 36640 49964 36678 50016
rect 36730 49964 36769 50016
rect 36640 49923 36769 49964
rect 36864 50023 37744 51031
rect 37852 51317 38161 51358
rect 37852 51265 37891 51317
rect 37943 51265 38071 51317
rect 38123 51265 38161 51317
rect 37852 51178 38161 51265
rect 37852 51122 37889 51178
rect 37945 51122 38069 51178
rect 38125 51122 38161 51178
rect 37852 50843 38161 51122
rect 37852 50791 37891 50843
rect 37943 50791 38071 50843
rect 38123 50791 38161 50843
rect 37852 50750 38161 50791
rect 38269 50553 38864 51399
rect 38269 50501 38330 50553
rect 38382 50501 38541 50553
rect 38593 50501 38752 50553
rect 38804 50501 38864 50553
rect 36864 49971 36961 50023
rect 37013 49971 37172 50023
rect 37224 49971 37384 50023
rect 37436 49971 37595 50023
rect 37647 49971 37744 50023
rect 35131 49739 35332 49791
rect 35384 49739 35543 49791
rect 35595 49739 35754 49791
rect 35806 49739 35965 49791
rect 36017 49739 36176 49791
rect 36228 49739 36415 49791
rect 35131 49515 36415 49739
rect 35131 49463 35332 49515
rect 35384 49463 35543 49515
rect 35595 49463 35754 49515
rect 35806 49463 35965 49515
rect 36017 49463 36176 49515
rect 36228 49463 36415 49515
rect 35131 49055 36415 49463
rect 35131 49003 35332 49055
rect 35384 49003 35543 49055
rect 35595 49003 35754 49055
rect 35806 49003 35965 49055
rect 36017 49003 36176 49055
rect 36228 49003 36415 49055
rect 36640 49290 36769 49331
rect 36640 49238 36678 49290
rect 36730 49238 36769 49290
rect 36640 49147 36769 49238
rect 36640 49091 36676 49147
rect 36732 49114 36769 49147
rect 36864 49283 37744 49971
rect 37852 50263 38161 50304
rect 37852 50211 37891 50263
rect 37943 50211 38071 50263
rect 38123 50211 38161 50263
rect 37852 49932 38161 50211
rect 37852 49876 37889 49932
rect 37945 49876 38069 49932
rect 38125 49876 38161 49932
rect 37852 49789 38161 49876
rect 37852 49737 37891 49789
rect 37943 49737 38071 49789
rect 38123 49737 38161 49789
rect 37852 49696 38161 49737
rect 38269 49655 38864 50501
rect 38269 49599 38328 49655
rect 38384 49599 38539 49655
rect 38595 49599 38750 49655
rect 38806 49599 38864 49655
rect 36864 49231 36961 49283
rect 37013 49231 37172 49283
rect 37224 49231 37384 49283
rect 37436 49231 37595 49283
rect 37647 49231 37744 49283
rect 36732 49091 36768 49114
rect 36640 49052 36768 49091
rect 35131 48755 36415 49003
rect 35131 48699 35218 48755
rect 35274 48699 35428 48755
rect 35484 48699 35639 48755
rect 35695 48699 35851 48755
rect 35907 48699 36062 48755
rect 36118 48699 36272 48755
rect 36328 48699 36415 48755
rect 35131 48451 36415 48699
rect 35131 48399 35332 48451
rect 35384 48399 35543 48451
rect 35595 48399 35754 48451
rect 35806 48399 35965 48451
rect 36017 48399 36176 48451
rect 36228 48399 36415 48451
rect 35131 47991 36415 48399
rect 36640 48363 36768 48402
rect 36640 48307 36676 48363
rect 36732 48340 36768 48363
rect 36732 48307 36769 48340
rect 36640 48216 36769 48307
rect 36640 48164 36678 48216
rect 36730 48164 36769 48216
rect 36640 48123 36769 48164
rect 36864 48223 37744 49231
rect 37852 49517 38161 49558
rect 37852 49465 37891 49517
rect 37943 49465 38071 49517
rect 38123 49465 38161 49517
rect 37852 49378 38161 49465
rect 37852 49322 37889 49378
rect 37945 49322 38069 49378
rect 38125 49322 38161 49378
rect 37852 49043 38161 49322
rect 37852 48991 37891 49043
rect 37943 48991 38071 49043
rect 38123 48991 38161 49043
rect 37852 48950 38161 48991
rect 38269 48753 38864 49599
rect 38269 48701 38330 48753
rect 38382 48701 38541 48753
rect 38593 48701 38752 48753
rect 38804 48701 38864 48753
rect 36864 48171 36961 48223
rect 37013 48171 37172 48223
rect 37224 48171 37384 48223
rect 37436 48171 37595 48223
rect 37647 48171 37744 48223
rect 35131 47939 35332 47991
rect 35384 47939 35543 47991
rect 35595 47939 35754 47991
rect 35806 47939 35965 47991
rect 36017 47939 36176 47991
rect 36228 47939 36415 47991
rect 35131 47715 36415 47939
rect 35131 47663 35332 47715
rect 35384 47663 35543 47715
rect 35595 47663 35754 47715
rect 35806 47663 35965 47715
rect 36017 47663 36176 47715
rect 36228 47663 36415 47715
rect 35131 47255 36415 47663
rect 35131 47203 35332 47255
rect 35384 47203 35543 47255
rect 35595 47203 35754 47255
rect 35806 47203 35965 47255
rect 36017 47203 36176 47255
rect 36228 47203 36415 47255
rect 36640 47490 36769 47531
rect 36640 47438 36678 47490
rect 36730 47438 36769 47490
rect 36640 47347 36769 47438
rect 36640 47291 36676 47347
rect 36732 47314 36769 47347
rect 36864 47483 37744 48171
rect 37852 48463 38161 48504
rect 37852 48411 37891 48463
rect 37943 48411 38071 48463
rect 38123 48411 38161 48463
rect 37852 48132 38161 48411
rect 37852 48076 37889 48132
rect 37945 48076 38069 48132
rect 38125 48076 38161 48132
rect 37852 47989 38161 48076
rect 37852 47937 37891 47989
rect 37943 47937 38071 47989
rect 38123 47937 38161 47989
rect 37852 47896 38161 47937
rect 38269 47855 38864 48701
rect 38269 47799 38328 47855
rect 38384 47799 38539 47855
rect 38595 47799 38750 47855
rect 38806 47799 38864 47855
rect 36864 47431 36961 47483
rect 37013 47431 37172 47483
rect 37224 47431 37384 47483
rect 37436 47431 37595 47483
rect 37647 47431 37744 47483
rect 36732 47291 36768 47314
rect 36640 47252 36768 47291
rect 35131 46955 36415 47203
rect 35131 46899 35218 46955
rect 35274 46899 35428 46955
rect 35484 46899 35639 46955
rect 35695 46899 35851 46955
rect 35907 46899 36062 46955
rect 36118 46899 36272 46955
rect 36328 46899 36415 46955
rect 35131 46651 36415 46899
rect 35131 46599 35332 46651
rect 35384 46599 35543 46651
rect 35595 46599 35754 46651
rect 35806 46599 35965 46651
rect 36017 46599 36176 46651
rect 36228 46599 36415 46651
rect 35131 46191 36415 46599
rect 36640 46563 36768 46602
rect 36640 46507 36676 46563
rect 36732 46540 36768 46563
rect 36732 46507 36769 46540
rect 36640 46416 36769 46507
rect 36640 46364 36678 46416
rect 36730 46364 36769 46416
rect 36640 46323 36769 46364
rect 36864 46423 37744 47431
rect 37852 47717 38161 47758
rect 37852 47665 37891 47717
rect 37943 47665 38071 47717
rect 38123 47665 38161 47717
rect 37852 47578 38161 47665
rect 37852 47522 37889 47578
rect 37945 47522 38069 47578
rect 38125 47522 38161 47578
rect 37852 47243 38161 47522
rect 37852 47191 37891 47243
rect 37943 47191 38071 47243
rect 38123 47191 38161 47243
rect 37852 47150 38161 47191
rect 38269 46953 38864 47799
rect 38269 46901 38330 46953
rect 38382 46901 38541 46953
rect 38593 46901 38752 46953
rect 38804 46901 38864 46953
rect 36864 46371 36961 46423
rect 37013 46371 37172 46423
rect 37224 46371 37384 46423
rect 37436 46371 37595 46423
rect 37647 46371 37744 46423
rect 35131 46139 35332 46191
rect 35384 46139 35543 46191
rect 35595 46139 35754 46191
rect 35806 46139 35965 46191
rect 36017 46139 36176 46191
rect 36228 46139 36415 46191
rect 35131 45915 36415 46139
rect 35131 45863 35332 45915
rect 35384 45863 35543 45915
rect 35595 45863 35754 45915
rect 35806 45863 35965 45915
rect 36017 45863 36176 45915
rect 36228 45863 36415 45915
rect 35131 45455 36415 45863
rect 35131 45403 35332 45455
rect 35384 45403 35543 45455
rect 35595 45403 35754 45455
rect 35806 45403 35965 45455
rect 36017 45403 36176 45455
rect 36228 45403 36415 45455
rect 36640 45690 36769 45731
rect 36640 45638 36678 45690
rect 36730 45638 36769 45690
rect 36640 45547 36769 45638
rect 36640 45491 36676 45547
rect 36732 45514 36769 45547
rect 36864 45683 37744 46371
rect 37852 46663 38161 46704
rect 37852 46611 37891 46663
rect 37943 46611 38071 46663
rect 38123 46611 38161 46663
rect 37852 46332 38161 46611
rect 37852 46276 37889 46332
rect 37945 46276 38069 46332
rect 38125 46276 38161 46332
rect 37852 46189 38161 46276
rect 37852 46137 37891 46189
rect 37943 46137 38071 46189
rect 38123 46137 38161 46189
rect 37852 46096 38161 46137
rect 38269 46055 38864 46901
rect 38269 45999 38328 46055
rect 38384 45999 38539 46055
rect 38595 45999 38750 46055
rect 38806 45999 38864 46055
rect 36864 45631 36961 45683
rect 37013 45631 37172 45683
rect 37224 45631 37384 45683
rect 37436 45631 37595 45683
rect 37647 45631 37744 45683
rect 36732 45491 36768 45514
rect 36640 45452 36768 45491
rect 35131 45155 36415 45403
rect 35131 45099 35218 45155
rect 35274 45099 35428 45155
rect 35484 45099 35639 45155
rect 35695 45099 35851 45155
rect 35907 45099 36062 45155
rect 36118 45099 36272 45155
rect 36328 45099 36415 45155
rect 35131 44851 36415 45099
rect 35131 44799 35332 44851
rect 35384 44799 35543 44851
rect 35595 44799 35754 44851
rect 35806 44799 35965 44851
rect 36017 44799 36176 44851
rect 36228 44799 36415 44851
rect 35131 44391 36415 44799
rect 36640 44763 36768 44802
rect 36640 44707 36676 44763
rect 36732 44740 36768 44763
rect 36732 44707 36769 44740
rect 36640 44616 36769 44707
rect 36640 44564 36678 44616
rect 36730 44564 36769 44616
rect 36640 44523 36769 44564
rect 36864 44623 37744 45631
rect 37852 45917 38161 45958
rect 37852 45865 37891 45917
rect 37943 45865 38071 45917
rect 38123 45865 38161 45917
rect 37852 45778 38161 45865
rect 37852 45722 37889 45778
rect 37945 45722 38069 45778
rect 38125 45722 38161 45778
rect 37852 45443 38161 45722
rect 37852 45391 37891 45443
rect 37943 45391 38071 45443
rect 38123 45391 38161 45443
rect 37852 45350 38161 45391
rect 38269 45153 38864 45999
rect 38269 45101 38330 45153
rect 38382 45101 38541 45153
rect 38593 45101 38752 45153
rect 38804 45101 38864 45153
rect 36864 44571 36961 44623
rect 37013 44571 37172 44623
rect 37224 44571 37384 44623
rect 37436 44571 37595 44623
rect 37647 44571 37744 44623
rect 35131 44339 35332 44391
rect 35384 44339 35543 44391
rect 35595 44339 35754 44391
rect 35806 44339 35965 44391
rect 36017 44339 36176 44391
rect 36228 44339 36415 44391
rect 35131 44115 36415 44339
rect 35131 44063 35332 44115
rect 35384 44063 35543 44115
rect 35595 44063 35754 44115
rect 35806 44063 35965 44115
rect 36017 44063 36176 44115
rect 36228 44063 36415 44115
rect 35131 43655 36415 44063
rect 35131 43603 35332 43655
rect 35384 43603 35543 43655
rect 35595 43603 35754 43655
rect 35806 43603 35965 43655
rect 36017 43603 36176 43655
rect 36228 43603 36415 43655
rect 36640 43890 36769 43931
rect 36640 43838 36678 43890
rect 36730 43838 36769 43890
rect 36640 43747 36769 43838
rect 36640 43691 36676 43747
rect 36732 43714 36769 43747
rect 36864 43883 37744 44571
rect 37852 44863 38161 44904
rect 37852 44811 37891 44863
rect 37943 44811 38071 44863
rect 38123 44811 38161 44863
rect 37852 44532 38161 44811
rect 37852 44476 37889 44532
rect 37945 44476 38069 44532
rect 38125 44476 38161 44532
rect 37852 44389 38161 44476
rect 37852 44337 37891 44389
rect 37943 44337 38071 44389
rect 38123 44337 38161 44389
rect 37852 44296 38161 44337
rect 38269 44255 38864 45101
rect 38269 44199 38328 44255
rect 38384 44199 38539 44255
rect 38595 44199 38750 44255
rect 38806 44199 38864 44255
rect 36864 43831 36961 43883
rect 37013 43831 37172 43883
rect 37224 43831 37384 43883
rect 37436 43831 37595 43883
rect 37647 43831 37744 43883
rect 36732 43691 36768 43714
rect 36640 43652 36768 43691
rect 35131 43355 36415 43603
rect 35131 43299 35218 43355
rect 35274 43299 35428 43355
rect 35484 43299 35639 43355
rect 35695 43299 35851 43355
rect 35907 43299 36062 43355
rect 36118 43299 36272 43355
rect 36328 43299 36415 43355
rect 35131 43051 36415 43299
rect 35131 42999 35332 43051
rect 35384 42999 35543 43051
rect 35595 42999 35754 43051
rect 35806 42999 35965 43051
rect 36017 42999 36176 43051
rect 36228 42999 36415 43051
rect 35131 42591 36415 42999
rect 36640 42963 36768 43002
rect 36640 42907 36676 42963
rect 36732 42940 36768 42963
rect 36732 42907 36769 42940
rect 36640 42816 36769 42907
rect 36640 42764 36678 42816
rect 36730 42764 36769 42816
rect 36640 42723 36769 42764
rect 36864 42823 37744 43831
rect 37852 44117 38161 44158
rect 37852 44065 37891 44117
rect 37943 44065 38071 44117
rect 38123 44065 38161 44117
rect 37852 43978 38161 44065
rect 37852 43922 37889 43978
rect 37945 43922 38069 43978
rect 38125 43922 38161 43978
rect 37852 43643 38161 43922
rect 37852 43591 37891 43643
rect 37943 43591 38071 43643
rect 38123 43591 38161 43643
rect 37852 43550 38161 43591
rect 38269 43353 38864 44199
rect 38269 43301 38330 43353
rect 38382 43301 38541 43353
rect 38593 43301 38752 43353
rect 38804 43301 38864 43353
rect 36864 42771 36961 42823
rect 37013 42771 37172 42823
rect 37224 42771 37384 42823
rect 37436 42771 37595 42823
rect 37647 42771 37744 42823
rect 35131 42539 35332 42591
rect 35384 42539 35543 42591
rect 35595 42539 35754 42591
rect 35806 42539 35965 42591
rect 36017 42539 36176 42591
rect 36228 42539 36415 42591
rect 35131 42315 36415 42539
rect 35131 42263 35332 42315
rect 35384 42263 35543 42315
rect 35595 42263 35754 42315
rect 35806 42263 35965 42315
rect 36017 42263 36176 42315
rect 36228 42263 36415 42315
rect 35131 41855 36415 42263
rect 35131 41803 35332 41855
rect 35384 41803 35543 41855
rect 35595 41803 35754 41855
rect 35806 41803 35965 41855
rect 36017 41803 36176 41855
rect 36228 41803 36415 41855
rect 36640 42090 36769 42131
rect 36640 42038 36678 42090
rect 36730 42038 36769 42090
rect 36640 41947 36769 42038
rect 36640 41891 36676 41947
rect 36732 41914 36769 41947
rect 36864 42083 37744 42771
rect 37852 43063 38161 43104
rect 37852 43011 37891 43063
rect 37943 43011 38071 43063
rect 38123 43011 38161 43063
rect 37852 42732 38161 43011
rect 37852 42676 37889 42732
rect 37945 42676 38069 42732
rect 38125 42676 38161 42732
rect 37852 42589 38161 42676
rect 37852 42537 37891 42589
rect 37943 42537 38071 42589
rect 38123 42537 38161 42589
rect 37852 42496 38161 42537
rect 38269 42455 38864 43301
rect 38269 42399 38328 42455
rect 38384 42399 38539 42455
rect 38595 42399 38750 42455
rect 38806 42399 38864 42455
rect 36864 42031 36961 42083
rect 37013 42031 37172 42083
rect 37224 42031 37384 42083
rect 37436 42031 37595 42083
rect 37647 42031 37744 42083
rect 36732 41891 36768 41914
rect 36640 41852 36768 41891
rect 35131 41555 36415 41803
rect 35131 41499 35218 41555
rect 35274 41499 35428 41555
rect 35484 41499 35639 41555
rect 35695 41499 35851 41555
rect 35907 41499 36062 41555
rect 36118 41499 36272 41555
rect 36328 41499 36415 41555
rect 35131 41251 36415 41499
rect 35131 41199 35332 41251
rect 35384 41199 35543 41251
rect 35595 41199 35754 41251
rect 35806 41199 35965 41251
rect 36017 41199 36176 41251
rect 36228 41199 36415 41251
rect 35131 40791 36415 41199
rect 36640 41163 36768 41202
rect 36640 41107 36676 41163
rect 36732 41140 36768 41163
rect 36732 41107 36769 41140
rect 36640 41016 36769 41107
rect 36640 40964 36678 41016
rect 36730 40964 36769 41016
rect 36640 40923 36769 40964
rect 36864 41023 37744 42031
rect 37852 42317 38161 42358
rect 37852 42265 37891 42317
rect 37943 42265 38071 42317
rect 38123 42265 38161 42317
rect 37852 42178 38161 42265
rect 37852 42122 37889 42178
rect 37945 42122 38069 42178
rect 38125 42122 38161 42178
rect 37852 41843 38161 42122
rect 37852 41791 37891 41843
rect 37943 41791 38071 41843
rect 38123 41791 38161 41843
rect 37852 41750 38161 41791
rect 38269 41553 38864 42399
rect 38269 41501 38330 41553
rect 38382 41501 38541 41553
rect 38593 41501 38752 41553
rect 38804 41501 38864 41553
rect 36864 40971 36961 41023
rect 37013 40971 37172 41023
rect 37224 40971 37384 41023
rect 37436 40971 37595 41023
rect 37647 40971 37744 41023
rect 35131 40739 35332 40791
rect 35384 40739 35543 40791
rect 35595 40739 35754 40791
rect 35806 40739 35965 40791
rect 36017 40739 36176 40791
rect 36228 40739 36415 40791
rect 35131 40515 36415 40739
rect 35131 40463 35332 40515
rect 35384 40463 35543 40515
rect 35595 40463 35754 40515
rect 35806 40463 35965 40515
rect 36017 40463 36176 40515
rect 36228 40463 36415 40515
rect 35131 40055 36415 40463
rect 35131 40003 35332 40055
rect 35384 40003 35543 40055
rect 35595 40003 35754 40055
rect 35806 40003 35965 40055
rect 36017 40003 36176 40055
rect 36228 40003 36415 40055
rect 36640 40290 36769 40331
rect 36640 40238 36678 40290
rect 36730 40238 36769 40290
rect 36640 40147 36769 40238
rect 36640 40091 36676 40147
rect 36732 40114 36769 40147
rect 36864 40283 37744 40971
rect 37852 41263 38161 41304
rect 37852 41211 37891 41263
rect 37943 41211 38071 41263
rect 38123 41211 38161 41263
rect 37852 40932 38161 41211
rect 37852 40876 37889 40932
rect 37945 40876 38069 40932
rect 38125 40876 38161 40932
rect 37852 40789 38161 40876
rect 37852 40737 37891 40789
rect 37943 40737 38071 40789
rect 38123 40737 38161 40789
rect 37852 40696 38161 40737
rect 38269 40655 38864 41501
rect 38269 40599 38328 40655
rect 38384 40599 38539 40655
rect 38595 40599 38750 40655
rect 38806 40599 38864 40655
rect 36864 40231 36961 40283
rect 37013 40231 37172 40283
rect 37224 40231 37384 40283
rect 37436 40231 37595 40283
rect 37647 40231 37744 40283
rect 36732 40091 36768 40114
rect 36640 40052 36768 40091
rect 35131 39755 36415 40003
rect 35131 39699 35218 39755
rect 35274 39699 35428 39755
rect 35484 39699 35639 39755
rect 35695 39699 35851 39755
rect 35907 39699 36062 39755
rect 36118 39699 36272 39755
rect 36328 39699 36415 39755
rect 35131 39451 36415 39699
rect 35131 39399 35332 39451
rect 35384 39399 35543 39451
rect 35595 39399 35754 39451
rect 35806 39399 35965 39451
rect 36017 39399 36176 39451
rect 36228 39399 36415 39451
rect 35131 38991 36415 39399
rect 36640 39363 36768 39402
rect 36640 39307 36676 39363
rect 36732 39340 36768 39363
rect 36732 39307 36769 39340
rect 36640 39216 36769 39307
rect 36640 39164 36678 39216
rect 36730 39164 36769 39216
rect 36640 39123 36769 39164
rect 36864 39223 37744 40231
rect 37852 40517 38161 40558
rect 37852 40465 37891 40517
rect 37943 40465 38071 40517
rect 38123 40465 38161 40517
rect 37852 40378 38161 40465
rect 37852 40322 37889 40378
rect 37945 40322 38069 40378
rect 38125 40322 38161 40378
rect 37852 40043 38161 40322
rect 37852 39991 37891 40043
rect 37943 39991 38071 40043
rect 38123 39991 38161 40043
rect 37852 39950 38161 39991
rect 38269 39753 38864 40599
rect 38269 39701 38330 39753
rect 38382 39701 38541 39753
rect 38593 39701 38752 39753
rect 38804 39701 38864 39753
rect 36864 39171 36961 39223
rect 37013 39171 37172 39223
rect 37224 39171 37384 39223
rect 37436 39171 37595 39223
rect 37647 39171 37744 39223
rect 35131 38939 35332 38991
rect 35384 38939 35543 38991
rect 35595 38939 35754 38991
rect 35806 38939 35965 38991
rect 36017 38939 36176 38991
rect 36228 38939 36415 38991
rect 35131 38715 36415 38939
rect 35131 38663 35332 38715
rect 35384 38663 35543 38715
rect 35595 38663 35754 38715
rect 35806 38663 35965 38715
rect 36017 38663 36176 38715
rect 36228 38663 36415 38715
rect 35131 38255 36415 38663
rect 35131 38203 35332 38255
rect 35384 38203 35543 38255
rect 35595 38203 35754 38255
rect 35806 38203 35965 38255
rect 36017 38203 36176 38255
rect 36228 38203 36415 38255
rect 36640 38490 36769 38531
rect 36640 38438 36678 38490
rect 36730 38438 36769 38490
rect 36640 38347 36769 38438
rect 36640 38291 36676 38347
rect 36732 38314 36769 38347
rect 36864 38483 37744 39171
rect 37852 39463 38161 39504
rect 37852 39411 37891 39463
rect 37943 39411 38071 39463
rect 38123 39411 38161 39463
rect 37852 39132 38161 39411
rect 37852 39076 37889 39132
rect 37945 39076 38069 39132
rect 38125 39076 38161 39132
rect 37852 38989 38161 39076
rect 37852 38937 37891 38989
rect 37943 38937 38071 38989
rect 38123 38937 38161 38989
rect 37852 38896 38161 38937
rect 38269 38855 38864 39701
rect 38269 38799 38328 38855
rect 38384 38799 38539 38855
rect 38595 38799 38750 38855
rect 38806 38799 38864 38855
rect 36864 38431 36961 38483
rect 37013 38431 37172 38483
rect 37224 38431 37384 38483
rect 37436 38431 37595 38483
rect 37647 38431 37744 38483
rect 36732 38291 36768 38314
rect 36640 38252 36768 38291
rect 35131 37955 36415 38203
rect 35131 37899 35218 37955
rect 35274 37899 35428 37955
rect 35484 37899 35639 37955
rect 35695 37899 35851 37955
rect 35907 37899 36062 37955
rect 36118 37899 36272 37955
rect 36328 37899 36415 37955
rect 35131 37651 36415 37899
rect 35131 37599 35332 37651
rect 35384 37599 35543 37651
rect 35595 37599 35754 37651
rect 35806 37599 35965 37651
rect 36017 37599 36176 37651
rect 36228 37599 36415 37651
rect 35131 37191 36415 37599
rect 36640 37563 36768 37602
rect 36640 37507 36676 37563
rect 36732 37540 36768 37563
rect 36732 37507 36769 37540
rect 36640 37416 36769 37507
rect 36640 37364 36678 37416
rect 36730 37364 36769 37416
rect 36640 37323 36769 37364
rect 36864 37423 37744 38431
rect 37852 38717 38161 38758
rect 37852 38665 37891 38717
rect 37943 38665 38071 38717
rect 38123 38665 38161 38717
rect 37852 38578 38161 38665
rect 37852 38522 37889 38578
rect 37945 38522 38069 38578
rect 38125 38522 38161 38578
rect 37852 38243 38161 38522
rect 37852 38191 37891 38243
rect 37943 38191 38071 38243
rect 38123 38191 38161 38243
rect 37852 38150 38161 38191
rect 38269 37953 38864 38799
rect 38269 37901 38330 37953
rect 38382 37901 38541 37953
rect 38593 37901 38752 37953
rect 38804 37901 38864 37953
rect 36864 37371 36961 37423
rect 37013 37371 37172 37423
rect 37224 37371 37384 37423
rect 37436 37371 37595 37423
rect 37647 37371 37744 37423
rect 35131 37139 35332 37191
rect 35384 37139 35543 37191
rect 35595 37139 35754 37191
rect 35806 37139 35965 37191
rect 36017 37139 36176 37191
rect 36228 37139 36415 37191
rect 35131 36915 36415 37139
rect 35131 36863 35332 36915
rect 35384 36863 35543 36915
rect 35595 36863 35754 36915
rect 35806 36863 35965 36915
rect 36017 36863 36176 36915
rect 36228 36863 36415 36915
rect 35131 36455 36415 36863
rect 35131 36403 35332 36455
rect 35384 36403 35543 36455
rect 35595 36403 35754 36455
rect 35806 36403 35965 36455
rect 36017 36403 36176 36455
rect 36228 36403 36415 36455
rect 36640 36690 36769 36731
rect 36640 36638 36678 36690
rect 36730 36638 36769 36690
rect 36864 36683 37744 37371
rect 37852 37663 38161 37704
rect 37852 37611 37891 37663
rect 37943 37611 38071 37663
rect 38123 37611 38161 37663
rect 37852 37332 38161 37611
rect 37852 37276 37889 37332
rect 37945 37276 38069 37332
rect 38125 37276 38161 37332
rect 37852 37189 38161 37276
rect 37852 37137 37891 37189
rect 37943 37137 38071 37189
rect 38123 37137 38161 37189
rect 37852 37096 38161 37137
rect 38269 37055 38864 37901
rect 38269 36999 38328 37055
rect 38384 36999 38539 37055
rect 38595 36999 38750 37055
rect 38806 36999 38864 37055
rect 36864 36650 36961 36683
rect 36640 36547 36769 36638
rect 36640 36491 36676 36547
rect 36732 36514 36769 36547
rect 36863 36631 36961 36650
rect 37013 36631 37172 36683
rect 37224 36631 37384 36683
rect 37436 36631 37595 36683
rect 37647 36631 37744 36683
rect 36732 36491 36768 36514
rect 36640 36452 36768 36491
rect 35131 36155 36415 36403
rect 35131 36099 35218 36155
rect 35274 36099 35428 36155
rect 35484 36099 35639 36155
rect 35695 36099 35851 36155
rect 35907 36099 36062 36155
rect 36118 36099 36272 36155
rect 36328 36099 36415 36155
rect 35131 35976 36415 36099
rect 36863 35976 37744 36631
rect 37852 36917 38161 36958
rect 37852 36865 37891 36917
rect 37943 36865 38071 36917
rect 38123 36865 38161 36917
rect 37852 36778 38161 36865
rect 37852 36722 37889 36778
rect 37945 36722 38069 36778
rect 38125 36722 38161 36778
rect 37852 36443 38161 36722
rect 37852 36391 37891 36443
rect 37943 36391 38071 36443
rect 38123 36391 38161 36443
rect 37852 36350 38161 36391
rect 38269 36153 38864 36999
rect 38269 36101 38330 36153
rect 38382 36101 38541 36153
rect 38593 36101 38752 36153
rect 38804 36101 38864 36153
rect 38269 35976 38864 36101
rect 38967 64899 39050 64940
rect 39106 64899 39230 64955
rect 39286 64899 39619 64955
rect 40214 64953 40524 65078
rect 40214 64940 40253 64953
rect 38967 63155 39619 64899
rect 40215 64901 40253 64940
rect 40305 64901 40433 64953
rect 40485 64901 40524 64953
rect 39736 64715 39865 64756
rect 39736 64663 39775 64715
rect 39827 64663 39865 64715
rect 39736 64332 39865 64663
rect 39736 64276 39773 64332
rect 39829 64276 39865 64332
rect 39736 64237 39865 64276
rect 39956 64563 40084 64602
rect 39956 64507 39992 64563
rect 40048 64541 40084 64563
rect 40048 64507 40085 64541
rect 39956 64500 40085 64507
rect 39956 64448 39994 64500
rect 40046 64448 40085 64500
rect 39956 64314 40085 64448
rect 39956 64262 39994 64314
rect 40046 64262 40085 64314
rect 39956 64221 40085 64262
rect 40215 64055 40524 64901
rect 40717 64955 41317 65078
rect 40717 64899 40777 64955
rect 40833 64899 40988 64955
rect 41044 64899 41199 64955
rect 41255 64899 41317 64955
rect 40717 64826 41317 64899
rect 40215 63999 40251 64055
rect 40307 63999 40431 64055
rect 40487 63999 40524 64055
rect 39736 63778 39865 63817
rect 39736 63722 39773 63778
rect 39829 63722 39865 63778
rect 39736 63391 39865 63722
rect 39956 63792 40085 63833
rect 39956 63740 39994 63792
rect 40046 63740 40085 63792
rect 39956 63606 40085 63740
rect 39956 63554 39994 63606
rect 40046 63554 40085 63606
rect 39956 63547 40085 63554
rect 39956 63491 39992 63547
rect 40048 63513 40085 63547
rect 40048 63491 40084 63513
rect 39956 63452 40084 63491
rect 39736 63339 39775 63391
rect 39827 63339 39865 63391
rect 39736 63298 39865 63339
rect 38967 63099 39050 63155
rect 39106 63099 39230 63155
rect 39286 63099 39619 63155
rect 38967 61355 39619 63099
rect 40215 63153 40524 63999
rect 40215 63101 40253 63153
rect 40305 63101 40433 63153
rect 40485 63101 40524 63153
rect 39736 62915 39865 62956
rect 39736 62863 39775 62915
rect 39827 62863 39865 62915
rect 39736 62532 39865 62863
rect 39736 62476 39773 62532
rect 39829 62476 39865 62532
rect 39736 62437 39865 62476
rect 39956 62763 40084 62802
rect 39956 62707 39992 62763
rect 40048 62741 40084 62763
rect 40048 62707 40085 62741
rect 39956 62700 40085 62707
rect 39956 62648 39994 62700
rect 40046 62648 40085 62700
rect 39956 62514 40085 62648
rect 39956 62462 39994 62514
rect 40046 62462 40085 62514
rect 39956 62421 40085 62462
rect 40215 62255 40524 63101
rect 40215 62199 40251 62255
rect 40307 62199 40431 62255
rect 40487 62199 40524 62255
rect 39736 61978 39865 62017
rect 39736 61922 39773 61978
rect 39829 61922 39865 61978
rect 39736 61591 39865 61922
rect 39956 61992 40085 62033
rect 39956 61940 39994 61992
rect 40046 61940 40085 61992
rect 39956 61806 40085 61940
rect 39956 61754 39994 61806
rect 40046 61754 40085 61806
rect 39956 61747 40085 61754
rect 39956 61691 39992 61747
rect 40048 61713 40085 61747
rect 40048 61691 40084 61713
rect 39956 61652 40084 61691
rect 39736 61539 39775 61591
rect 39827 61539 39865 61591
rect 39736 61498 39865 61539
rect 38967 61299 39050 61355
rect 39106 61299 39230 61355
rect 39286 61299 39619 61355
rect 38967 59555 39619 61299
rect 40215 61353 40524 62199
rect 40215 61301 40253 61353
rect 40305 61301 40433 61353
rect 40485 61301 40524 61353
rect 39736 61115 39865 61156
rect 39736 61063 39775 61115
rect 39827 61063 39865 61115
rect 39736 60732 39865 61063
rect 39736 60676 39773 60732
rect 39829 60676 39865 60732
rect 39736 60637 39865 60676
rect 39956 60963 40084 61002
rect 39956 60907 39992 60963
rect 40048 60941 40084 60963
rect 40048 60907 40085 60941
rect 39956 60900 40085 60907
rect 39956 60848 39994 60900
rect 40046 60848 40085 60900
rect 39956 60714 40085 60848
rect 39956 60662 39994 60714
rect 40046 60662 40085 60714
rect 39956 60621 40085 60662
rect 40215 60455 40524 61301
rect 40215 60399 40251 60455
rect 40307 60399 40431 60455
rect 40487 60399 40524 60455
rect 39736 60178 39865 60217
rect 39736 60122 39773 60178
rect 39829 60122 39865 60178
rect 39736 59791 39865 60122
rect 39956 60192 40085 60233
rect 39956 60140 39994 60192
rect 40046 60140 40085 60192
rect 39956 60006 40085 60140
rect 39956 59954 39994 60006
rect 40046 59954 40085 60006
rect 39956 59947 40085 59954
rect 39956 59891 39992 59947
rect 40048 59913 40085 59947
rect 40048 59891 40084 59913
rect 39956 59852 40084 59891
rect 39736 59739 39775 59791
rect 39827 59739 39865 59791
rect 39736 59698 39865 59739
rect 38967 59499 39050 59555
rect 39106 59499 39230 59555
rect 39286 59499 39619 59555
rect 38967 57755 39619 59499
rect 40215 59553 40524 60399
rect 40215 59501 40253 59553
rect 40305 59501 40433 59553
rect 40485 59501 40524 59553
rect 39736 59315 39865 59356
rect 39736 59263 39775 59315
rect 39827 59263 39865 59315
rect 39736 58932 39865 59263
rect 39736 58876 39773 58932
rect 39829 58876 39865 58932
rect 39736 58837 39865 58876
rect 39956 59163 40084 59202
rect 39956 59107 39992 59163
rect 40048 59141 40084 59163
rect 40048 59107 40085 59141
rect 39956 59100 40085 59107
rect 39956 59048 39994 59100
rect 40046 59048 40085 59100
rect 39956 58914 40085 59048
rect 39956 58862 39994 58914
rect 40046 58862 40085 58914
rect 39956 58821 40085 58862
rect 40215 58655 40524 59501
rect 40215 58599 40251 58655
rect 40307 58599 40431 58655
rect 40487 58599 40524 58655
rect 39736 58378 39865 58417
rect 39736 58322 39773 58378
rect 39829 58322 39865 58378
rect 39736 57991 39865 58322
rect 39956 58392 40085 58433
rect 39956 58340 39994 58392
rect 40046 58340 40085 58392
rect 39956 58206 40085 58340
rect 39956 58154 39994 58206
rect 40046 58154 40085 58206
rect 39956 58147 40085 58154
rect 39956 58091 39992 58147
rect 40048 58113 40085 58147
rect 40048 58091 40084 58113
rect 39956 58052 40084 58091
rect 39736 57939 39775 57991
rect 39827 57939 39865 57991
rect 39736 57898 39865 57939
rect 38967 57699 39050 57755
rect 39106 57699 39230 57755
rect 39286 57699 39619 57755
rect 38967 55955 39619 57699
rect 40215 57753 40524 58599
rect 40215 57701 40253 57753
rect 40305 57701 40433 57753
rect 40485 57701 40524 57753
rect 39736 57515 39865 57556
rect 39736 57463 39775 57515
rect 39827 57463 39865 57515
rect 39736 57132 39865 57463
rect 39736 57076 39773 57132
rect 39829 57076 39865 57132
rect 39736 57037 39865 57076
rect 39956 57363 40084 57402
rect 39956 57307 39992 57363
rect 40048 57341 40084 57363
rect 40048 57307 40085 57341
rect 39956 57300 40085 57307
rect 39956 57248 39994 57300
rect 40046 57248 40085 57300
rect 39956 57114 40085 57248
rect 39956 57062 39994 57114
rect 40046 57062 40085 57114
rect 39956 57021 40085 57062
rect 40215 56855 40524 57701
rect 40215 56799 40251 56855
rect 40307 56799 40431 56855
rect 40487 56799 40524 56855
rect 39736 56578 39865 56617
rect 39736 56522 39773 56578
rect 39829 56522 39865 56578
rect 39736 56191 39865 56522
rect 39956 56592 40085 56633
rect 39956 56540 39994 56592
rect 40046 56540 40085 56592
rect 39956 56406 40085 56540
rect 39956 56354 39994 56406
rect 40046 56354 40085 56406
rect 39956 56347 40085 56354
rect 39956 56291 39992 56347
rect 40048 56313 40085 56347
rect 40048 56291 40084 56313
rect 39956 56252 40084 56291
rect 39736 56139 39775 56191
rect 39827 56139 39865 56191
rect 39736 56098 39865 56139
rect 38967 55899 39050 55955
rect 39106 55899 39230 55955
rect 39286 55899 39619 55955
rect 38967 54155 39619 55899
rect 40215 55953 40524 56799
rect 40215 55901 40253 55953
rect 40305 55901 40433 55953
rect 40485 55901 40524 55953
rect 39736 55715 39865 55756
rect 39736 55663 39775 55715
rect 39827 55663 39865 55715
rect 39736 55332 39865 55663
rect 39736 55276 39773 55332
rect 39829 55276 39865 55332
rect 39736 55237 39865 55276
rect 39956 55563 40084 55602
rect 39956 55507 39992 55563
rect 40048 55541 40084 55563
rect 40048 55507 40085 55541
rect 39956 55500 40085 55507
rect 39956 55448 39994 55500
rect 40046 55448 40085 55500
rect 39956 55314 40085 55448
rect 39956 55262 39994 55314
rect 40046 55262 40085 55314
rect 39956 55221 40085 55262
rect 40215 55055 40524 55901
rect 40215 54999 40251 55055
rect 40307 54999 40431 55055
rect 40487 54999 40524 55055
rect 39736 54778 39865 54817
rect 39736 54722 39773 54778
rect 39829 54722 39865 54778
rect 39736 54391 39865 54722
rect 39956 54792 40085 54833
rect 39956 54740 39994 54792
rect 40046 54740 40085 54792
rect 39956 54606 40085 54740
rect 39956 54554 39994 54606
rect 40046 54554 40085 54606
rect 39956 54547 40085 54554
rect 39956 54491 39992 54547
rect 40048 54513 40085 54547
rect 40048 54491 40084 54513
rect 39956 54452 40084 54491
rect 39736 54339 39775 54391
rect 39827 54339 39865 54391
rect 39736 54298 39865 54339
rect 38967 54099 39050 54155
rect 39106 54099 39230 54155
rect 39286 54099 39619 54155
rect 38967 52355 39619 54099
rect 40215 54153 40524 54999
rect 40215 54101 40253 54153
rect 40305 54101 40433 54153
rect 40485 54101 40524 54153
rect 39736 53915 39865 53956
rect 39736 53863 39775 53915
rect 39827 53863 39865 53915
rect 39736 53532 39865 53863
rect 39736 53476 39773 53532
rect 39829 53476 39865 53532
rect 39736 53437 39865 53476
rect 39956 53763 40084 53802
rect 39956 53707 39992 53763
rect 40048 53741 40084 53763
rect 40048 53707 40085 53741
rect 39956 53700 40085 53707
rect 39956 53648 39994 53700
rect 40046 53648 40085 53700
rect 39956 53514 40085 53648
rect 39956 53462 39994 53514
rect 40046 53462 40085 53514
rect 39956 53421 40085 53462
rect 40215 53255 40524 54101
rect 40215 53199 40251 53255
rect 40307 53199 40431 53255
rect 40487 53199 40524 53255
rect 39736 52978 39865 53017
rect 39736 52922 39773 52978
rect 39829 52922 39865 52978
rect 39736 52591 39865 52922
rect 39956 52992 40085 53033
rect 39956 52940 39994 52992
rect 40046 52940 40085 52992
rect 39956 52806 40085 52940
rect 39956 52754 39994 52806
rect 40046 52754 40085 52806
rect 39956 52747 40085 52754
rect 39956 52691 39992 52747
rect 40048 52713 40085 52747
rect 40048 52691 40084 52713
rect 39956 52652 40084 52691
rect 39736 52539 39775 52591
rect 39827 52539 39865 52591
rect 39736 52498 39865 52539
rect 38967 52299 39050 52355
rect 39106 52299 39230 52355
rect 39286 52299 39619 52355
rect 38967 50555 39619 52299
rect 40215 52353 40524 53199
rect 40215 52301 40253 52353
rect 40305 52301 40433 52353
rect 40485 52301 40524 52353
rect 39736 52115 39865 52156
rect 39736 52063 39775 52115
rect 39827 52063 39865 52115
rect 39736 51732 39865 52063
rect 39736 51676 39773 51732
rect 39829 51676 39865 51732
rect 39736 51637 39865 51676
rect 39956 51963 40084 52002
rect 39956 51907 39992 51963
rect 40048 51941 40084 51963
rect 40048 51907 40085 51941
rect 39956 51900 40085 51907
rect 39956 51848 39994 51900
rect 40046 51848 40085 51900
rect 39956 51714 40085 51848
rect 39956 51662 39994 51714
rect 40046 51662 40085 51714
rect 39956 51621 40085 51662
rect 40215 51455 40524 52301
rect 40215 51399 40251 51455
rect 40307 51399 40431 51455
rect 40487 51399 40524 51455
rect 39736 51178 39865 51217
rect 39736 51122 39773 51178
rect 39829 51122 39865 51178
rect 39736 50791 39865 51122
rect 39956 51192 40085 51233
rect 39956 51140 39994 51192
rect 40046 51140 40085 51192
rect 39956 51006 40085 51140
rect 39956 50954 39994 51006
rect 40046 50954 40085 51006
rect 39956 50947 40085 50954
rect 39956 50891 39992 50947
rect 40048 50913 40085 50947
rect 40048 50891 40084 50913
rect 39956 50852 40084 50891
rect 39736 50739 39775 50791
rect 39827 50739 39865 50791
rect 39736 50698 39865 50739
rect 38967 50499 39050 50555
rect 39106 50499 39230 50555
rect 39286 50499 39619 50555
rect 38967 48755 39619 50499
rect 40215 50553 40524 51399
rect 40215 50501 40253 50553
rect 40305 50501 40433 50553
rect 40485 50501 40524 50553
rect 39736 50315 39865 50356
rect 39736 50263 39775 50315
rect 39827 50263 39865 50315
rect 39736 49932 39865 50263
rect 39736 49876 39773 49932
rect 39829 49876 39865 49932
rect 39736 49837 39865 49876
rect 39956 50163 40084 50202
rect 39956 50107 39992 50163
rect 40048 50141 40084 50163
rect 40048 50107 40085 50141
rect 39956 50100 40085 50107
rect 39956 50048 39994 50100
rect 40046 50048 40085 50100
rect 39956 49914 40085 50048
rect 39956 49862 39994 49914
rect 40046 49862 40085 49914
rect 39956 49821 40085 49862
rect 40215 49655 40524 50501
rect 40215 49599 40251 49655
rect 40307 49599 40431 49655
rect 40487 49599 40524 49655
rect 39736 49378 39865 49417
rect 39736 49322 39773 49378
rect 39829 49322 39865 49378
rect 39736 48991 39865 49322
rect 39956 49392 40085 49433
rect 39956 49340 39994 49392
rect 40046 49340 40085 49392
rect 39956 49206 40085 49340
rect 39956 49154 39994 49206
rect 40046 49154 40085 49206
rect 39956 49147 40085 49154
rect 39956 49091 39992 49147
rect 40048 49113 40085 49147
rect 40048 49091 40084 49113
rect 39956 49052 40084 49091
rect 39736 48939 39775 48991
rect 39827 48939 39865 48991
rect 39736 48898 39865 48939
rect 38967 48699 39050 48755
rect 39106 48699 39230 48755
rect 39286 48699 39619 48755
rect 38967 46955 39619 48699
rect 40215 48753 40524 49599
rect 40215 48701 40253 48753
rect 40305 48701 40433 48753
rect 40485 48701 40524 48753
rect 39736 48515 39865 48556
rect 39736 48463 39775 48515
rect 39827 48463 39865 48515
rect 39736 48132 39865 48463
rect 39736 48076 39773 48132
rect 39829 48076 39865 48132
rect 39736 48037 39865 48076
rect 39956 48363 40084 48402
rect 39956 48307 39992 48363
rect 40048 48341 40084 48363
rect 40048 48307 40085 48341
rect 39956 48300 40085 48307
rect 39956 48248 39994 48300
rect 40046 48248 40085 48300
rect 39956 48114 40085 48248
rect 39956 48062 39994 48114
rect 40046 48062 40085 48114
rect 39956 48021 40085 48062
rect 40215 47855 40524 48701
rect 40215 47799 40251 47855
rect 40307 47799 40431 47855
rect 40487 47799 40524 47855
rect 39736 47578 39865 47617
rect 39736 47522 39773 47578
rect 39829 47522 39865 47578
rect 39736 47191 39865 47522
rect 39956 47592 40085 47633
rect 39956 47540 39994 47592
rect 40046 47540 40085 47592
rect 39956 47406 40085 47540
rect 39956 47354 39994 47406
rect 40046 47354 40085 47406
rect 39956 47347 40085 47354
rect 39956 47291 39992 47347
rect 40048 47313 40085 47347
rect 40048 47291 40084 47313
rect 39956 47252 40084 47291
rect 39736 47139 39775 47191
rect 39827 47139 39865 47191
rect 39736 47098 39865 47139
rect 38967 46899 39050 46955
rect 39106 46899 39230 46955
rect 39286 46899 39619 46955
rect 38967 45155 39619 46899
rect 40215 46953 40524 47799
rect 40215 46901 40253 46953
rect 40305 46901 40433 46953
rect 40485 46901 40524 46953
rect 39736 46715 39865 46756
rect 39736 46663 39775 46715
rect 39827 46663 39865 46715
rect 39736 46332 39865 46663
rect 39736 46276 39773 46332
rect 39829 46276 39865 46332
rect 39736 46237 39865 46276
rect 39956 46563 40084 46602
rect 39956 46507 39992 46563
rect 40048 46541 40084 46563
rect 40048 46507 40085 46541
rect 39956 46500 40085 46507
rect 39956 46448 39994 46500
rect 40046 46448 40085 46500
rect 39956 46314 40085 46448
rect 39956 46262 39994 46314
rect 40046 46262 40085 46314
rect 39956 46221 40085 46262
rect 40215 46055 40524 46901
rect 40215 45999 40251 46055
rect 40307 45999 40431 46055
rect 40487 45999 40524 46055
rect 39736 45778 39865 45817
rect 39736 45722 39773 45778
rect 39829 45722 39865 45778
rect 39736 45391 39865 45722
rect 39956 45792 40085 45833
rect 39956 45740 39994 45792
rect 40046 45740 40085 45792
rect 39956 45606 40085 45740
rect 39956 45554 39994 45606
rect 40046 45554 40085 45606
rect 39956 45547 40085 45554
rect 39956 45491 39992 45547
rect 40048 45513 40085 45547
rect 40048 45491 40084 45513
rect 39956 45452 40084 45491
rect 39736 45339 39775 45391
rect 39827 45339 39865 45391
rect 39736 45298 39865 45339
rect 38967 45099 39050 45155
rect 39106 45099 39230 45155
rect 39286 45099 39619 45155
rect 38967 43355 39619 45099
rect 40215 45153 40524 45999
rect 40215 45101 40253 45153
rect 40305 45101 40433 45153
rect 40485 45101 40524 45153
rect 39736 44915 39865 44956
rect 39736 44863 39775 44915
rect 39827 44863 39865 44915
rect 39736 44532 39865 44863
rect 39736 44476 39773 44532
rect 39829 44476 39865 44532
rect 39736 44437 39865 44476
rect 39956 44763 40084 44802
rect 39956 44707 39992 44763
rect 40048 44741 40084 44763
rect 40048 44707 40085 44741
rect 39956 44700 40085 44707
rect 39956 44648 39994 44700
rect 40046 44648 40085 44700
rect 39956 44514 40085 44648
rect 39956 44462 39994 44514
rect 40046 44462 40085 44514
rect 39956 44421 40085 44462
rect 40215 44255 40524 45101
rect 40215 44199 40251 44255
rect 40307 44199 40431 44255
rect 40487 44199 40524 44255
rect 39736 43978 39865 44017
rect 39736 43922 39773 43978
rect 39829 43922 39865 43978
rect 39736 43591 39865 43922
rect 39956 43992 40085 44033
rect 39956 43940 39994 43992
rect 40046 43940 40085 43992
rect 39956 43806 40085 43940
rect 39956 43754 39994 43806
rect 40046 43754 40085 43806
rect 39956 43747 40085 43754
rect 39956 43691 39992 43747
rect 40048 43713 40085 43747
rect 40048 43691 40084 43713
rect 39956 43652 40084 43691
rect 39736 43539 39775 43591
rect 39827 43539 39865 43591
rect 39736 43498 39865 43539
rect 38967 43299 39050 43355
rect 39106 43299 39230 43355
rect 39286 43299 39619 43355
rect 38967 41555 39619 43299
rect 40215 43353 40524 44199
rect 40215 43301 40253 43353
rect 40305 43301 40433 43353
rect 40485 43301 40524 43353
rect 39736 43115 39865 43156
rect 39736 43063 39775 43115
rect 39827 43063 39865 43115
rect 39736 42732 39865 43063
rect 39736 42676 39773 42732
rect 39829 42676 39865 42732
rect 39736 42637 39865 42676
rect 39956 42963 40084 43002
rect 39956 42907 39992 42963
rect 40048 42941 40084 42963
rect 40048 42907 40085 42941
rect 39956 42900 40085 42907
rect 39956 42848 39994 42900
rect 40046 42848 40085 42900
rect 39956 42714 40085 42848
rect 39956 42662 39994 42714
rect 40046 42662 40085 42714
rect 39956 42621 40085 42662
rect 40215 42455 40524 43301
rect 40215 42399 40251 42455
rect 40307 42399 40431 42455
rect 40487 42399 40524 42455
rect 39736 42178 39865 42217
rect 39736 42122 39773 42178
rect 39829 42122 39865 42178
rect 39736 41791 39865 42122
rect 39956 42192 40085 42233
rect 39956 42140 39994 42192
rect 40046 42140 40085 42192
rect 39956 42006 40085 42140
rect 39956 41954 39994 42006
rect 40046 41954 40085 42006
rect 39956 41947 40085 41954
rect 39956 41891 39992 41947
rect 40048 41913 40085 41947
rect 40048 41891 40084 41913
rect 39956 41852 40084 41891
rect 39736 41739 39775 41791
rect 39827 41739 39865 41791
rect 39736 41698 39865 41739
rect 38967 41499 39050 41555
rect 39106 41499 39230 41555
rect 39286 41499 39619 41555
rect 38967 39755 39619 41499
rect 40215 41553 40524 42399
rect 40215 41501 40253 41553
rect 40305 41501 40433 41553
rect 40485 41501 40524 41553
rect 39736 41315 39865 41356
rect 39736 41263 39775 41315
rect 39827 41263 39865 41315
rect 39736 40932 39865 41263
rect 39736 40876 39773 40932
rect 39829 40876 39865 40932
rect 39736 40837 39865 40876
rect 39956 41163 40084 41202
rect 39956 41107 39992 41163
rect 40048 41141 40084 41163
rect 40048 41107 40085 41141
rect 39956 41100 40085 41107
rect 39956 41048 39994 41100
rect 40046 41048 40085 41100
rect 39956 40914 40085 41048
rect 39956 40862 39994 40914
rect 40046 40862 40085 40914
rect 39956 40821 40085 40862
rect 40215 40655 40524 41501
rect 40215 40599 40251 40655
rect 40307 40599 40431 40655
rect 40487 40599 40524 40655
rect 39736 40378 39865 40417
rect 39736 40322 39773 40378
rect 39829 40322 39865 40378
rect 39736 39991 39865 40322
rect 39956 40392 40085 40433
rect 39956 40340 39994 40392
rect 40046 40340 40085 40392
rect 39956 40206 40085 40340
rect 39956 40154 39994 40206
rect 40046 40154 40085 40206
rect 39956 40147 40085 40154
rect 39956 40091 39992 40147
rect 40048 40113 40085 40147
rect 40048 40091 40084 40113
rect 39956 40052 40084 40091
rect 39736 39939 39775 39991
rect 39827 39939 39865 39991
rect 39736 39898 39865 39939
rect 38967 39699 39050 39755
rect 39106 39699 39230 39755
rect 39286 39699 39619 39755
rect 38967 37955 39619 39699
rect 40215 39753 40524 40599
rect 40215 39701 40253 39753
rect 40305 39701 40433 39753
rect 40485 39701 40524 39753
rect 39736 39515 39865 39556
rect 39736 39463 39775 39515
rect 39827 39463 39865 39515
rect 39736 39132 39865 39463
rect 39736 39076 39773 39132
rect 39829 39076 39865 39132
rect 39736 39037 39865 39076
rect 39956 39363 40084 39402
rect 39956 39307 39992 39363
rect 40048 39341 40084 39363
rect 40048 39307 40085 39341
rect 39956 39300 40085 39307
rect 39956 39248 39994 39300
rect 40046 39248 40085 39300
rect 39956 39114 40085 39248
rect 39956 39062 39994 39114
rect 40046 39062 40085 39114
rect 39956 39021 40085 39062
rect 40215 38855 40524 39701
rect 40215 38799 40251 38855
rect 40307 38799 40431 38855
rect 40487 38799 40524 38855
rect 39736 38578 39865 38617
rect 39736 38522 39773 38578
rect 39829 38522 39865 38578
rect 39736 38191 39865 38522
rect 39956 38592 40085 38633
rect 39956 38540 39994 38592
rect 40046 38540 40085 38592
rect 39956 38406 40085 38540
rect 39956 38354 39994 38406
rect 40046 38354 40085 38406
rect 39956 38347 40085 38354
rect 39956 38291 39992 38347
rect 40048 38313 40085 38347
rect 40048 38291 40084 38313
rect 39956 38252 40084 38291
rect 39736 38139 39775 38191
rect 39827 38139 39865 38191
rect 39736 38098 39865 38139
rect 38967 37899 39050 37955
rect 39106 37899 39230 37955
rect 39286 37899 39619 37955
rect 38967 36155 39619 37899
rect 40215 37953 40524 38799
rect 40215 37901 40253 37953
rect 40305 37901 40433 37953
rect 40485 37901 40524 37953
rect 39736 37715 39865 37756
rect 39736 37663 39775 37715
rect 39827 37663 39865 37715
rect 39736 37332 39865 37663
rect 39736 37276 39773 37332
rect 39829 37276 39865 37332
rect 39736 37237 39865 37276
rect 39956 37563 40084 37602
rect 39956 37507 39992 37563
rect 40048 37541 40084 37563
rect 40048 37507 40085 37541
rect 39956 37500 40085 37507
rect 39956 37448 39994 37500
rect 40046 37448 40085 37500
rect 39956 37314 40085 37448
rect 39956 37262 39994 37314
rect 40046 37262 40085 37314
rect 39956 37221 40085 37262
rect 40215 37055 40524 37901
rect 40215 36999 40251 37055
rect 40307 36999 40431 37055
rect 40487 36999 40524 37055
rect 39736 36778 39865 36817
rect 39736 36722 39773 36778
rect 39829 36722 39865 36778
rect 39736 36391 39865 36722
rect 39956 36792 40085 36833
rect 39956 36740 39994 36792
rect 40046 36740 40085 36792
rect 39956 36606 40085 36740
rect 39956 36554 39994 36606
rect 40046 36554 40085 36606
rect 39956 36547 40085 36554
rect 39956 36491 39992 36547
rect 40048 36513 40085 36547
rect 40048 36491 40084 36513
rect 39956 36452 40084 36491
rect 39736 36339 39775 36391
rect 39827 36339 39865 36391
rect 39736 36298 39865 36339
rect 38967 36099 39050 36155
rect 39106 36099 39230 36155
rect 39286 36099 39619 36155
rect 38967 35976 39619 36099
rect 40215 36153 40524 36999
rect 40215 36101 40253 36153
rect 40305 36101 40433 36153
rect 40485 36101 40524 36153
rect 40215 35976 40524 36101
rect 40718 35976 40939 64826
rect 41095 35976 41317 64826
rect 41473 36096 41695 65091
rect 41851 64954 42072 65091
rect 41851 64898 41881 64954
rect 42041 64898 42072 64954
rect 41851 64715 42072 64898
rect 41851 64663 41935 64715
rect 41987 64663 42072 64715
rect 41851 63391 42072 64663
rect 41851 63339 41935 63391
rect 41987 63339 42072 63391
rect 41851 62915 42072 63339
rect 41851 62863 41935 62915
rect 41987 62863 42072 62915
rect 41851 61591 42072 62863
rect 41851 61539 41935 61591
rect 41987 61539 42072 61591
rect 41851 61115 42072 61539
rect 41851 61063 41935 61115
rect 41987 61063 42072 61115
rect 41851 59791 42072 61063
rect 41851 59739 41935 59791
rect 41987 59739 42072 59791
rect 41851 59315 42072 59739
rect 41851 59263 41935 59315
rect 41987 59263 42072 59315
rect 41851 57991 42072 59263
rect 41851 57939 41935 57991
rect 41987 57939 42072 57991
rect 41851 57515 42072 57939
rect 41851 57463 41935 57515
rect 41987 57463 42072 57515
rect 41851 56191 42072 57463
rect 41851 56139 41935 56191
rect 41987 56139 42072 56191
rect 41851 55715 42072 56139
rect 41851 55663 41935 55715
rect 41987 55663 42072 55715
rect 41851 54391 42072 55663
rect 41851 54339 41935 54391
rect 41987 54339 42072 54391
rect 41851 53915 42072 54339
rect 41851 53863 41935 53915
rect 41987 53863 42072 53915
rect 41851 52591 42072 53863
rect 41851 52539 41935 52591
rect 41987 52539 42072 52591
rect 41851 52115 42072 52539
rect 41851 52063 41935 52115
rect 41987 52063 42072 52115
rect 41851 50791 42072 52063
rect 41851 50739 41935 50791
rect 41987 50739 42072 50791
rect 41851 50315 42072 50739
rect 41851 50263 41935 50315
rect 41987 50263 42072 50315
rect 41851 48991 42072 50263
rect 41851 48939 41935 48991
rect 41987 48939 42072 48991
rect 41851 48515 42072 48939
rect 41851 48463 41935 48515
rect 41987 48463 42072 48515
rect 41851 47191 42072 48463
rect 41851 47139 41935 47191
rect 41987 47139 42072 47191
rect 41851 46715 42072 47139
rect 41851 46663 41935 46715
rect 41987 46663 42072 46715
rect 41851 45391 42072 46663
rect 41851 45339 41935 45391
rect 41987 45339 42072 45391
rect 41851 44915 42072 45339
rect 41851 44863 41935 44915
rect 41987 44863 42072 44915
rect 41851 43591 42072 44863
rect 41851 43539 41935 43591
rect 41987 43539 42072 43591
rect 41851 43115 42072 43539
rect 41851 43063 41935 43115
rect 41987 43063 42072 43115
rect 41851 41791 42072 43063
rect 41851 41739 41935 41791
rect 41987 41739 42072 41791
rect 41851 41315 42072 41739
rect 41851 41263 41935 41315
rect 41987 41263 42072 41315
rect 41851 39991 42072 41263
rect 41851 39939 41935 39991
rect 41987 39939 42072 39991
rect 41851 39515 42072 39939
rect 41851 39463 41935 39515
rect 41987 39463 42072 39515
rect 41851 38191 42072 39463
rect 41851 38139 41935 38191
rect 41987 38139 42072 38191
rect 41851 37715 42072 38139
rect 41851 37663 41935 37715
rect 41987 37663 42072 37715
rect 41851 36391 42072 37663
rect 41851 36339 41935 36391
rect 41987 36339 42072 36391
rect 41851 36096 42072 36339
rect 42229 64484 42450 65091
rect 42229 64432 42312 64484
rect 42364 64432 42450 64484
rect 42229 63622 42450 64432
rect 42229 63570 42312 63622
rect 42364 63570 42450 63622
rect 42229 62684 42450 63570
rect 42229 62632 42312 62684
rect 42364 62632 42450 62684
rect 42229 61822 42450 62632
rect 42229 61770 42312 61822
rect 42364 61770 42450 61822
rect 42229 60884 42450 61770
rect 42229 60832 42312 60884
rect 42364 60832 42450 60884
rect 42229 60022 42450 60832
rect 42229 59970 42312 60022
rect 42364 59970 42450 60022
rect 42229 59084 42450 59970
rect 42229 59032 42312 59084
rect 42364 59032 42450 59084
rect 42229 58222 42450 59032
rect 42229 58170 42312 58222
rect 42364 58170 42450 58222
rect 42229 36096 42450 58170
rect 36863 35881 37743 35976
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 36863 35786 37743 35825
rect 41472 35963 41695 36096
rect 41472 35761 41694 35963
rect 41850 35778 42072 36096
rect 42228 35963 42450 36096
rect 42606 57284 42828 65091
rect 42606 57232 42690 57284
rect 42742 57232 42828 57284
rect 42606 56422 42828 57232
rect 42606 56370 42690 56422
rect 42742 56370 42828 56422
rect 42606 55484 42828 56370
rect 42606 55432 42690 55484
rect 42742 55432 42828 55484
rect 42606 54622 42828 55432
rect 42606 54570 42690 54622
rect 42742 54570 42828 54622
rect 42606 53684 42828 54570
rect 42606 53632 42690 53684
rect 42742 53632 42828 53684
rect 42606 52822 42828 53632
rect 42606 52770 42690 52822
rect 42742 52770 42828 52822
rect 42606 51884 42828 52770
rect 42606 51832 42690 51884
rect 42742 51832 42828 51884
rect 42606 51022 42828 51832
rect 42606 50970 42690 51022
rect 42742 50970 42828 51022
rect 42606 36085 42828 50970
rect 42984 50084 43205 65091
rect 42984 50032 43068 50084
rect 43120 50032 43205 50084
rect 42984 49222 43205 50032
rect 42984 49170 43068 49222
rect 43120 49170 43205 49222
rect 42984 48284 43205 49170
rect 42984 48232 43068 48284
rect 43120 48232 43205 48284
rect 42984 47422 43205 48232
rect 42984 47370 43068 47422
rect 43120 47370 43205 47422
rect 42984 46484 43205 47370
rect 42984 46432 43068 46484
rect 43120 46432 43205 46484
rect 42984 45622 43205 46432
rect 42984 45570 43068 45622
rect 43120 45570 43205 45622
rect 42984 44684 43205 45570
rect 42984 44632 43068 44684
rect 43120 44632 43205 44684
rect 42984 43822 43205 44632
rect 42984 43770 43068 43822
rect 43120 43770 43205 43822
rect 42984 36096 43205 43770
rect 42603 35963 42828 36085
rect 38596 35532 41694 35761
rect 38596 35516 38817 35532
rect 27387 34968 27478 35024
rect 27534 34968 27690 35024
rect 27746 34968 27828 35024
rect 27387 34960 27828 34968
rect 27387 34596 27469 34960
rect 27729 34806 27828 34960
rect 27746 34750 27828 34806
rect 27729 34596 27828 34750
rect 27387 34588 27828 34596
rect 27387 34532 27478 34588
rect 27534 34532 27690 34588
rect 27746 34532 27828 34588
rect 27387 33432 27828 34532
rect 27387 33380 27476 33432
rect 27528 33380 27688 33432
rect 27740 33380 27828 33432
rect 27387 33215 27828 33380
rect 31615 35287 38817 35516
rect 41850 35425 42072 35509
rect 31615 33349 31836 35287
rect 39077 35197 42072 35425
rect 39077 35171 39298 35197
rect 31970 34943 39298 35171
rect 42228 35090 42449 35963
rect 31970 33349 32192 34943
rect 39755 34861 42449 35090
rect 39755 34675 39977 34861
rect 42603 34754 42825 35963
rect 38301 34491 39977 34675
rect 37201 34446 39977 34491
rect 40106 34526 42825 34754
rect 37201 34263 38523 34446
rect 40106 34312 40328 34526
rect 42983 34419 43205 36096
rect 43362 42884 43583 65091
rect 43703 64953 44564 65853
rect 48789 65833 49990 66376
rect 48789 65781 48828 65833
rect 48880 65781 49039 65833
rect 49091 65781 49250 65833
rect 49302 65781 49461 65833
rect 49513 65781 49990 65833
rect 48789 65370 49990 65781
rect 48789 65318 48828 65370
rect 48880 65318 49039 65370
rect 49091 65318 49250 65370
rect 49302 65318 49461 65370
rect 49513 65318 49990 65370
rect 43703 64940 43790 64953
rect 43362 42832 43445 42884
rect 43497 42832 43583 42884
rect 43362 42022 43583 42832
rect 43362 41970 43445 42022
rect 43497 41970 43583 42022
rect 43362 41084 43583 41970
rect 43362 41032 43445 41084
rect 43497 41032 43583 41084
rect 43362 40222 43583 41032
rect 43362 40170 43445 40222
rect 43497 40170 43583 40222
rect 43362 39284 43583 40170
rect 43362 39232 43445 39284
rect 43497 39232 43583 39284
rect 43362 38422 43583 39232
rect 43362 38370 43445 38422
rect 43497 38370 43583 38422
rect 43362 37484 43583 38370
rect 43362 37432 43445 37484
rect 43497 37432 43583 37484
rect 43362 36622 43583 37432
rect 43362 36570 43445 36622
rect 43497 36570 43583 36622
rect 43362 36085 43583 36570
rect 37201 33360 37423 34263
rect 38642 34156 40328 34312
rect 37557 34084 40328 34156
rect 40458 34190 43205 34419
rect 43359 35963 43583 36085
rect 43704 64901 43790 64940
rect 43842 64901 44001 64953
rect 44053 64901 44213 64953
rect 44265 64901 44424 64953
rect 44476 64940 44564 64953
rect 44758 64955 45384 65078
rect 44476 64901 44563 64940
rect 43704 64055 44563 64901
rect 43704 63999 43788 64055
rect 43844 63999 43999 64055
rect 44055 63999 44211 64055
rect 44267 63999 44422 64055
rect 44478 63999 44563 64055
rect 43704 63153 44563 63999
rect 43704 63101 43790 63153
rect 43842 63101 44001 63153
rect 44053 63101 44213 63153
rect 44265 63101 44424 63153
rect 44476 63101 44563 63153
rect 43704 62255 44563 63101
rect 43704 62199 43788 62255
rect 43844 62199 43999 62255
rect 44055 62199 44211 62255
rect 44267 62199 44422 62255
rect 44478 62199 44563 62255
rect 43704 61353 44563 62199
rect 43704 61301 43790 61353
rect 43842 61301 44001 61353
rect 44053 61301 44213 61353
rect 44265 61301 44424 61353
rect 44476 61301 44563 61353
rect 43704 60455 44563 61301
rect 43704 60399 43788 60455
rect 43844 60399 43999 60455
rect 44055 60399 44211 60455
rect 44267 60399 44422 60455
rect 44478 60399 44563 60455
rect 43704 59553 44563 60399
rect 43704 59501 43790 59553
rect 43842 59501 44001 59553
rect 44053 59501 44213 59553
rect 44265 59501 44424 59553
rect 44476 59501 44563 59553
rect 43704 58655 44563 59501
rect 43704 58599 43788 58655
rect 43844 58599 43999 58655
rect 44055 58599 44211 58655
rect 44267 58599 44422 58655
rect 44478 58599 44563 58655
rect 43704 57753 44563 58599
rect 43704 57701 43790 57753
rect 43842 57701 44001 57753
rect 44053 57701 44213 57753
rect 44265 57701 44424 57753
rect 44476 57701 44563 57753
rect 43704 56855 44563 57701
rect 43704 56799 43788 56855
rect 43844 56799 43999 56855
rect 44055 56799 44211 56855
rect 44267 56799 44422 56855
rect 44478 56799 44563 56855
rect 43704 55953 44563 56799
rect 43704 55901 43790 55953
rect 43842 55901 44001 55953
rect 44053 55901 44213 55953
rect 44265 55901 44424 55953
rect 44476 55901 44563 55953
rect 43704 55055 44563 55901
rect 43704 54999 43788 55055
rect 43844 54999 43999 55055
rect 44055 54999 44211 55055
rect 44267 54999 44422 55055
rect 44478 54999 44563 55055
rect 43704 54153 44563 54999
rect 43704 54101 43790 54153
rect 43842 54101 44001 54153
rect 44053 54101 44213 54153
rect 44265 54101 44424 54153
rect 44476 54101 44563 54153
rect 43704 53255 44563 54101
rect 43704 53199 43788 53255
rect 43844 53199 43999 53255
rect 44055 53199 44211 53255
rect 44267 53199 44422 53255
rect 44478 53199 44563 53255
rect 43704 52353 44563 53199
rect 43704 52301 43790 52353
rect 43842 52301 44001 52353
rect 44053 52301 44213 52353
rect 44265 52301 44424 52353
rect 44476 52301 44563 52353
rect 43704 51455 44563 52301
rect 43704 51399 43788 51455
rect 43844 51399 43999 51455
rect 44055 51399 44211 51455
rect 44267 51399 44422 51455
rect 44478 51399 44563 51455
rect 43704 50553 44563 51399
rect 43704 50501 43790 50553
rect 43842 50501 44001 50553
rect 44053 50501 44213 50553
rect 44265 50501 44424 50553
rect 44476 50501 44563 50553
rect 43704 49655 44563 50501
rect 43704 49599 43788 49655
rect 43844 49599 43999 49655
rect 44055 49599 44211 49655
rect 44267 49599 44422 49655
rect 44478 49599 44563 49655
rect 43704 48753 44563 49599
rect 43704 48701 43790 48753
rect 43842 48701 44001 48753
rect 44053 48701 44213 48753
rect 44265 48701 44424 48753
rect 44476 48701 44563 48753
rect 43704 47855 44563 48701
rect 43704 47799 43788 47855
rect 43844 47799 43999 47855
rect 44055 47799 44211 47855
rect 44267 47799 44422 47855
rect 44478 47799 44563 47855
rect 43704 46953 44563 47799
rect 43704 46901 43790 46953
rect 43842 46901 44001 46953
rect 44053 46901 44213 46953
rect 44265 46901 44424 46953
rect 44476 46901 44563 46953
rect 43704 46055 44563 46901
rect 43704 45999 43788 46055
rect 43844 45999 43999 46055
rect 44055 45999 44211 46055
rect 44267 45999 44422 46055
rect 44478 45999 44563 46055
rect 43704 45153 44563 45999
rect 43704 45101 43790 45153
rect 43842 45101 44001 45153
rect 44053 45101 44213 45153
rect 44265 45101 44424 45153
rect 44476 45101 44563 45153
rect 43704 44255 44563 45101
rect 43704 44199 43788 44255
rect 43844 44199 43999 44255
rect 44055 44199 44211 44255
rect 44267 44199 44422 44255
rect 44478 44199 44563 44255
rect 43704 43353 44563 44199
rect 43704 43301 43790 43353
rect 43842 43301 44001 43353
rect 44053 43301 44213 43353
rect 44265 43301 44424 43353
rect 44476 43301 44563 43353
rect 43704 42455 44563 43301
rect 43704 42399 43788 42455
rect 43844 42399 43999 42455
rect 44055 42399 44211 42455
rect 44267 42399 44422 42455
rect 44478 42399 44563 42455
rect 43704 41553 44563 42399
rect 43704 41501 43790 41553
rect 43842 41501 44001 41553
rect 44053 41501 44213 41553
rect 44265 41501 44424 41553
rect 44476 41501 44563 41553
rect 43704 40655 44563 41501
rect 43704 40599 43788 40655
rect 43844 40599 43999 40655
rect 44055 40599 44211 40655
rect 44267 40599 44422 40655
rect 44478 40599 44563 40655
rect 43704 39753 44563 40599
rect 43704 39701 43790 39753
rect 43842 39701 44001 39753
rect 44053 39701 44213 39753
rect 44265 39701 44424 39753
rect 44476 39701 44563 39753
rect 43704 38855 44563 39701
rect 43704 38799 43788 38855
rect 43844 38799 43999 38855
rect 44055 38799 44211 38855
rect 44267 38799 44422 38855
rect 44478 38799 44563 38855
rect 43704 37953 44563 38799
rect 43704 37901 43790 37953
rect 43842 37901 44001 37953
rect 44053 37901 44213 37953
rect 44265 37901 44424 37953
rect 44476 37901 44563 37953
rect 43704 37055 44563 37901
rect 43704 36999 43788 37055
rect 43844 36999 43999 37055
rect 44055 36999 44211 37055
rect 44267 36999 44422 37055
rect 44478 36999 44563 37055
rect 43704 36153 44563 36999
rect 43704 36101 43790 36153
rect 43842 36101 44001 36153
rect 44053 36101 44213 36153
rect 44265 36101 44424 36153
rect 44476 36101 44563 36153
rect 43704 35976 44563 36101
rect 44758 64899 44832 64955
rect 44888 64899 45043 64955
rect 45099 64899 45254 64955
rect 45310 64899 45384 64955
rect 44758 64491 45384 64899
rect 44758 64439 44939 64491
rect 44991 64439 45151 64491
rect 45203 64439 45384 64491
rect 44758 63615 45384 64439
rect 44758 63563 44939 63615
rect 44991 63563 45151 63615
rect 45203 63563 45384 63615
rect 44758 63155 45384 63563
rect 44758 63099 44832 63155
rect 44888 63099 45043 63155
rect 45099 63099 45254 63155
rect 45310 63099 45384 63155
rect 44758 62691 45384 63099
rect 44758 62639 44939 62691
rect 44991 62639 45151 62691
rect 45203 62639 45384 62691
rect 44758 61815 45384 62639
rect 44758 61763 44939 61815
rect 44991 61763 45151 61815
rect 45203 61763 45384 61815
rect 44758 61355 45384 61763
rect 44758 61299 44832 61355
rect 44888 61299 45043 61355
rect 45099 61299 45254 61355
rect 45310 61299 45384 61355
rect 44758 60891 45384 61299
rect 44758 60839 44939 60891
rect 44991 60839 45151 60891
rect 45203 60839 45384 60891
rect 44758 60015 45384 60839
rect 44758 59963 44939 60015
rect 44991 59963 45151 60015
rect 45203 59963 45384 60015
rect 44758 59555 45384 59963
rect 44758 59499 44832 59555
rect 44888 59499 45043 59555
rect 45099 59499 45254 59555
rect 45310 59499 45384 59555
rect 44758 59091 45384 59499
rect 44758 59039 44939 59091
rect 44991 59039 45151 59091
rect 45203 59039 45384 59091
rect 44758 58215 45384 59039
rect 44758 58163 44939 58215
rect 44991 58163 45151 58215
rect 45203 58163 45384 58215
rect 44758 57755 45384 58163
rect 44758 57699 44832 57755
rect 44888 57699 45043 57755
rect 45099 57699 45254 57755
rect 45310 57699 45384 57755
rect 44758 57291 45384 57699
rect 44758 57239 44939 57291
rect 44991 57239 45151 57291
rect 45203 57239 45384 57291
rect 44758 56415 45384 57239
rect 44758 56363 44939 56415
rect 44991 56363 45151 56415
rect 45203 56363 45384 56415
rect 44758 55955 45384 56363
rect 44758 55899 44832 55955
rect 44888 55899 45043 55955
rect 45099 55899 45254 55955
rect 45310 55899 45384 55955
rect 44758 55491 45384 55899
rect 44758 55439 44939 55491
rect 44991 55439 45151 55491
rect 45203 55439 45384 55491
rect 44758 54615 45384 55439
rect 44758 54563 44939 54615
rect 44991 54563 45151 54615
rect 45203 54563 45384 54615
rect 44758 54155 45384 54563
rect 44758 54099 44832 54155
rect 44888 54099 45043 54155
rect 45099 54099 45254 54155
rect 45310 54099 45384 54155
rect 44758 53691 45384 54099
rect 44758 53639 44939 53691
rect 44991 53639 45151 53691
rect 45203 53639 45384 53691
rect 44758 52815 45384 53639
rect 44758 52763 44939 52815
rect 44991 52763 45151 52815
rect 45203 52763 45384 52815
rect 44758 52355 45384 52763
rect 44758 52299 44832 52355
rect 44888 52299 45043 52355
rect 45099 52299 45254 52355
rect 45310 52299 45384 52355
rect 44758 51891 45384 52299
rect 44758 51839 44939 51891
rect 44991 51839 45151 51891
rect 45203 51839 45384 51891
rect 44758 51015 45384 51839
rect 44758 50963 44939 51015
rect 44991 50963 45151 51015
rect 45203 50963 45384 51015
rect 44758 50555 45384 50963
rect 44758 50499 44832 50555
rect 44888 50499 45043 50555
rect 45099 50499 45254 50555
rect 45310 50499 45384 50555
rect 44758 50091 45384 50499
rect 44758 50039 44939 50091
rect 44991 50039 45151 50091
rect 45203 50039 45384 50091
rect 44758 49215 45384 50039
rect 44758 49163 44939 49215
rect 44991 49163 45151 49215
rect 45203 49163 45384 49215
rect 44758 48755 45384 49163
rect 44758 48699 44832 48755
rect 44888 48699 45043 48755
rect 45099 48699 45254 48755
rect 45310 48699 45384 48755
rect 44758 48291 45384 48699
rect 44758 48239 44939 48291
rect 44991 48239 45151 48291
rect 45203 48239 45384 48291
rect 44758 47415 45384 48239
rect 44758 47363 44939 47415
rect 44991 47363 45151 47415
rect 45203 47363 45384 47415
rect 44758 46955 45384 47363
rect 44758 46899 44832 46955
rect 44888 46899 45043 46955
rect 45099 46899 45254 46955
rect 45310 46899 45384 46955
rect 44758 46491 45384 46899
rect 44758 46439 44939 46491
rect 44991 46439 45151 46491
rect 45203 46439 45384 46491
rect 44758 45615 45384 46439
rect 44758 45563 44939 45615
rect 44991 45563 45151 45615
rect 45203 45563 45384 45615
rect 44758 45155 45384 45563
rect 44758 45099 44832 45155
rect 44888 45099 45043 45155
rect 45099 45099 45254 45155
rect 45310 45099 45384 45155
rect 44758 44691 45384 45099
rect 44758 44639 44939 44691
rect 44991 44639 45151 44691
rect 45203 44639 45384 44691
rect 44758 43815 45384 44639
rect 44758 43763 44939 43815
rect 44991 43763 45151 43815
rect 45203 43763 45384 43815
rect 44758 43355 45384 43763
rect 44758 43299 44832 43355
rect 44888 43299 45043 43355
rect 45099 43299 45254 43355
rect 45310 43299 45384 43355
rect 44758 42891 45384 43299
rect 44758 42839 44939 42891
rect 44991 42839 45151 42891
rect 45203 42839 45384 42891
rect 44758 42015 45384 42839
rect 44758 41963 44939 42015
rect 44991 41963 45151 42015
rect 45203 41963 45384 42015
rect 44758 41555 45384 41963
rect 44758 41499 44832 41555
rect 44888 41499 45043 41555
rect 45099 41499 45254 41555
rect 45310 41499 45384 41555
rect 44758 41091 45384 41499
rect 44758 41039 44939 41091
rect 44991 41039 45151 41091
rect 45203 41039 45384 41091
rect 44758 40215 45384 41039
rect 44758 40163 44939 40215
rect 44991 40163 45151 40215
rect 45203 40163 45384 40215
rect 44758 39755 45384 40163
rect 44758 39699 44832 39755
rect 44888 39699 45043 39755
rect 45099 39699 45254 39755
rect 45310 39699 45384 39755
rect 44758 39291 45384 39699
rect 44758 39239 44939 39291
rect 44991 39239 45151 39291
rect 45203 39239 45384 39291
rect 44758 38415 45384 39239
rect 44758 38363 44939 38415
rect 44991 38363 45151 38415
rect 45203 38363 45384 38415
rect 44758 37955 45384 38363
rect 44758 37899 44832 37955
rect 44888 37899 45043 37955
rect 45099 37899 45254 37955
rect 45310 37899 45384 37955
rect 44758 37491 45384 37899
rect 44758 37439 44939 37491
rect 44991 37439 45151 37491
rect 45203 37439 45384 37491
rect 44758 36615 45384 37439
rect 44758 36563 44939 36615
rect 44991 36563 45151 36615
rect 45203 36563 45384 36615
rect 44758 36155 45384 36563
rect 44758 36099 44832 36155
rect 44888 36099 45043 36155
rect 45099 36099 45254 36155
rect 45310 36099 45384 36155
rect 44758 35976 45384 36099
rect 45514 64375 45735 65091
rect 45514 64323 45597 64375
rect 45649 64323 45735 64375
rect 45514 57175 45735 64323
rect 45514 57123 45597 57175
rect 45649 57123 45735 57175
rect 45514 49975 45735 57123
rect 45514 49923 45597 49975
rect 45649 49923 45735 49975
rect 45514 42775 45735 49923
rect 45514 42723 45597 42775
rect 45649 42723 45735 42775
rect 45514 36096 45735 42723
rect 37557 33927 38863 34084
rect 40458 33977 40679 34190
rect 43359 34083 43580 35963
rect 45513 35842 45735 36096
rect 37557 33349 37778 33927
rect 38993 33748 40679 33977
rect 40809 33855 43580 34083
rect 44646 35614 45735 35842
rect 45891 63731 46113 65091
rect 45891 63679 45975 63731
rect 46027 63679 46113 63731
rect 45891 56531 46113 63679
rect 45891 56479 45975 56531
rect 46027 56479 46113 56531
rect 45891 49331 46113 56479
rect 45891 49279 45975 49331
rect 46027 49279 46113 49331
rect 45891 42131 46113 49279
rect 45891 42079 45975 42131
rect 46027 42079 46113 42131
rect 45891 35963 46113 42079
rect 46269 62575 46491 65091
rect 46269 62523 46353 62575
rect 46405 62523 46491 62575
rect 46269 55375 46491 62523
rect 46269 55323 46353 55375
rect 46405 55323 46491 55375
rect 46269 48175 46491 55323
rect 46269 48123 46353 48175
rect 46405 48123 46491 48175
rect 46269 40975 46491 48123
rect 46269 40923 46353 40975
rect 46405 40923 46491 40975
rect 46269 36096 46491 40923
rect 46268 35963 46491 36096
rect 46647 61931 46868 65091
rect 46647 61879 46731 61931
rect 46783 61879 46868 61931
rect 46647 54731 46868 61879
rect 46647 54679 46731 54731
rect 46783 54679 46868 54731
rect 46647 47531 46868 54679
rect 46647 47479 46731 47531
rect 46783 47479 46868 47531
rect 46647 40331 46868 47479
rect 46647 40279 46731 40331
rect 46783 40279 46868 40331
rect 46647 36085 46868 40279
rect 38993 33360 39215 33748
rect 40809 33625 41031 33855
rect 39349 33397 41031 33625
rect 44646 33576 44867 35614
rect 45891 35507 46112 35963
rect 44997 35278 46112 35507
rect 46268 35681 46490 35963
rect 46268 35453 46501 35681
rect 44997 33576 45219 35278
rect 46279 33576 46501 35453
rect 46646 35346 46868 36085
rect 47025 60775 47246 65091
rect 47025 60723 47108 60775
rect 47160 60723 47246 60775
rect 47025 53575 47246 60723
rect 47025 53523 47108 53575
rect 47160 53523 47246 53575
rect 47025 46375 47246 53523
rect 47025 46323 47108 46375
rect 47160 46323 47246 46375
rect 47025 39175 47246 46323
rect 47025 39123 47108 39175
rect 47160 39123 47246 39175
rect 47025 36085 47246 39123
rect 47402 60131 47624 65091
rect 47402 60079 47486 60131
rect 47538 60079 47624 60131
rect 47402 52931 47624 60079
rect 47402 52879 47486 52931
rect 47538 52879 47624 52931
rect 47402 45731 47624 52879
rect 47402 45679 47486 45731
rect 47538 45679 47624 45731
rect 47402 38531 47624 45679
rect 47402 38479 47486 38531
rect 47538 38479 47624 38531
rect 47025 35963 47248 36085
rect 46631 35117 46868 35346
rect 46631 33564 46852 35117
rect 47026 34836 47248 35963
rect 47402 35963 47624 38479
rect 47780 58975 48002 65091
rect 47780 58923 47864 58975
rect 47916 58923 48002 58975
rect 47780 51775 48002 58923
rect 47780 51723 47864 51775
rect 47916 51723 48002 51775
rect 47780 44575 48002 51723
rect 47780 44523 47864 44575
rect 47916 44523 48002 44575
rect 47780 37375 48002 44523
rect 47780 37323 47864 37375
rect 47916 37323 48002 37375
rect 47780 36096 48002 37323
rect 48158 58331 48379 65091
rect 48789 65078 49990 65318
rect 50098 65855 50913 65946
rect 50098 65799 50135 65855
rect 50191 65799 50346 65855
rect 50402 65799 50557 65855
rect 50613 65799 50768 65855
rect 50824 65799 50913 65855
rect 50098 65635 50913 65799
rect 50098 65583 50137 65635
rect 50189 65583 50348 65635
rect 50400 65583 50559 65635
rect 50611 65583 50770 65635
rect 50822 65583 50913 65635
rect 48789 64955 49991 65078
rect 48789 64940 48836 64955
rect 48790 64899 48836 64940
rect 48892 64899 49046 64955
rect 49102 64899 49257 64955
rect 49313 64899 49469 64955
rect 49525 64899 49680 64955
rect 49736 64899 49890 64955
rect 49946 64899 49991 64955
rect 50098 64953 50913 65583
rect 52226 65853 54354 66376
rect 52226 65801 52576 65853
rect 52628 65801 52787 65853
rect 52839 65801 52998 65853
rect 53050 65801 53209 65853
rect 53261 65801 53419 65853
rect 53471 65801 53630 65853
rect 53682 65801 53841 65853
rect 53893 65801 54052 65853
rect 54104 65801 54263 65853
rect 54315 65801 54354 65853
rect 52226 65635 54354 65801
rect 52226 65583 52576 65635
rect 52628 65583 52787 65635
rect 52839 65583 52998 65635
rect 53050 65583 53209 65635
rect 53261 65583 53419 65635
rect 53471 65583 53630 65635
rect 53682 65583 53841 65635
rect 53893 65583 54052 65635
rect 54104 65583 54263 65635
rect 54315 65583 54354 65635
rect 52226 65418 54354 65583
rect 51042 65372 52015 65411
rect 51042 65316 51079 65372
rect 51135 65316 51290 65372
rect 51346 65316 51501 65372
rect 51557 65316 51712 65372
rect 51768 65316 51923 65372
rect 51979 65316 52015 65372
rect 51042 65278 52015 65316
rect 52226 65366 52576 65418
rect 52628 65366 52787 65418
rect 52839 65366 52998 65418
rect 53050 65366 53209 65418
rect 53261 65366 53419 65418
rect 53471 65366 53630 65418
rect 53682 65366 53841 65418
rect 53893 65366 54052 65418
rect 54104 65366 54263 65418
rect 54315 65366 54354 65418
rect 50098 64940 50346 64953
rect 48790 64654 49991 64899
rect 48790 64602 48943 64654
rect 48995 64602 49154 64654
rect 49206 64602 49365 64654
rect 49417 64602 49576 64654
rect 49628 64602 49787 64654
rect 49839 64602 49991 64654
rect 48557 64549 48687 64588
rect 48557 64493 48594 64549
rect 48650 64493 48687 64549
rect 48557 64331 48687 64493
rect 48557 64275 48594 64331
rect 48650 64275 48687 64331
rect 48557 64237 48687 64275
rect 48790 64191 49991 64602
rect 48790 64139 48943 64191
rect 48995 64139 49154 64191
rect 49206 64139 49365 64191
rect 49417 64139 49576 64191
rect 49628 64139 49787 64191
rect 49839 64139 49991 64191
rect 48790 63915 49991 64139
rect 48790 63863 48943 63915
rect 48995 63863 49154 63915
rect 49206 63863 49365 63915
rect 49417 63863 49576 63915
rect 49628 63863 49787 63915
rect 49839 63863 49991 63915
rect 48557 63779 48687 63817
rect 48557 63723 48594 63779
rect 48650 63723 48687 63779
rect 48557 63561 48687 63723
rect 48557 63505 48594 63561
rect 48650 63505 48687 63561
rect 48557 63466 48687 63505
rect 48790 63452 49991 63863
rect 48790 63400 48943 63452
rect 48995 63400 49154 63452
rect 49206 63400 49365 63452
rect 49417 63400 49576 63452
rect 49628 63400 49787 63452
rect 49839 63400 49991 63452
rect 48790 63155 49991 63400
rect 48790 63099 48836 63155
rect 48892 63099 49046 63155
rect 49102 63099 49257 63155
rect 49313 63099 49469 63155
rect 49525 63099 49680 63155
rect 49736 63099 49890 63155
rect 49946 63099 49991 63155
rect 48790 62854 49991 63099
rect 48790 62802 48943 62854
rect 48995 62802 49154 62854
rect 49206 62802 49365 62854
rect 49417 62802 49576 62854
rect 49628 62802 49787 62854
rect 49839 62802 49991 62854
rect 48557 62749 48687 62788
rect 48557 62693 48594 62749
rect 48650 62693 48687 62749
rect 48557 62531 48687 62693
rect 48557 62475 48594 62531
rect 48650 62475 48687 62531
rect 48557 62437 48687 62475
rect 48790 62391 49991 62802
rect 48790 62339 48943 62391
rect 48995 62339 49154 62391
rect 49206 62339 49365 62391
rect 49417 62339 49576 62391
rect 49628 62339 49787 62391
rect 49839 62339 49991 62391
rect 48790 62115 49991 62339
rect 48790 62063 48943 62115
rect 48995 62063 49154 62115
rect 49206 62063 49365 62115
rect 49417 62063 49576 62115
rect 49628 62063 49787 62115
rect 49839 62063 49991 62115
rect 48557 61979 48687 62017
rect 48557 61923 48594 61979
rect 48650 61923 48687 61979
rect 48557 61761 48687 61923
rect 48557 61705 48594 61761
rect 48650 61705 48687 61761
rect 48557 61666 48687 61705
rect 48790 61652 49991 62063
rect 48790 61600 48943 61652
rect 48995 61600 49154 61652
rect 49206 61600 49365 61652
rect 49417 61600 49576 61652
rect 49628 61600 49787 61652
rect 49839 61600 49991 61652
rect 48790 61355 49991 61600
rect 48790 61299 48836 61355
rect 48892 61299 49046 61355
rect 49102 61299 49257 61355
rect 49313 61299 49469 61355
rect 49525 61299 49680 61355
rect 49736 61299 49890 61355
rect 49946 61299 49991 61355
rect 48790 61054 49991 61299
rect 48790 61002 48943 61054
rect 48995 61002 49154 61054
rect 49206 61002 49365 61054
rect 49417 61002 49576 61054
rect 49628 61002 49787 61054
rect 49839 61002 49991 61054
rect 48557 60949 48687 60988
rect 48557 60893 48594 60949
rect 48650 60893 48687 60949
rect 48557 60731 48687 60893
rect 48557 60675 48594 60731
rect 48650 60675 48687 60731
rect 48557 60637 48687 60675
rect 48790 60591 49991 61002
rect 48790 60539 48943 60591
rect 48995 60539 49154 60591
rect 49206 60539 49365 60591
rect 49417 60539 49576 60591
rect 49628 60539 49787 60591
rect 49839 60539 49991 60591
rect 48790 60315 49991 60539
rect 48790 60263 48943 60315
rect 48995 60263 49154 60315
rect 49206 60263 49365 60315
rect 49417 60263 49576 60315
rect 49628 60263 49787 60315
rect 49839 60263 49991 60315
rect 48557 60179 48687 60217
rect 48557 60123 48594 60179
rect 48650 60123 48687 60179
rect 48557 59961 48687 60123
rect 48557 59905 48594 59961
rect 48650 59905 48687 59961
rect 48557 59866 48687 59905
rect 48790 59852 49991 60263
rect 48790 59800 48943 59852
rect 48995 59800 49154 59852
rect 49206 59800 49365 59852
rect 49417 59800 49576 59852
rect 49628 59800 49787 59852
rect 49839 59800 49991 59852
rect 48790 59555 49991 59800
rect 48790 59499 48836 59555
rect 48892 59499 49046 59555
rect 49102 59499 49257 59555
rect 49313 59499 49469 59555
rect 49525 59499 49680 59555
rect 49736 59499 49890 59555
rect 49946 59499 49991 59555
rect 48790 59254 49991 59499
rect 48790 59202 48943 59254
rect 48995 59202 49154 59254
rect 49206 59202 49365 59254
rect 49417 59202 49576 59254
rect 49628 59202 49787 59254
rect 49839 59202 49991 59254
rect 48557 59149 48687 59188
rect 48557 59093 48594 59149
rect 48650 59093 48687 59149
rect 48557 58931 48687 59093
rect 48557 58875 48594 58931
rect 48650 58875 48687 58931
rect 48557 58837 48687 58875
rect 48790 58791 49991 59202
rect 48790 58739 48943 58791
rect 48995 58739 49154 58791
rect 49206 58739 49365 58791
rect 49417 58739 49576 58791
rect 49628 58739 49787 58791
rect 49839 58739 49991 58791
rect 48790 58515 49991 58739
rect 48790 58463 48943 58515
rect 48995 58463 49154 58515
rect 49206 58463 49365 58515
rect 49417 58463 49576 58515
rect 49628 58463 49787 58515
rect 49839 58463 49991 58515
rect 48158 58279 48241 58331
rect 48293 58279 48379 58331
rect 48158 51131 48379 58279
rect 48557 58379 48687 58417
rect 48557 58323 48594 58379
rect 48650 58323 48687 58379
rect 48557 58161 48687 58323
rect 48557 58105 48594 58161
rect 48650 58105 48687 58161
rect 48557 58066 48687 58105
rect 48790 58052 49991 58463
rect 48790 58000 48943 58052
rect 48995 58000 49154 58052
rect 49206 58000 49365 58052
rect 49417 58000 49576 58052
rect 49628 58000 49787 58052
rect 49839 58000 49991 58052
rect 48790 57755 49991 58000
rect 48790 57699 48836 57755
rect 48892 57699 49046 57755
rect 49102 57699 49257 57755
rect 49313 57699 49469 57755
rect 49525 57699 49680 57755
rect 49736 57699 49890 57755
rect 49946 57699 49991 57755
rect 48790 57454 49991 57699
rect 48790 57402 48943 57454
rect 48995 57402 49154 57454
rect 49206 57402 49365 57454
rect 49417 57402 49576 57454
rect 49628 57402 49787 57454
rect 49839 57402 49991 57454
rect 48557 57349 48687 57388
rect 48557 57293 48594 57349
rect 48650 57293 48687 57349
rect 48557 57131 48687 57293
rect 48557 57075 48594 57131
rect 48650 57075 48687 57131
rect 48557 57037 48687 57075
rect 48790 56991 49991 57402
rect 48790 56939 48943 56991
rect 48995 56939 49154 56991
rect 49206 56939 49365 56991
rect 49417 56939 49576 56991
rect 49628 56939 49787 56991
rect 49839 56939 49991 56991
rect 48790 56715 49991 56939
rect 48790 56663 48943 56715
rect 48995 56663 49154 56715
rect 49206 56663 49365 56715
rect 49417 56663 49576 56715
rect 49628 56663 49787 56715
rect 49839 56663 49991 56715
rect 48557 56579 48687 56617
rect 48557 56523 48594 56579
rect 48650 56523 48687 56579
rect 48557 56361 48687 56523
rect 48557 56305 48594 56361
rect 48650 56305 48687 56361
rect 48557 56266 48687 56305
rect 48790 56252 49991 56663
rect 48790 56200 48943 56252
rect 48995 56200 49154 56252
rect 49206 56200 49365 56252
rect 49417 56200 49576 56252
rect 49628 56200 49787 56252
rect 49839 56200 49991 56252
rect 48790 55955 49991 56200
rect 48790 55899 48836 55955
rect 48892 55899 49046 55955
rect 49102 55899 49257 55955
rect 49313 55899 49469 55955
rect 49525 55899 49680 55955
rect 49736 55899 49890 55955
rect 49946 55899 49991 55955
rect 48790 55654 49991 55899
rect 48790 55602 48943 55654
rect 48995 55602 49154 55654
rect 49206 55602 49365 55654
rect 49417 55602 49576 55654
rect 49628 55602 49787 55654
rect 49839 55602 49991 55654
rect 48557 55549 48687 55588
rect 48557 55493 48594 55549
rect 48650 55493 48687 55549
rect 48557 55331 48687 55493
rect 48557 55275 48594 55331
rect 48650 55275 48687 55331
rect 48557 55237 48687 55275
rect 48790 55191 49991 55602
rect 48790 55139 48943 55191
rect 48995 55139 49154 55191
rect 49206 55139 49365 55191
rect 49417 55139 49576 55191
rect 49628 55139 49787 55191
rect 49839 55139 49991 55191
rect 48790 54915 49991 55139
rect 48790 54863 48943 54915
rect 48995 54863 49154 54915
rect 49206 54863 49365 54915
rect 49417 54863 49576 54915
rect 49628 54863 49787 54915
rect 49839 54863 49991 54915
rect 48557 54779 48687 54817
rect 48557 54723 48594 54779
rect 48650 54723 48687 54779
rect 48557 54561 48687 54723
rect 48557 54505 48594 54561
rect 48650 54505 48687 54561
rect 48557 54466 48687 54505
rect 48790 54452 49991 54863
rect 48790 54400 48943 54452
rect 48995 54400 49154 54452
rect 49206 54400 49365 54452
rect 49417 54400 49576 54452
rect 49628 54400 49787 54452
rect 49839 54400 49991 54452
rect 48790 54155 49991 54400
rect 48790 54099 48836 54155
rect 48892 54099 49046 54155
rect 49102 54099 49257 54155
rect 49313 54099 49469 54155
rect 49525 54099 49680 54155
rect 49736 54099 49890 54155
rect 49946 54099 49991 54155
rect 48790 53854 49991 54099
rect 48790 53802 48943 53854
rect 48995 53802 49154 53854
rect 49206 53802 49365 53854
rect 49417 53802 49576 53854
rect 49628 53802 49787 53854
rect 49839 53802 49991 53854
rect 48557 53749 48687 53788
rect 48557 53693 48594 53749
rect 48650 53693 48687 53749
rect 48557 53531 48687 53693
rect 48557 53475 48594 53531
rect 48650 53475 48687 53531
rect 48557 53437 48687 53475
rect 48790 53391 49991 53802
rect 48790 53339 48943 53391
rect 48995 53339 49154 53391
rect 49206 53339 49365 53391
rect 49417 53339 49576 53391
rect 49628 53339 49787 53391
rect 49839 53339 49991 53391
rect 48790 53115 49991 53339
rect 48790 53063 48943 53115
rect 48995 53063 49154 53115
rect 49206 53063 49365 53115
rect 49417 53063 49576 53115
rect 49628 53063 49787 53115
rect 49839 53063 49991 53115
rect 48557 52979 48687 53017
rect 48557 52923 48594 52979
rect 48650 52923 48687 52979
rect 48557 52761 48687 52923
rect 48557 52705 48594 52761
rect 48650 52705 48687 52761
rect 48557 52666 48687 52705
rect 48790 52652 49991 53063
rect 48790 52600 48943 52652
rect 48995 52600 49154 52652
rect 49206 52600 49365 52652
rect 49417 52600 49576 52652
rect 49628 52600 49787 52652
rect 49839 52600 49991 52652
rect 48790 52355 49991 52600
rect 48790 52299 48836 52355
rect 48892 52299 49046 52355
rect 49102 52299 49257 52355
rect 49313 52299 49469 52355
rect 49525 52299 49680 52355
rect 49736 52299 49890 52355
rect 49946 52299 49991 52355
rect 48790 52054 49991 52299
rect 48790 52002 48943 52054
rect 48995 52002 49154 52054
rect 49206 52002 49365 52054
rect 49417 52002 49576 52054
rect 49628 52002 49787 52054
rect 49839 52002 49991 52054
rect 48557 51949 48687 51988
rect 48557 51893 48594 51949
rect 48650 51893 48687 51949
rect 48557 51731 48687 51893
rect 48557 51675 48594 51731
rect 48650 51675 48687 51731
rect 48557 51637 48687 51675
rect 48790 51591 49991 52002
rect 48790 51539 48943 51591
rect 48995 51539 49154 51591
rect 49206 51539 49365 51591
rect 49417 51539 49576 51591
rect 49628 51539 49787 51591
rect 49839 51539 49991 51591
rect 48790 51315 49991 51539
rect 48790 51263 48943 51315
rect 48995 51263 49154 51315
rect 49206 51263 49365 51315
rect 49417 51263 49576 51315
rect 49628 51263 49787 51315
rect 49839 51263 49991 51315
rect 48158 51079 48241 51131
rect 48293 51079 48379 51131
rect 48158 43931 48379 51079
rect 48557 51179 48687 51217
rect 48557 51123 48594 51179
rect 48650 51123 48687 51179
rect 48557 50961 48687 51123
rect 48557 50905 48594 50961
rect 48650 50905 48687 50961
rect 48557 50866 48687 50905
rect 48790 50852 49991 51263
rect 48790 50800 48943 50852
rect 48995 50800 49154 50852
rect 49206 50800 49365 50852
rect 49417 50800 49576 50852
rect 49628 50800 49787 50852
rect 49839 50800 49991 50852
rect 48790 50555 49991 50800
rect 48790 50499 48836 50555
rect 48892 50499 49046 50555
rect 49102 50499 49257 50555
rect 49313 50499 49469 50555
rect 49525 50499 49680 50555
rect 49736 50499 49890 50555
rect 49946 50499 49991 50555
rect 48790 50254 49991 50499
rect 48790 50202 48943 50254
rect 48995 50202 49154 50254
rect 49206 50202 49365 50254
rect 49417 50202 49576 50254
rect 49628 50202 49787 50254
rect 49839 50202 49991 50254
rect 48557 50149 48687 50188
rect 48557 50093 48594 50149
rect 48650 50093 48687 50149
rect 48557 49931 48687 50093
rect 48557 49875 48594 49931
rect 48650 49875 48687 49931
rect 48557 49837 48687 49875
rect 48790 49791 49991 50202
rect 48790 49739 48943 49791
rect 48995 49739 49154 49791
rect 49206 49739 49365 49791
rect 49417 49739 49576 49791
rect 49628 49739 49787 49791
rect 49839 49739 49991 49791
rect 48790 49515 49991 49739
rect 48790 49463 48943 49515
rect 48995 49463 49154 49515
rect 49206 49463 49365 49515
rect 49417 49463 49576 49515
rect 49628 49463 49787 49515
rect 49839 49463 49991 49515
rect 48557 49379 48687 49417
rect 48557 49323 48594 49379
rect 48650 49323 48687 49379
rect 48557 49161 48687 49323
rect 48557 49105 48594 49161
rect 48650 49105 48687 49161
rect 48557 49066 48687 49105
rect 48790 49052 49991 49463
rect 48790 49000 48943 49052
rect 48995 49000 49154 49052
rect 49206 49000 49365 49052
rect 49417 49000 49576 49052
rect 49628 49000 49787 49052
rect 49839 49000 49991 49052
rect 48790 48755 49991 49000
rect 48790 48699 48836 48755
rect 48892 48699 49046 48755
rect 49102 48699 49257 48755
rect 49313 48699 49469 48755
rect 49525 48699 49680 48755
rect 49736 48699 49890 48755
rect 49946 48699 49991 48755
rect 48790 48454 49991 48699
rect 48790 48402 48943 48454
rect 48995 48402 49154 48454
rect 49206 48402 49365 48454
rect 49417 48402 49576 48454
rect 49628 48402 49787 48454
rect 49839 48402 49991 48454
rect 48557 48349 48687 48388
rect 48557 48293 48594 48349
rect 48650 48293 48687 48349
rect 48557 48131 48687 48293
rect 48557 48075 48594 48131
rect 48650 48075 48687 48131
rect 48557 48037 48687 48075
rect 48790 47991 49991 48402
rect 48790 47939 48943 47991
rect 48995 47939 49154 47991
rect 49206 47939 49365 47991
rect 49417 47939 49576 47991
rect 49628 47939 49787 47991
rect 49839 47939 49991 47991
rect 48790 47715 49991 47939
rect 48790 47663 48943 47715
rect 48995 47663 49154 47715
rect 49206 47663 49365 47715
rect 49417 47663 49576 47715
rect 49628 47663 49787 47715
rect 49839 47663 49991 47715
rect 48557 47579 48687 47617
rect 48557 47523 48594 47579
rect 48650 47523 48687 47579
rect 48557 47361 48687 47523
rect 48557 47305 48594 47361
rect 48650 47305 48687 47361
rect 48557 47266 48687 47305
rect 48790 47252 49991 47663
rect 48790 47200 48943 47252
rect 48995 47200 49154 47252
rect 49206 47200 49365 47252
rect 49417 47200 49576 47252
rect 49628 47200 49787 47252
rect 49839 47200 49991 47252
rect 48790 46955 49991 47200
rect 48790 46899 48836 46955
rect 48892 46899 49046 46955
rect 49102 46899 49257 46955
rect 49313 46899 49469 46955
rect 49525 46899 49680 46955
rect 49736 46899 49890 46955
rect 49946 46899 49991 46955
rect 48790 46654 49991 46899
rect 48790 46602 48943 46654
rect 48995 46602 49154 46654
rect 49206 46602 49365 46654
rect 49417 46602 49576 46654
rect 49628 46602 49787 46654
rect 49839 46602 49991 46654
rect 48557 46549 48687 46588
rect 48557 46493 48594 46549
rect 48650 46493 48687 46549
rect 48557 46331 48687 46493
rect 48557 46275 48594 46331
rect 48650 46275 48687 46331
rect 48557 46237 48687 46275
rect 48790 46191 49991 46602
rect 48790 46139 48943 46191
rect 48995 46139 49154 46191
rect 49206 46139 49365 46191
rect 49417 46139 49576 46191
rect 49628 46139 49787 46191
rect 49839 46139 49991 46191
rect 48790 45915 49991 46139
rect 48790 45863 48943 45915
rect 48995 45863 49154 45915
rect 49206 45863 49365 45915
rect 49417 45863 49576 45915
rect 49628 45863 49787 45915
rect 49839 45863 49991 45915
rect 48557 45779 48687 45817
rect 48557 45723 48594 45779
rect 48650 45723 48687 45779
rect 48557 45561 48687 45723
rect 48557 45505 48594 45561
rect 48650 45505 48687 45561
rect 48557 45466 48687 45505
rect 48790 45452 49991 45863
rect 48790 45400 48943 45452
rect 48995 45400 49154 45452
rect 49206 45400 49365 45452
rect 49417 45400 49576 45452
rect 49628 45400 49787 45452
rect 49839 45400 49991 45452
rect 48790 45155 49991 45400
rect 48790 45099 48836 45155
rect 48892 45099 49046 45155
rect 49102 45099 49257 45155
rect 49313 45099 49469 45155
rect 49525 45099 49680 45155
rect 49736 45099 49890 45155
rect 49946 45099 49991 45155
rect 48790 44854 49991 45099
rect 48790 44802 48943 44854
rect 48995 44802 49154 44854
rect 49206 44802 49365 44854
rect 49417 44802 49576 44854
rect 49628 44802 49787 44854
rect 49839 44802 49991 44854
rect 48557 44749 48687 44788
rect 48557 44693 48594 44749
rect 48650 44693 48687 44749
rect 48557 44531 48687 44693
rect 48557 44475 48594 44531
rect 48650 44475 48687 44531
rect 48557 44437 48687 44475
rect 48790 44391 49991 44802
rect 48790 44339 48943 44391
rect 48995 44339 49154 44391
rect 49206 44339 49365 44391
rect 49417 44339 49576 44391
rect 49628 44339 49787 44391
rect 49839 44339 49991 44391
rect 48790 44115 49991 44339
rect 48790 44063 48943 44115
rect 48995 44063 49154 44115
rect 49206 44063 49365 44115
rect 49417 44063 49576 44115
rect 49628 44063 49787 44115
rect 49839 44063 49991 44115
rect 48158 43879 48241 43931
rect 48293 43879 48379 43931
rect 48158 36731 48379 43879
rect 48557 43979 48687 44017
rect 48557 43923 48594 43979
rect 48650 43923 48687 43979
rect 48557 43761 48687 43923
rect 48557 43705 48594 43761
rect 48650 43705 48687 43761
rect 48557 43666 48687 43705
rect 48790 43652 49991 44063
rect 48790 43600 48943 43652
rect 48995 43600 49154 43652
rect 49206 43600 49365 43652
rect 49417 43600 49576 43652
rect 49628 43600 49787 43652
rect 49839 43600 49991 43652
rect 48790 43355 49991 43600
rect 48790 43299 48836 43355
rect 48892 43299 49046 43355
rect 49102 43299 49257 43355
rect 49313 43299 49469 43355
rect 49525 43299 49680 43355
rect 49736 43299 49890 43355
rect 49946 43299 49991 43355
rect 48790 43054 49991 43299
rect 48790 43002 48943 43054
rect 48995 43002 49154 43054
rect 49206 43002 49365 43054
rect 49417 43002 49576 43054
rect 49628 43002 49787 43054
rect 49839 43002 49991 43054
rect 48557 42949 48687 42988
rect 48557 42893 48594 42949
rect 48650 42893 48687 42949
rect 48557 42731 48687 42893
rect 48557 42675 48594 42731
rect 48650 42675 48687 42731
rect 48557 42637 48687 42675
rect 48790 42591 49991 43002
rect 48790 42539 48943 42591
rect 48995 42539 49154 42591
rect 49206 42539 49365 42591
rect 49417 42539 49576 42591
rect 49628 42539 49787 42591
rect 49839 42539 49991 42591
rect 48790 42315 49991 42539
rect 48790 42263 48943 42315
rect 48995 42263 49154 42315
rect 49206 42263 49365 42315
rect 49417 42263 49576 42315
rect 49628 42263 49787 42315
rect 49839 42263 49991 42315
rect 48557 42179 48687 42217
rect 48557 42123 48594 42179
rect 48650 42123 48687 42179
rect 48557 41961 48687 42123
rect 48557 41905 48594 41961
rect 48650 41905 48687 41961
rect 48557 41866 48687 41905
rect 48790 41852 49991 42263
rect 48790 41800 48943 41852
rect 48995 41800 49154 41852
rect 49206 41800 49365 41852
rect 49417 41800 49576 41852
rect 49628 41800 49787 41852
rect 49839 41800 49991 41852
rect 48790 41555 49991 41800
rect 48790 41499 48836 41555
rect 48892 41499 49046 41555
rect 49102 41499 49257 41555
rect 49313 41499 49469 41555
rect 49525 41499 49680 41555
rect 49736 41499 49890 41555
rect 49946 41499 49991 41555
rect 48790 41254 49991 41499
rect 48790 41202 48943 41254
rect 48995 41202 49154 41254
rect 49206 41202 49365 41254
rect 49417 41202 49576 41254
rect 49628 41202 49787 41254
rect 49839 41202 49991 41254
rect 48557 41149 48687 41188
rect 48557 41093 48594 41149
rect 48650 41093 48687 41149
rect 48557 40931 48687 41093
rect 48557 40875 48594 40931
rect 48650 40875 48687 40931
rect 48557 40837 48687 40875
rect 48790 40791 49991 41202
rect 48790 40739 48943 40791
rect 48995 40739 49154 40791
rect 49206 40739 49365 40791
rect 49417 40739 49576 40791
rect 49628 40739 49787 40791
rect 49839 40739 49991 40791
rect 48790 40515 49991 40739
rect 48790 40463 48943 40515
rect 48995 40463 49154 40515
rect 49206 40463 49365 40515
rect 49417 40463 49576 40515
rect 49628 40463 49787 40515
rect 49839 40463 49991 40515
rect 48557 40379 48687 40417
rect 48557 40323 48594 40379
rect 48650 40323 48687 40379
rect 48557 40161 48687 40323
rect 48557 40105 48594 40161
rect 48650 40105 48687 40161
rect 48557 40066 48687 40105
rect 48790 40052 49991 40463
rect 48790 40000 48943 40052
rect 48995 40000 49154 40052
rect 49206 40000 49365 40052
rect 49417 40000 49576 40052
rect 49628 40000 49787 40052
rect 49839 40000 49991 40052
rect 48790 39755 49991 40000
rect 48790 39699 48836 39755
rect 48892 39699 49046 39755
rect 49102 39699 49257 39755
rect 49313 39699 49469 39755
rect 49525 39699 49680 39755
rect 49736 39699 49890 39755
rect 49946 39699 49991 39755
rect 48790 39454 49991 39699
rect 48790 39402 48943 39454
rect 48995 39402 49154 39454
rect 49206 39402 49365 39454
rect 49417 39402 49576 39454
rect 49628 39402 49787 39454
rect 49839 39402 49991 39454
rect 48557 39349 48687 39388
rect 48557 39293 48594 39349
rect 48650 39293 48687 39349
rect 48557 39131 48687 39293
rect 48557 39075 48594 39131
rect 48650 39075 48687 39131
rect 48557 39037 48687 39075
rect 48790 38991 49991 39402
rect 48790 38939 48943 38991
rect 48995 38939 49154 38991
rect 49206 38939 49365 38991
rect 49417 38939 49576 38991
rect 49628 38939 49787 38991
rect 49839 38939 49991 38991
rect 48790 38715 49991 38939
rect 48790 38663 48943 38715
rect 48995 38663 49154 38715
rect 49206 38663 49365 38715
rect 49417 38663 49576 38715
rect 49628 38663 49787 38715
rect 49839 38663 49991 38715
rect 48557 38579 48687 38617
rect 48557 38523 48594 38579
rect 48650 38523 48687 38579
rect 48557 38361 48687 38523
rect 48557 38305 48594 38361
rect 48650 38305 48687 38361
rect 48557 38266 48687 38305
rect 48790 38252 49991 38663
rect 48790 38200 48943 38252
rect 48995 38200 49154 38252
rect 49206 38200 49365 38252
rect 49417 38200 49576 38252
rect 49628 38200 49787 38252
rect 49839 38200 49991 38252
rect 48790 37955 49991 38200
rect 48790 37899 48836 37955
rect 48892 37899 49046 37955
rect 49102 37899 49257 37955
rect 49313 37899 49469 37955
rect 49525 37899 49680 37955
rect 49736 37899 49890 37955
rect 49946 37899 49991 37955
rect 48790 37654 49991 37899
rect 48790 37602 48943 37654
rect 48995 37602 49154 37654
rect 49206 37602 49365 37654
rect 49417 37602 49576 37654
rect 49628 37602 49787 37654
rect 49839 37602 49991 37654
rect 48557 37549 48687 37588
rect 48557 37493 48594 37549
rect 48650 37493 48687 37549
rect 48557 37331 48687 37493
rect 48557 37275 48594 37331
rect 48650 37275 48687 37331
rect 48557 37237 48687 37275
rect 48790 37191 49991 37602
rect 48790 37139 48943 37191
rect 48995 37139 49154 37191
rect 49206 37139 49365 37191
rect 49417 37139 49576 37191
rect 49628 37139 49787 37191
rect 49839 37139 49991 37191
rect 48790 36915 49991 37139
rect 48790 36863 48943 36915
rect 48995 36863 49154 36915
rect 49206 36863 49365 36915
rect 49417 36863 49576 36915
rect 49628 36863 49787 36915
rect 49839 36863 49991 36915
rect 48158 36679 48241 36731
rect 48293 36679 48379 36731
rect 48158 36096 48379 36679
rect 48557 36779 48687 36817
rect 48557 36723 48594 36779
rect 48650 36723 48687 36779
rect 48557 36561 48687 36723
rect 48557 36505 48594 36561
rect 48650 36505 48687 36561
rect 48557 36466 48687 36505
rect 47779 35963 48002 36096
rect 47402 35171 47623 35963
rect 47779 35507 48001 35963
rect 48157 35842 48379 36096
rect 48790 36452 49991 36863
rect 48790 36400 48943 36452
rect 48995 36400 49154 36452
rect 49206 36400 49365 36452
rect 49417 36400 49576 36452
rect 49628 36400 49787 36452
rect 49839 36400 49991 36452
rect 48790 36155 49991 36400
rect 48790 36099 48836 36155
rect 48892 36099 49046 36155
rect 49102 36099 49257 36155
rect 49313 36099 49469 36155
rect 49525 36099 49680 36155
rect 49736 36099 49890 36155
rect 49946 36099 49991 36155
rect 48790 35976 49991 36099
rect 50099 64901 50346 64940
rect 50398 64901 50557 64953
rect 50609 64901 50768 64953
rect 50820 64901 50913 64953
rect 52226 65078 54354 65366
rect 54758 65853 55638 66376
rect 54758 65801 54855 65853
rect 54907 65801 55066 65853
rect 55118 65801 55278 65853
rect 55330 65801 55489 65853
rect 55541 65801 55638 65853
rect 52226 64955 54355 65078
rect 52226 64940 52314 64955
rect 50099 64491 50913 64901
rect 52227 64899 52314 64940
rect 52370 64899 52525 64955
rect 52581 64899 52736 64955
rect 52792 64899 52946 64955
rect 53002 64899 53157 64955
rect 53213 64899 53369 64955
rect 53425 64899 53580 64955
rect 53636 64899 53790 64955
rect 53846 64899 54001 64955
rect 54057 64899 54212 64955
rect 54268 64899 54355 64955
rect 50099 64439 50300 64491
rect 50352 64439 50511 64491
rect 50563 64439 50722 64491
rect 50774 64439 50913 64491
rect 50099 64055 50913 64439
rect 51034 64729 51344 64770
rect 51034 64677 51073 64729
rect 51125 64677 51253 64729
rect 51305 64677 51344 64729
rect 51034 64515 51344 64677
rect 51034 64459 51071 64515
rect 51127 64459 51251 64515
rect 51307 64459 51344 64515
rect 51034 64386 51344 64459
rect 51796 64722 52106 64763
rect 51796 64670 51835 64722
rect 51887 64670 52015 64722
rect 52067 64670 52106 64722
rect 51796 64515 52106 64670
rect 51796 64459 51833 64515
rect 51889 64459 52013 64515
rect 52069 64459 52106 64515
rect 51796 64259 52106 64459
rect 51796 64207 51835 64259
rect 51887 64207 52015 64259
rect 52067 64207 52106 64259
rect 51796 64167 52106 64207
rect 50099 64053 50161 64055
rect 50217 64053 50372 64055
rect 50099 64001 50138 64053
rect 50217 64001 50318 64053
rect 50370 64001 50372 64053
rect 50099 63999 50161 64001
rect 50217 63999 50372 64001
rect 50428 63999 50584 64055
rect 50640 63999 50795 64055
rect 50851 63999 50913 64055
rect 50099 63615 50913 63999
rect 52227 64053 54355 64899
rect 52227 64001 52316 64053
rect 52368 64001 52527 64053
rect 52579 64001 52738 64053
rect 52790 64001 52948 64053
rect 53000 64001 53159 64053
rect 53211 64001 53371 64053
rect 53423 64001 53582 64053
rect 53634 64001 53792 64053
rect 53844 64001 54003 64053
rect 54055 64001 54214 64053
rect 54266 64001 54355 64053
rect 51796 63847 52106 63887
rect 51796 63795 51835 63847
rect 51887 63795 52015 63847
rect 52067 63795 52106 63847
rect 50099 63563 50300 63615
rect 50352 63563 50511 63615
rect 50563 63563 50722 63615
rect 50774 63563 50913 63615
rect 50099 63153 50913 63563
rect 51034 63595 51344 63668
rect 51034 63539 51071 63595
rect 51127 63539 51251 63595
rect 51307 63539 51344 63595
rect 51034 63377 51344 63539
rect 51034 63325 51073 63377
rect 51125 63325 51253 63377
rect 51305 63325 51344 63377
rect 51034 63284 51344 63325
rect 51796 63595 52106 63795
rect 51796 63539 51833 63595
rect 51889 63539 52013 63595
rect 52069 63539 52106 63595
rect 51796 63384 52106 63539
rect 51796 63332 51835 63384
rect 51887 63332 52015 63384
rect 52067 63332 52106 63384
rect 51796 63291 52106 63332
rect 50099 63101 50346 63153
rect 50398 63101 50557 63153
rect 50609 63101 50768 63153
rect 50820 63101 50913 63153
rect 50099 62691 50913 63101
rect 52227 63155 54355 64001
rect 52227 63099 52314 63155
rect 52370 63099 52525 63155
rect 52581 63099 52736 63155
rect 52792 63099 52946 63155
rect 53002 63099 53157 63155
rect 53213 63099 53369 63155
rect 53425 63099 53580 63155
rect 53636 63099 53790 63155
rect 53846 63099 54001 63155
rect 54057 63099 54212 63155
rect 54268 63099 54355 63155
rect 50099 62639 50300 62691
rect 50352 62639 50511 62691
rect 50563 62639 50722 62691
rect 50774 62639 50913 62691
rect 50099 62255 50913 62639
rect 51034 62929 51344 62970
rect 51034 62877 51073 62929
rect 51125 62877 51253 62929
rect 51305 62877 51344 62929
rect 51034 62715 51344 62877
rect 51034 62659 51071 62715
rect 51127 62659 51251 62715
rect 51307 62659 51344 62715
rect 51034 62586 51344 62659
rect 51796 62922 52106 62963
rect 51796 62870 51835 62922
rect 51887 62870 52015 62922
rect 52067 62870 52106 62922
rect 51796 62715 52106 62870
rect 51796 62659 51833 62715
rect 51889 62659 52013 62715
rect 52069 62659 52106 62715
rect 51796 62459 52106 62659
rect 51796 62407 51835 62459
rect 51887 62407 52015 62459
rect 52067 62407 52106 62459
rect 51796 62367 52106 62407
rect 50099 62253 50161 62255
rect 50217 62253 50372 62255
rect 50099 62201 50138 62253
rect 50217 62201 50318 62253
rect 50370 62201 50372 62253
rect 50099 62199 50161 62201
rect 50217 62199 50372 62201
rect 50428 62199 50584 62255
rect 50640 62199 50795 62255
rect 50851 62199 50913 62255
rect 50099 61815 50913 62199
rect 52227 62253 54355 63099
rect 52227 62201 52316 62253
rect 52368 62201 52527 62253
rect 52579 62201 52738 62253
rect 52790 62201 52948 62253
rect 53000 62201 53159 62253
rect 53211 62201 53371 62253
rect 53423 62201 53582 62253
rect 53634 62201 53792 62253
rect 53844 62201 54003 62253
rect 54055 62201 54214 62253
rect 54266 62201 54355 62253
rect 51796 62047 52106 62087
rect 51796 61995 51835 62047
rect 51887 61995 52015 62047
rect 52067 61995 52106 62047
rect 50099 61763 50300 61815
rect 50352 61763 50511 61815
rect 50563 61763 50722 61815
rect 50774 61763 50913 61815
rect 50099 61353 50913 61763
rect 51034 61795 51344 61868
rect 51034 61739 51071 61795
rect 51127 61739 51251 61795
rect 51307 61739 51344 61795
rect 51034 61577 51344 61739
rect 51034 61525 51073 61577
rect 51125 61525 51253 61577
rect 51305 61525 51344 61577
rect 51034 61484 51344 61525
rect 51796 61795 52106 61995
rect 51796 61739 51833 61795
rect 51889 61739 52013 61795
rect 52069 61739 52106 61795
rect 51796 61584 52106 61739
rect 51796 61532 51835 61584
rect 51887 61532 52015 61584
rect 52067 61532 52106 61584
rect 51796 61491 52106 61532
rect 50099 61301 50346 61353
rect 50398 61301 50557 61353
rect 50609 61301 50768 61353
rect 50820 61301 50913 61353
rect 50099 60891 50913 61301
rect 52227 61355 54355 62201
rect 52227 61299 52314 61355
rect 52370 61299 52525 61355
rect 52581 61299 52736 61355
rect 52792 61299 52946 61355
rect 53002 61299 53157 61355
rect 53213 61299 53369 61355
rect 53425 61299 53580 61355
rect 53636 61299 53790 61355
rect 53846 61299 54001 61355
rect 54057 61299 54212 61355
rect 54268 61299 54355 61355
rect 50099 60839 50300 60891
rect 50352 60839 50511 60891
rect 50563 60839 50722 60891
rect 50774 60839 50913 60891
rect 50099 60455 50913 60839
rect 51034 61129 51344 61170
rect 51034 61077 51073 61129
rect 51125 61077 51253 61129
rect 51305 61077 51344 61129
rect 51034 60915 51344 61077
rect 51034 60859 51071 60915
rect 51127 60859 51251 60915
rect 51307 60859 51344 60915
rect 51034 60786 51344 60859
rect 51796 61122 52106 61163
rect 51796 61070 51835 61122
rect 51887 61070 52015 61122
rect 52067 61070 52106 61122
rect 51796 60915 52106 61070
rect 51796 60859 51833 60915
rect 51889 60859 52013 60915
rect 52069 60859 52106 60915
rect 51796 60659 52106 60859
rect 51796 60607 51835 60659
rect 51887 60607 52015 60659
rect 52067 60607 52106 60659
rect 51796 60567 52106 60607
rect 50099 60453 50161 60455
rect 50217 60453 50372 60455
rect 50099 60401 50138 60453
rect 50217 60401 50318 60453
rect 50370 60401 50372 60453
rect 50099 60399 50161 60401
rect 50217 60399 50372 60401
rect 50428 60399 50584 60455
rect 50640 60399 50795 60455
rect 50851 60399 50913 60455
rect 50099 60015 50913 60399
rect 52227 60453 54355 61299
rect 52227 60401 52316 60453
rect 52368 60401 52527 60453
rect 52579 60401 52738 60453
rect 52790 60401 52948 60453
rect 53000 60401 53159 60453
rect 53211 60401 53371 60453
rect 53423 60401 53582 60453
rect 53634 60401 53792 60453
rect 53844 60401 54003 60453
rect 54055 60401 54214 60453
rect 54266 60401 54355 60453
rect 51796 60247 52106 60287
rect 51796 60195 51835 60247
rect 51887 60195 52015 60247
rect 52067 60195 52106 60247
rect 50099 59963 50300 60015
rect 50352 59963 50511 60015
rect 50563 59963 50722 60015
rect 50774 59963 50913 60015
rect 50099 59553 50913 59963
rect 51034 59995 51344 60068
rect 51034 59939 51071 59995
rect 51127 59939 51251 59995
rect 51307 59939 51344 59995
rect 51034 59777 51344 59939
rect 51034 59725 51073 59777
rect 51125 59725 51253 59777
rect 51305 59725 51344 59777
rect 51034 59684 51344 59725
rect 51796 59995 52106 60195
rect 51796 59939 51833 59995
rect 51889 59939 52013 59995
rect 52069 59939 52106 59995
rect 51796 59784 52106 59939
rect 51796 59732 51835 59784
rect 51887 59732 52015 59784
rect 52067 59732 52106 59784
rect 51796 59691 52106 59732
rect 50099 59501 50346 59553
rect 50398 59501 50557 59553
rect 50609 59501 50768 59553
rect 50820 59501 50913 59553
rect 50099 59091 50913 59501
rect 52227 59555 54355 60401
rect 52227 59499 52314 59555
rect 52370 59499 52525 59555
rect 52581 59499 52736 59555
rect 52792 59499 52946 59555
rect 53002 59499 53157 59555
rect 53213 59499 53369 59555
rect 53425 59499 53580 59555
rect 53636 59499 53790 59555
rect 53846 59499 54001 59555
rect 54057 59499 54212 59555
rect 54268 59499 54355 59555
rect 50099 59039 50300 59091
rect 50352 59039 50511 59091
rect 50563 59039 50722 59091
rect 50774 59039 50913 59091
rect 50099 58655 50913 59039
rect 51034 59329 51344 59370
rect 51034 59277 51073 59329
rect 51125 59277 51253 59329
rect 51305 59277 51344 59329
rect 51034 59115 51344 59277
rect 51034 59059 51071 59115
rect 51127 59059 51251 59115
rect 51307 59059 51344 59115
rect 51034 58986 51344 59059
rect 51796 59322 52106 59363
rect 51796 59270 51835 59322
rect 51887 59270 52015 59322
rect 52067 59270 52106 59322
rect 51796 59115 52106 59270
rect 51796 59059 51833 59115
rect 51889 59059 52013 59115
rect 52069 59059 52106 59115
rect 51796 58859 52106 59059
rect 51796 58807 51835 58859
rect 51887 58807 52015 58859
rect 52067 58807 52106 58859
rect 51796 58767 52106 58807
rect 50099 58653 50161 58655
rect 50217 58653 50372 58655
rect 50099 58601 50138 58653
rect 50217 58601 50318 58653
rect 50370 58601 50372 58653
rect 50099 58599 50161 58601
rect 50217 58599 50372 58601
rect 50428 58599 50584 58655
rect 50640 58599 50795 58655
rect 50851 58599 50913 58655
rect 50099 58215 50913 58599
rect 52227 58653 54355 59499
rect 52227 58601 52316 58653
rect 52368 58601 52527 58653
rect 52579 58601 52738 58653
rect 52790 58601 52948 58653
rect 53000 58601 53159 58653
rect 53211 58601 53371 58653
rect 53423 58601 53582 58653
rect 53634 58601 53792 58653
rect 53844 58601 54003 58653
rect 54055 58601 54214 58653
rect 54266 58601 54355 58653
rect 51796 58447 52106 58487
rect 51796 58395 51835 58447
rect 51887 58395 52015 58447
rect 52067 58395 52106 58447
rect 50099 58163 50300 58215
rect 50352 58163 50511 58215
rect 50563 58163 50722 58215
rect 50774 58163 50913 58215
rect 50099 57753 50913 58163
rect 51034 58195 51344 58268
rect 51034 58139 51071 58195
rect 51127 58139 51251 58195
rect 51307 58139 51344 58195
rect 51034 57977 51344 58139
rect 51034 57925 51073 57977
rect 51125 57925 51253 57977
rect 51305 57925 51344 57977
rect 51034 57884 51344 57925
rect 51796 58195 52106 58395
rect 51796 58139 51833 58195
rect 51889 58139 52013 58195
rect 52069 58139 52106 58195
rect 51796 57984 52106 58139
rect 51796 57932 51835 57984
rect 51887 57932 52015 57984
rect 52067 57932 52106 57984
rect 51796 57891 52106 57932
rect 50099 57701 50346 57753
rect 50398 57701 50557 57753
rect 50609 57701 50768 57753
rect 50820 57701 50913 57753
rect 50099 57291 50913 57701
rect 52227 57755 54355 58601
rect 52227 57699 52314 57755
rect 52370 57699 52525 57755
rect 52581 57699 52736 57755
rect 52792 57699 52946 57755
rect 53002 57699 53157 57755
rect 53213 57699 53369 57755
rect 53425 57699 53580 57755
rect 53636 57699 53790 57755
rect 53846 57699 54001 57755
rect 54057 57699 54212 57755
rect 54268 57699 54355 57755
rect 50099 57239 50300 57291
rect 50352 57239 50511 57291
rect 50563 57239 50722 57291
rect 50774 57239 50913 57291
rect 50099 56855 50913 57239
rect 51034 57529 51344 57570
rect 51034 57477 51073 57529
rect 51125 57477 51253 57529
rect 51305 57477 51344 57529
rect 51034 57315 51344 57477
rect 51034 57259 51071 57315
rect 51127 57259 51251 57315
rect 51307 57259 51344 57315
rect 51034 57186 51344 57259
rect 51796 57522 52106 57563
rect 51796 57470 51835 57522
rect 51887 57470 52015 57522
rect 52067 57470 52106 57522
rect 51796 57315 52106 57470
rect 51796 57259 51833 57315
rect 51889 57259 52013 57315
rect 52069 57259 52106 57315
rect 51796 57059 52106 57259
rect 51796 57007 51835 57059
rect 51887 57007 52015 57059
rect 52067 57007 52106 57059
rect 51796 56967 52106 57007
rect 50099 56853 50161 56855
rect 50217 56853 50372 56855
rect 50099 56801 50138 56853
rect 50217 56801 50318 56853
rect 50370 56801 50372 56853
rect 50099 56799 50161 56801
rect 50217 56799 50372 56801
rect 50428 56799 50584 56855
rect 50640 56799 50795 56855
rect 50851 56799 50913 56855
rect 50099 56415 50913 56799
rect 52227 56853 54355 57699
rect 52227 56801 52316 56853
rect 52368 56801 52527 56853
rect 52579 56801 52738 56853
rect 52790 56801 52948 56853
rect 53000 56801 53159 56853
rect 53211 56801 53371 56853
rect 53423 56801 53582 56853
rect 53634 56801 53792 56853
rect 53844 56801 54003 56853
rect 54055 56801 54214 56853
rect 54266 56801 54355 56853
rect 51796 56647 52106 56687
rect 51796 56595 51835 56647
rect 51887 56595 52015 56647
rect 52067 56595 52106 56647
rect 50099 56363 50300 56415
rect 50352 56363 50511 56415
rect 50563 56363 50722 56415
rect 50774 56363 50913 56415
rect 50099 55953 50913 56363
rect 51034 56395 51344 56468
rect 51034 56339 51071 56395
rect 51127 56339 51251 56395
rect 51307 56339 51344 56395
rect 51034 56177 51344 56339
rect 51034 56125 51073 56177
rect 51125 56125 51253 56177
rect 51305 56125 51344 56177
rect 51034 56084 51344 56125
rect 51796 56395 52106 56595
rect 51796 56339 51833 56395
rect 51889 56339 52013 56395
rect 52069 56339 52106 56395
rect 51796 56184 52106 56339
rect 51796 56132 51835 56184
rect 51887 56132 52015 56184
rect 52067 56132 52106 56184
rect 51796 56091 52106 56132
rect 50099 55901 50346 55953
rect 50398 55901 50557 55953
rect 50609 55901 50768 55953
rect 50820 55901 50913 55953
rect 50099 55491 50913 55901
rect 52227 55955 54355 56801
rect 52227 55899 52314 55955
rect 52370 55899 52525 55955
rect 52581 55899 52736 55955
rect 52792 55899 52946 55955
rect 53002 55899 53157 55955
rect 53213 55899 53369 55955
rect 53425 55899 53580 55955
rect 53636 55899 53790 55955
rect 53846 55899 54001 55955
rect 54057 55899 54212 55955
rect 54268 55899 54355 55955
rect 50099 55439 50300 55491
rect 50352 55439 50511 55491
rect 50563 55439 50722 55491
rect 50774 55439 50913 55491
rect 50099 55055 50913 55439
rect 51034 55729 51344 55770
rect 51034 55677 51073 55729
rect 51125 55677 51253 55729
rect 51305 55677 51344 55729
rect 51034 55515 51344 55677
rect 51034 55459 51071 55515
rect 51127 55459 51251 55515
rect 51307 55459 51344 55515
rect 51034 55386 51344 55459
rect 51796 55722 52106 55763
rect 51796 55670 51835 55722
rect 51887 55670 52015 55722
rect 52067 55670 52106 55722
rect 51796 55515 52106 55670
rect 51796 55459 51833 55515
rect 51889 55459 52013 55515
rect 52069 55459 52106 55515
rect 51796 55259 52106 55459
rect 51796 55207 51835 55259
rect 51887 55207 52015 55259
rect 52067 55207 52106 55259
rect 51796 55167 52106 55207
rect 50099 55053 50161 55055
rect 50217 55053 50372 55055
rect 50099 55001 50138 55053
rect 50217 55001 50318 55053
rect 50370 55001 50372 55053
rect 50099 54999 50161 55001
rect 50217 54999 50372 55001
rect 50428 54999 50584 55055
rect 50640 54999 50795 55055
rect 50851 54999 50913 55055
rect 50099 54615 50913 54999
rect 52227 55053 54355 55899
rect 52227 55001 52316 55053
rect 52368 55001 52527 55053
rect 52579 55001 52738 55053
rect 52790 55001 52948 55053
rect 53000 55001 53159 55053
rect 53211 55001 53371 55053
rect 53423 55001 53582 55053
rect 53634 55001 53792 55053
rect 53844 55001 54003 55053
rect 54055 55001 54214 55053
rect 54266 55001 54355 55053
rect 51796 54847 52106 54887
rect 51796 54795 51835 54847
rect 51887 54795 52015 54847
rect 52067 54795 52106 54847
rect 50099 54563 50300 54615
rect 50352 54563 50511 54615
rect 50563 54563 50722 54615
rect 50774 54563 50913 54615
rect 50099 54153 50913 54563
rect 51034 54595 51344 54668
rect 51034 54539 51071 54595
rect 51127 54539 51251 54595
rect 51307 54539 51344 54595
rect 51034 54377 51344 54539
rect 51034 54325 51073 54377
rect 51125 54325 51253 54377
rect 51305 54325 51344 54377
rect 51034 54284 51344 54325
rect 51796 54595 52106 54795
rect 51796 54539 51833 54595
rect 51889 54539 52013 54595
rect 52069 54539 52106 54595
rect 51796 54384 52106 54539
rect 51796 54332 51835 54384
rect 51887 54332 52015 54384
rect 52067 54332 52106 54384
rect 51796 54291 52106 54332
rect 50099 54101 50346 54153
rect 50398 54101 50557 54153
rect 50609 54101 50768 54153
rect 50820 54101 50913 54153
rect 50099 53691 50913 54101
rect 52227 54155 54355 55001
rect 52227 54099 52314 54155
rect 52370 54099 52525 54155
rect 52581 54099 52736 54155
rect 52792 54099 52946 54155
rect 53002 54099 53157 54155
rect 53213 54099 53369 54155
rect 53425 54099 53580 54155
rect 53636 54099 53790 54155
rect 53846 54099 54001 54155
rect 54057 54099 54212 54155
rect 54268 54099 54355 54155
rect 50099 53639 50300 53691
rect 50352 53639 50511 53691
rect 50563 53639 50722 53691
rect 50774 53639 50913 53691
rect 50099 53255 50913 53639
rect 51034 53929 51344 53970
rect 51034 53877 51073 53929
rect 51125 53877 51253 53929
rect 51305 53877 51344 53929
rect 51034 53715 51344 53877
rect 51034 53659 51071 53715
rect 51127 53659 51251 53715
rect 51307 53659 51344 53715
rect 51034 53586 51344 53659
rect 51796 53922 52106 53963
rect 51796 53870 51835 53922
rect 51887 53870 52015 53922
rect 52067 53870 52106 53922
rect 51796 53715 52106 53870
rect 51796 53659 51833 53715
rect 51889 53659 52013 53715
rect 52069 53659 52106 53715
rect 51796 53459 52106 53659
rect 51796 53407 51835 53459
rect 51887 53407 52015 53459
rect 52067 53407 52106 53459
rect 51796 53367 52106 53407
rect 50099 53253 50161 53255
rect 50217 53253 50372 53255
rect 50099 53201 50138 53253
rect 50217 53201 50318 53253
rect 50370 53201 50372 53253
rect 50099 53199 50161 53201
rect 50217 53199 50372 53201
rect 50428 53199 50584 53255
rect 50640 53199 50795 53255
rect 50851 53199 50913 53255
rect 50099 52815 50913 53199
rect 52227 53253 54355 54099
rect 52227 53201 52316 53253
rect 52368 53201 52527 53253
rect 52579 53201 52738 53253
rect 52790 53201 52948 53253
rect 53000 53201 53159 53253
rect 53211 53201 53371 53253
rect 53423 53201 53582 53253
rect 53634 53201 53792 53253
rect 53844 53201 54003 53253
rect 54055 53201 54214 53253
rect 54266 53201 54355 53253
rect 51796 53047 52106 53087
rect 51796 52995 51835 53047
rect 51887 52995 52015 53047
rect 52067 52995 52106 53047
rect 50099 52763 50300 52815
rect 50352 52763 50511 52815
rect 50563 52763 50722 52815
rect 50774 52763 50913 52815
rect 50099 52353 50913 52763
rect 51034 52795 51344 52868
rect 51034 52739 51071 52795
rect 51127 52739 51251 52795
rect 51307 52739 51344 52795
rect 51034 52577 51344 52739
rect 51034 52525 51073 52577
rect 51125 52525 51253 52577
rect 51305 52525 51344 52577
rect 51034 52484 51344 52525
rect 51796 52795 52106 52995
rect 51796 52739 51833 52795
rect 51889 52739 52013 52795
rect 52069 52739 52106 52795
rect 51796 52584 52106 52739
rect 51796 52532 51835 52584
rect 51887 52532 52015 52584
rect 52067 52532 52106 52584
rect 51796 52491 52106 52532
rect 50099 52301 50346 52353
rect 50398 52301 50557 52353
rect 50609 52301 50768 52353
rect 50820 52301 50913 52353
rect 50099 51891 50913 52301
rect 52227 52355 54355 53201
rect 52227 52299 52314 52355
rect 52370 52299 52525 52355
rect 52581 52299 52736 52355
rect 52792 52299 52946 52355
rect 53002 52299 53157 52355
rect 53213 52299 53369 52355
rect 53425 52299 53580 52355
rect 53636 52299 53790 52355
rect 53846 52299 54001 52355
rect 54057 52299 54212 52355
rect 54268 52299 54355 52355
rect 50099 51839 50300 51891
rect 50352 51839 50511 51891
rect 50563 51839 50722 51891
rect 50774 51839 50913 51891
rect 50099 51455 50913 51839
rect 51034 52129 51344 52170
rect 51034 52077 51073 52129
rect 51125 52077 51253 52129
rect 51305 52077 51344 52129
rect 51034 51915 51344 52077
rect 51034 51859 51071 51915
rect 51127 51859 51251 51915
rect 51307 51859 51344 51915
rect 51034 51786 51344 51859
rect 51796 52122 52106 52163
rect 51796 52070 51835 52122
rect 51887 52070 52015 52122
rect 52067 52070 52106 52122
rect 51796 51915 52106 52070
rect 51796 51859 51833 51915
rect 51889 51859 52013 51915
rect 52069 51859 52106 51915
rect 51796 51659 52106 51859
rect 51796 51607 51835 51659
rect 51887 51607 52015 51659
rect 52067 51607 52106 51659
rect 51796 51567 52106 51607
rect 50099 51453 50161 51455
rect 50217 51453 50372 51455
rect 50099 51401 50138 51453
rect 50217 51401 50318 51453
rect 50370 51401 50372 51453
rect 50099 51399 50161 51401
rect 50217 51399 50372 51401
rect 50428 51399 50584 51455
rect 50640 51399 50795 51455
rect 50851 51399 50913 51455
rect 50099 51015 50913 51399
rect 52227 51453 54355 52299
rect 52227 51401 52316 51453
rect 52368 51401 52527 51453
rect 52579 51401 52738 51453
rect 52790 51401 52948 51453
rect 53000 51401 53159 51453
rect 53211 51401 53371 51453
rect 53423 51401 53582 51453
rect 53634 51401 53792 51453
rect 53844 51401 54003 51453
rect 54055 51401 54214 51453
rect 54266 51401 54355 51453
rect 51796 51247 52106 51287
rect 51796 51195 51835 51247
rect 51887 51195 52015 51247
rect 52067 51195 52106 51247
rect 50099 50963 50300 51015
rect 50352 50963 50511 51015
rect 50563 50963 50722 51015
rect 50774 50963 50913 51015
rect 50099 50553 50913 50963
rect 51034 50995 51344 51068
rect 51034 50939 51071 50995
rect 51127 50939 51251 50995
rect 51307 50939 51344 50995
rect 51034 50777 51344 50939
rect 51034 50725 51073 50777
rect 51125 50725 51253 50777
rect 51305 50725 51344 50777
rect 51034 50684 51344 50725
rect 51796 50995 52106 51195
rect 51796 50939 51833 50995
rect 51889 50939 52013 50995
rect 52069 50939 52106 50995
rect 51796 50784 52106 50939
rect 51796 50732 51835 50784
rect 51887 50732 52015 50784
rect 52067 50732 52106 50784
rect 51796 50691 52106 50732
rect 50099 50501 50346 50553
rect 50398 50501 50557 50553
rect 50609 50501 50768 50553
rect 50820 50501 50913 50553
rect 50099 50091 50913 50501
rect 52227 50555 54355 51401
rect 52227 50499 52314 50555
rect 52370 50499 52525 50555
rect 52581 50499 52736 50555
rect 52792 50499 52946 50555
rect 53002 50499 53157 50555
rect 53213 50499 53369 50555
rect 53425 50499 53580 50555
rect 53636 50499 53790 50555
rect 53846 50499 54001 50555
rect 54057 50499 54212 50555
rect 54268 50499 54355 50555
rect 50099 50039 50300 50091
rect 50352 50039 50511 50091
rect 50563 50039 50722 50091
rect 50774 50039 50913 50091
rect 50099 49655 50913 50039
rect 51034 50329 51344 50370
rect 51034 50277 51073 50329
rect 51125 50277 51253 50329
rect 51305 50277 51344 50329
rect 51034 50115 51344 50277
rect 51034 50059 51071 50115
rect 51127 50059 51251 50115
rect 51307 50059 51344 50115
rect 51034 49986 51344 50059
rect 51796 50322 52106 50363
rect 51796 50270 51835 50322
rect 51887 50270 52015 50322
rect 52067 50270 52106 50322
rect 51796 50115 52106 50270
rect 51796 50059 51833 50115
rect 51889 50059 52013 50115
rect 52069 50059 52106 50115
rect 51796 49859 52106 50059
rect 51796 49807 51835 49859
rect 51887 49807 52015 49859
rect 52067 49807 52106 49859
rect 51796 49767 52106 49807
rect 50099 49653 50161 49655
rect 50217 49653 50372 49655
rect 50099 49601 50138 49653
rect 50217 49601 50318 49653
rect 50370 49601 50372 49653
rect 50099 49599 50161 49601
rect 50217 49599 50372 49601
rect 50428 49599 50584 49655
rect 50640 49599 50795 49655
rect 50851 49599 50913 49655
rect 50099 49215 50913 49599
rect 52227 49653 54355 50499
rect 52227 49601 52316 49653
rect 52368 49601 52527 49653
rect 52579 49601 52738 49653
rect 52790 49601 52948 49653
rect 53000 49601 53159 49653
rect 53211 49601 53371 49653
rect 53423 49601 53582 49653
rect 53634 49601 53792 49653
rect 53844 49601 54003 49653
rect 54055 49601 54214 49653
rect 54266 49601 54355 49653
rect 51796 49447 52106 49487
rect 51796 49395 51835 49447
rect 51887 49395 52015 49447
rect 52067 49395 52106 49447
rect 50099 49163 50300 49215
rect 50352 49163 50511 49215
rect 50563 49163 50722 49215
rect 50774 49163 50913 49215
rect 50099 48753 50913 49163
rect 51034 49195 51344 49268
rect 51034 49139 51071 49195
rect 51127 49139 51251 49195
rect 51307 49139 51344 49195
rect 51034 48977 51344 49139
rect 51034 48925 51073 48977
rect 51125 48925 51253 48977
rect 51305 48925 51344 48977
rect 51034 48884 51344 48925
rect 51796 49195 52106 49395
rect 51796 49139 51833 49195
rect 51889 49139 52013 49195
rect 52069 49139 52106 49195
rect 51796 48984 52106 49139
rect 51796 48932 51835 48984
rect 51887 48932 52015 48984
rect 52067 48932 52106 48984
rect 51796 48891 52106 48932
rect 50099 48701 50346 48753
rect 50398 48701 50557 48753
rect 50609 48701 50768 48753
rect 50820 48701 50913 48753
rect 50099 48291 50913 48701
rect 52227 48755 54355 49601
rect 52227 48699 52314 48755
rect 52370 48699 52525 48755
rect 52581 48699 52736 48755
rect 52792 48699 52946 48755
rect 53002 48699 53157 48755
rect 53213 48699 53369 48755
rect 53425 48699 53580 48755
rect 53636 48699 53790 48755
rect 53846 48699 54001 48755
rect 54057 48699 54212 48755
rect 54268 48699 54355 48755
rect 50099 48239 50300 48291
rect 50352 48239 50511 48291
rect 50563 48239 50722 48291
rect 50774 48239 50913 48291
rect 50099 47855 50913 48239
rect 51034 48529 51344 48570
rect 51034 48477 51073 48529
rect 51125 48477 51253 48529
rect 51305 48477 51344 48529
rect 51034 48315 51344 48477
rect 51034 48259 51071 48315
rect 51127 48259 51251 48315
rect 51307 48259 51344 48315
rect 51034 48186 51344 48259
rect 51796 48522 52106 48563
rect 51796 48470 51835 48522
rect 51887 48470 52015 48522
rect 52067 48470 52106 48522
rect 51796 48315 52106 48470
rect 51796 48259 51833 48315
rect 51889 48259 52013 48315
rect 52069 48259 52106 48315
rect 51796 48059 52106 48259
rect 51796 48007 51835 48059
rect 51887 48007 52015 48059
rect 52067 48007 52106 48059
rect 51796 47967 52106 48007
rect 50099 47853 50161 47855
rect 50217 47853 50372 47855
rect 50099 47801 50138 47853
rect 50217 47801 50318 47853
rect 50370 47801 50372 47853
rect 50099 47799 50161 47801
rect 50217 47799 50372 47801
rect 50428 47799 50584 47855
rect 50640 47799 50795 47855
rect 50851 47799 50913 47855
rect 50099 47415 50913 47799
rect 52227 47853 54355 48699
rect 52227 47801 52316 47853
rect 52368 47801 52527 47853
rect 52579 47801 52738 47853
rect 52790 47801 52948 47853
rect 53000 47801 53159 47853
rect 53211 47801 53371 47853
rect 53423 47801 53582 47853
rect 53634 47801 53792 47853
rect 53844 47801 54003 47853
rect 54055 47801 54214 47853
rect 54266 47801 54355 47853
rect 51796 47647 52106 47687
rect 51796 47595 51835 47647
rect 51887 47595 52015 47647
rect 52067 47595 52106 47647
rect 50099 47363 50300 47415
rect 50352 47363 50511 47415
rect 50563 47363 50722 47415
rect 50774 47363 50913 47415
rect 50099 46953 50913 47363
rect 51034 47395 51344 47468
rect 51034 47339 51071 47395
rect 51127 47339 51251 47395
rect 51307 47339 51344 47395
rect 51034 47177 51344 47339
rect 51034 47125 51073 47177
rect 51125 47125 51253 47177
rect 51305 47125 51344 47177
rect 51034 47084 51344 47125
rect 51796 47395 52106 47595
rect 51796 47339 51833 47395
rect 51889 47339 52013 47395
rect 52069 47339 52106 47395
rect 51796 47184 52106 47339
rect 51796 47132 51835 47184
rect 51887 47132 52015 47184
rect 52067 47132 52106 47184
rect 51796 47091 52106 47132
rect 50099 46901 50346 46953
rect 50398 46901 50557 46953
rect 50609 46901 50768 46953
rect 50820 46901 50913 46953
rect 50099 46491 50913 46901
rect 52227 46955 54355 47801
rect 52227 46899 52314 46955
rect 52370 46899 52525 46955
rect 52581 46899 52736 46955
rect 52792 46899 52946 46955
rect 53002 46899 53157 46955
rect 53213 46899 53369 46955
rect 53425 46899 53580 46955
rect 53636 46899 53790 46955
rect 53846 46899 54001 46955
rect 54057 46899 54212 46955
rect 54268 46899 54355 46955
rect 50099 46439 50300 46491
rect 50352 46439 50511 46491
rect 50563 46439 50722 46491
rect 50774 46439 50913 46491
rect 50099 46055 50913 46439
rect 51034 46729 51344 46770
rect 51034 46677 51073 46729
rect 51125 46677 51253 46729
rect 51305 46677 51344 46729
rect 51034 46515 51344 46677
rect 51034 46459 51071 46515
rect 51127 46459 51251 46515
rect 51307 46459 51344 46515
rect 51034 46386 51344 46459
rect 51796 46722 52106 46763
rect 51796 46670 51835 46722
rect 51887 46670 52015 46722
rect 52067 46670 52106 46722
rect 51796 46515 52106 46670
rect 51796 46459 51833 46515
rect 51889 46459 52013 46515
rect 52069 46459 52106 46515
rect 51796 46259 52106 46459
rect 51796 46207 51835 46259
rect 51887 46207 52015 46259
rect 52067 46207 52106 46259
rect 51796 46167 52106 46207
rect 50099 46053 50161 46055
rect 50217 46053 50372 46055
rect 50099 46001 50138 46053
rect 50217 46001 50318 46053
rect 50370 46001 50372 46053
rect 50099 45999 50161 46001
rect 50217 45999 50372 46001
rect 50428 45999 50584 46055
rect 50640 45999 50795 46055
rect 50851 45999 50913 46055
rect 50099 45615 50913 45999
rect 52227 46053 54355 46899
rect 52227 46001 52316 46053
rect 52368 46001 52527 46053
rect 52579 46001 52738 46053
rect 52790 46001 52948 46053
rect 53000 46001 53159 46053
rect 53211 46001 53371 46053
rect 53423 46001 53582 46053
rect 53634 46001 53792 46053
rect 53844 46001 54003 46053
rect 54055 46001 54214 46053
rect 54266 46001 54355 46053
rect 51796 45847 52106 45887
rect 51796 45795 51835 45847
rect 51887 45795 52015 45847
rect 52067 45795 52106 45847
rect 50099 45563 50300 45615
rect 50352 45563 50511 45615
rect 50563 45563 50722 45615
rect 50774 45563 50913 45615
rect 50099 45153 50913 45563
rect 51034 45595 51344 45668
rect 51034 45539 51071 45595
rect 51127 45539 51251 45595
rect 51307 45539 51344 45595
rect 51034 45377 51344 45539
rect 51034 45325 51073 45377
rect 51125 45325 51253 45377
rect 51305 45325 51344 45377
rect 51034 45284 51344 45325
rect 51796 45595 52106 45795
rect 51796 45539 51833 45595
rect 51889 45539 52013 45595
rect 52069 45539 52106 45595
rect 51796 45384 52106 45539
rect 51796 45332 51835 45384
rect 51887 45332 52015 45384
rect 52067 45332 52106 45384
rect 51796 45291 52106 45332
rect 50099 45101 50346 45153
rect 50398 45101 50557 45153
rect 50609 45101 50768 45153
rect 50820 45101 50913 45153
rect 50099 44691 50913 45101
rect 52227 45155 54355 46001
rect 52227 45099 52314 45155
rect 52370 45099 52525 45155
rect 52581 45099 52736 45155
rect 52792 45099 52946 45155
rect 53002 45099 53157 45155
rect 53213 45099 53369 45155
rect 53425 45099 53580 45155
rect 53636 45099 53790 45155
rect 53846 45099 54001 45155
rect 54057 45099 54212 45155
rect 54268 45099 54355 45155
rect 50099 44639 50300 44691
rect 50352 44639 50511 44691
rect 50563 44639 50722 44691
rect 50774 44639 50913 44691
rect 50099 44255 50913 44639
rect 51034 44929 51344 44970
rect 51034 44877 51073 44929
rect 51125 44877 51253 44929
rect 51305 44877 51344 44929
rect 51034 44715 51344 44877
rect 51034 44659 51071 44715
rect 51127 44659 51251 44715
rect 51307 44659 51344 44715
rect 51034 44586 51344 44659
rect 51796 44922 52106 44963
rect 51796 44870 51835 44922
rect 51887 44870 52015 44922
rect 52067 44870 52106 44922
rect 51796 44715 52106 44870
rect 51796 44659 51833 44715
rect 51889 44659 52013 44715
rect 52069 44659 52106 44715
rect 51796 44459 52106 44659
rect 51796 44407 51835 44459
rect 51887 44407 52015 44459
rect 52067 44407 52106 44459
rect 51796 44367 52106 44407
rect 50099 44253 50161 44255
rect 50217 44253 50372 44255
rect 50099 44201 50138 44253
rect 50217 44201 50318 44253
rect 50370 44201 50372 44253
rect 50099 44199 50161 44201
rect 50217 44199 50372 44201
rect 50428 44199 50584 44255
rect 50640 44199 50795 44255
rect 50851 44199 50913 44255
rect 50099 43815 50913 44199
rect 52227 44253 54355 45099
rect 52227 44201 52316 44253
rect 52368 44201 52527 44253
rect 52579 44201 52738 44253
rect 52790 44201 52948 44253
rect 53000 44201 53159 44253
rect 53211 44201 53371 44253
rect 53423 44201 53582 44253
rect 53634 44201 53792 44253
rect 53844 44201 54003 44253
rect 54055 44201 54214 44253
rect 54266 44201 54355 44253
rect 51796 44047 52106 44087
rect 51796 43995 51835 44047
rect 51887 43995 52015 44047
rect 52067 43995 52106 44047
rect 50099 43763 50300 43815
rect 50352 43763 50511 43815
rect 50563 43763 50722 43815
rect 50774 43763 50913 43815
rect 50099 43353 50913 43763
rect 51034 43795 51344 43868
rect 51034 43739 51071 43795
rect 51127 43739 51251 43795
rect 51307 43739 51344 43795
rect 51034 43577 51344 43739
rect 51034 43525 51073 43577
rect 51125 43525 51253 43577
rect 51305 43525 51344 43577
rect 51034 43484 51344 43525
rect 51796 43795 52106 43995
rect 51796 43739 51833 43795
rect 51889 43739 52013 43795
rect 52069 43739 52106 43795
rect 51796 43584 52106 43739
rect 51796 43532 51835 43584
rect 51887 43532 52015 43584
rect 52067 43532 52106 43584
rect 51796 43491 52106 43532
rect 50099 43301 50346 43353
rect 50398 43301 50557 43353
rect 50609 43301 50768 43353
rect 50820 43301 50913 43353
rect 50099 42891 50913 43301
rect 52227 43355 54355 44201
rect 52227 43299 52314 43355
rect 52370 43299 52525 43355
rect 52581 43299 52736 43355
rect 52792 43299 52946 43355
rect 53002 43299 53157 43355
rect 53213 43299 53369 43355
rect 53425 43299 53580 43355
rect 53636 43299 53790 43355
rect 53846 43299 54001 43355
rect 54057 43299 54212 43355
rect 54268 43299 54355 43355
rect 50099 42839 50300 42891
rect 50352 42839 50511 42891
rect 50563 42839 50722 42891
rect 50774 42839 50913 42891
rect 50099 42455 50913 42839
rect 51034 43129 51344 43170
rect 51034 43077 51073 43129
rect 51125 43077 51253 43129
rect 51305 43077 51344 43129
rect 51034 42915 51344 43077
rect 51034 42859 51071 42915
rect 51127 42859 51251 42915
rect 51307 42859 51344 42915
rect 51034 42786 51344 42859
rect 51796 43122 52106 43163
rect 51796 43070 51835 43122
rect 51887 43070 52015 43122
rect 52067 43070 52106 43122
rect 51796 42915 52106 43070
rect 51796 42859 51833 42915
rect 51889 42859 52013 42915
rect 52069 42859 52106 42915
rect 51796 42659 52106 42859
rect 51796 42607 51835 42659
rect 51887 42607 52015 42659
rect 52067 42607 52106 42659
rect 51796 42567 52106 42607
rect 50099 42453 50161 42455
rect 50217 42453 50372 42455
rect 50099 42401 50138 42453
rect 50217 42401 50318 42453
rect 50370 42401 50372 42453
rect 50099 42399 50161 42401
rect 50217 42399 50372 42401
rect 50428 42399 50584 42455
rect 50640 42399 50795 42455
rect 50851 42399 50913 42455
rect 50099 42015 50913 42399
rect 52227 42453 54355 43299
rect 52227 42401 52316 42453
rect 52368 42401 52527 42453
rect 52579 42401 52738 42453
rect 52790 42401 52948 42453
rect 53000 42401 53159 42453
rect 53211 42401 53371 42453
rect 53423 42401 53582 42453
rect 53634 42401 53792 42453
rect 53844 42401 54003 42453
rect 54055 42401 54214 42453
rect 54266 42401 54355 42453
rect 51796 42247 52106 42287
rect 51796 42195 51835 42247
rect 51887 42195 52015 42247
rect 52067 42195 52106 42247
rect 50099 41963 50300 42015
rect 50352 41963 50511 42015
rect 50563 41963 50722 42015
rect 50774 41963 50913 42015
rect 50099 41553 50913 41963
rect 51034 41995 51344 42068
rect 51034 41939 51071 41995
rect 51127 41939 51251 41995
rect 51307 41939 51344 41995
rect 51034 41777 51344 41939
rect 51034 41725 51073 41777
rect 51125 41725 51253 41777
rect 51305 41725 51344 41777
rect 51034 41684 51344 41725
rect 51796 41995 52106 42195
rect 51796 41939 51833 41995
rect 51889 41939 52013 41995
rect 52069 41939 52106 41995
rect 51796 41784 52106 41939
rect 51796 41732 51835 41784
rect 51887 41732 52015 41784
rect 52067 41732 52106 41784
rect 51796 41691 52106 41732
rect 50099 41501 50346 41553
rect 50398 41501 50557 41553
rect 50609 41501 50768 41553
rect 50820 41501 50913 41553
rect 50099 41091 50913 41501
rect 52227 41555 54355 42401
rect 52227 41499 52314 41555
rect 52370 41499 52525 41555
rect 52581 41499 52736 41555
rect 52792 41499 52946 41555
rect 53002 41499 53157 41555
rect 53213 41499 53369 41555
rect 53425 41499 53580 41555
rect 53636 41499 53790 41555
rect 53846 41499 54001 41555
rect 54057 41499 54212 41555
rect 54268 41499 54355 41555
rect 50099 41039 50300 41091
rect 50352 41039 50511 41091
rect 50563 41039 50722 41091
rect 50774 41039 50913 41091
rect 50099 40655 50913 41039
rect 51034 41329 51344 41370
rect 51034 41277 51073 41329
rect 51125 41277 51253 41329
rect 51305 41277 51344 41329
rect 51034 41115 51344 41277
rect 51034 41059 51071 41115
rect 51127 41059 51251 41115
rect 51307 41059 51344 41115
rect 51034 40986 51344 41059
rect 51796 41322 52106 41363
rect 51796 41270 51835 41322
rect 51887 41270 52015 41322
rect 52067 41270 52106 41322
rect 51796 41115 52106 41270
rect 51796 41059 51833 41115
rect 51889 41059 52013 41115
rect 52069 41059 52106 41115
rect 51796 40859 52106 41059
rect 51796 40807 51835 40859
rect 51887 40807 52015 40859
rect 52067 40807 52106 40859
rect 51796 40767 52106 40807
rect 50099 40653 50161 40655
rect 50217 40653 50372 40655
rect 50099 40601 50138 40653
rect 50217 40601 50318 40653
rect 50370 40601 50372 40653
rect 50099 40599 50161 40601
rect 50217 40599 50372 40601
rect 50428 40599 50584 40655
rect 50640 40599 50795 40655
rect 50851 40599 50913 40655
rect 50099 40215 50913 40599
rect 52227 40653 54355 41499
rect 52227 40601 52316 40653
rect 52368 40601 52527 40653
rect 52579 40601 52738 40653
rect 52790 40601 52948 40653
rect 53000 40601 53159 40653
rect 53211 40601 53371 40653
rect 53423 40601 53582 40653
rect 53634 40601 53792 40653
rect 53844 40601 54003 40653
rect 54055 40601 54214 40653
rect 54266 40601 54355 40653
rect 51796 40447 52106 40487
rect 51796 40395 51835 40447
rect 51887 40395 52015 40447
rect 52067 40395 52106 40447
rect 50099 40163 50300 40215
rect 50352 40163 50511 40215
rect 50563 40163 50722 40215
rect 50774 40163 50913 40215
rect 50099 39753 50913 40163
rect 51034 40195 51344 40268
rect 51034 40139 51071 40195
rect 51127 40139 51251 40195
rect 51307 40139 51344 40195
rect 51034 39977 51344 40139
rect 51034 39925 51073 39977
rect 51125 39925 51253 39977
rect 51305 39925 51344 39977
rect 51034 39884 51344 39925
rect 51796 40195 52106 40395
rect 51796 40139 51833 40195
rect 51889 40139 52013 40195
rect 52069 40139 52106 40195
rect 51796 39984 52106 40139
rect 51796 39932 51835 39984
rect 51887 39932 52015 39984
rect 52067 39932 52106 39984
rect 51796 39891 52106 39932
rect 50099 39701 50346 39753
rect 50398 39701 50557 39753
rect 50609 39701 50768 39753
rect 50820 39701 50913 39753
rect 50099 39291 50913 39701
rect 52227 39755 54355 40601
rect 52227 39699 52314 39755
rect 52370 39699 52525 39755
rect 52581 39699 52736 39755
rect 52792 39699 52946 39755
rect 53002 39699 53157 39755
rect 53213 39699 53369 39755
rect 53425 39699 53580 39755
rect 53636 39699 53790 39755
rect 53846 39699 54001 39755
rect 54057 39699 54212 39755
rect 54268 39699 54355 39755
rect 50099 39239 50300 39291
rect 50352 39239 50511 39291
rect 50563 39239 50722 39291
rect 50774 39239 50913 39291
rect 50099 38855 50913 39239
rect 51034 39529 51344 39570
rect 51034 39477 51073 39529
rect 51125 39477 51253 39529
rect 51305 39477 51344 39529
rect 51034 39315 51344 39477
rect 51034 39259 51071 39315
rect 51127 39259 51251 39315
rect 51307 39259 51344 39315
rect 51034 39186 51344 39259
rect 51796 39522 52106 39563
rect 51796 39470 51835 39522
rect 51887 39470 52015 39522
rect 52067 39470 52106 39522
rect 51796 39315 52106 39470
rect 51796 39259 51833 39315
rect 51889 39259 52013 39315
rect 52069 39259 52106 39315
rect 51796 39059 52106 39259
rect 51796 39007 51835 39059
rect 51887 39007 52015 39059
rect 52067 39007 52106 39059
rect 51796 38967 52106 39007
rect 50099 38853 50161 38855
rect 50217 38853 50372 38855
rect 50099 38801 50138 38853
rect 50217 38801 50318 38853
rect 50370 38801 50372 38853
rect 50099 38799 50161 38801
rect 50217 38799 50372 38801
rect 50428 38799 50584 38855
rect 50640 38799 50795 38855
rect 50851 38799 50913 38855
rect 50099 38415 50913 38799
rect 52227 38853 54355 39699
rect 52227 38801 52316 38853
rect 52368 38801 52527 38853
rect 52579 38801 52738 38853
rect 52790 38801 52948 38853
rect 53000 38801 53159 38853
rect 53211 38801 53371 38853
rect 53423 38801 53582 38853
rect 53634 38801 53792 38853
rect 53844 38801 54003 38853
rect 54055 38801 54214 38853
rect 54266 38801 54355 38853
rect 51796 38647 52106 38687
rect 51796 38595 51835 38647
rect 51887 38595 52015 38647
rect 52067 38595 52106 38647
rect 50099 38363 50300 38415
rect 50352 38363 50511 38415
rect 50563 38363 50722 38415
rect 50774 38363 50913 38415
rect 50099 37953 50913 38363
rect 51034 38395 51344 38468
rect 51034 38339 51071 38395
rect 51127 38339 51251 38395
rect 51307 38339 51344 38395
rect 51034 38177 51344 38339
rect 51034 38125 51073 38177
rect 51125 38125 51253 38177
rect 51305 38125 51344 38177
rect 51034 38084 51344 38125
rect 51796 38395 52106 38595
rect 51796 38339 51833 38395
rect 51889 38339 52013 38395
rect 52069 38339 52106 38395
rect 51796 38184 52106 38339
rect 51796 38132 51835 38184
rect 51887 38132 52015 38184
rect 52067 38132 52106 38184
rect 51796 38091 52106 38132
rect 50099 37901 50346 37953
rect 50398 37901 50557 37953
rect 50609 37901 50768 37953
rect 50820 37901 50913 37953
rect 50099 37491 50913 37901
rect 52227 37955 54355 38801
rect 52227 37899 52314 37955
rect 52370 37899 52525 37955
rect 52581 37899 52736 37955
rect 52792 37899 52946 37955
rect 53002 37899 53157 37955
rect 53213 37899 53369 37955
rect 53425 37899 53580 37955
rect 53636 37899 53790 37955
rect 53846 37899 54001 37955
rect 54057 37899 54212 37955
rect 54268 37899 54355 37955
rect 50099 37439 50300 37491
rect 50352 37439 50511 37491
rect 50563 37439 50722 37491
rect 50774 37439 50913 37491
rect 50099 37055 50913 37439
rect 51034 37729 51344 37770
rect 51034 37677 51073 37729
rect 51125 37677 51253 37729
rect 51305 37677 51344 37729
rect 51034 37515 51344 37677
rect 51034 37459 51071 37515
rect 51127 37459 51251 37515
rect 51307 37459 51344 37515
rect 51034 37386 51344 37459
rect 51796 37722 52106 37763
rect 51796 37670 51835 37722
rect 51887 37670 52015 37722
rect 52067 37670 52106 37722
rect 51796 37515 52106 37670
rect 51796 37459 51833 37515
rect 51889 37459 52013 37515
rect 52069 37459 52106 37515
rect 51796 37259 52106 37459
rect 51796 37207 51835 37259
rect 51887 37207 52015 37259
rect 52067 37207 52106 37259
rect 51796 37167 52106 37207
rect 50099 37053 50161 37055
rect 50217 37053 50372 37055
rect 50099 37001 50138 37053
rect 50217 37001 50318 37053
rect 50370 37001 50372 37053
rect 50099 36999 50161 37001
rect 50217 36999 50372 37001
rect 50428 36999 50584 37055
rect 50640 36999 50795 37055
rect 50851 36999 50913 37055
rect 50099 36615 50913 36999
rect 52227 37053 54355 37899
rect 52227 37001 52316 37053
rect 52368 37001 52527 37053
rect 52579 37001 52738 37053
rect 52790 37001 52948 37053
rect 53000 37001 53159 37053
rect 53211 37001 53371 37053
rect 53423 37001 53582 37053
rect 53634 37001 53792 37053
rect 53844 37001 54003 37053
rect 54055 37001 54214 37053
rect 54266 37001 54355 37053
rect 51796 36847 52106 36887
rect 51796 36795 51835 36847
rect 51887 36795 52015 36847
rect 52067 36795 52106 36847
rect 50099 36563 50300 36615
rect 50352 36563 50511 36615
rect 50563 36563 50722 36615
rect 50774 36563 50913 36615
rect 50099 36153 50913 36563
rect 51034 36595 51344 36668
rect 51034 36539 51071 36595
rect 51127 36539 51251 36595
rect 51307 36539 51344 36595
rect 51034 36377 51344 36539
rect 51034 36325 51073 36377
rect 51125 36325 51253 36377
rect 51305 36325 51344 36377
rect 51034 36284 51344 36325
rect 51796 36595 52106 36795
rect 51796 36539 51833 36595
rect 51889 36539 52013 36595
rect 52069 36539 52106 36595
rect 51796 36384 52106 36539
rect 51796 36332 51835 36384
rect 51887 36332 52015 36384
rect 52067 36332 52106 36384
rect 51796 36291 52106 36332
rect 50099 36101 50346 36153
rect 50398 36101 50557 36153
rect 50609 36101 50768 36153
rect 50820 36101 50913 36153
rect 50099 35976 50913 36101
rect 52227 36155 54355 37001
rect 52227 36099 52314 36155
rect 52370 36099 52525 36155
rect 52581 36099 52736 36155
rect 52792 36099 52946 36155
rect 53002 36099 53157 36155
rect 53213 36099 53369 36155
rect 53425 36099 53580 36155
rect 53636 36099 53790 36155
rect 53846 36099 54001 36155
rect 54057 36099 54212 36155
rect 54268 36099 54355 36155
rect 52227 35976 54355 36099
rect 54758 64955 55638 65801
rect 55977 65855 57371 65894
rect 55977 65799 56013 65855
rect 56069 65799 56224 65855
rect 56280 65799 56435 65855
rect 56491 65799 56646 65855
rect 56702 65799 56857 65855
rect 56913 65799 57068 65855
rect 57124 65799 57279 65855
rect 57335 65799 57371 65855
rect 55977 65760 57371 65799
rect 54758 64899 54853 64955
rect 54909 64899 55064 64955
rect 55120 64899 55276 64955
rect 55332 64899 55487 64955
rect 55543 64899 55638 64955
rect 54758 64053 55638 64899
rect 54758 64001 54855 64053
rect 54907 64001 55066 64053
rect 55118 64001 55278 64053
rect 55330 64001 55489 64053
rect 55541 64001 55638 64053
rect 54758 63155 55638 64001
rect 55977 64055 57371 64094
rect 55977 63999 56013 64055
rect 56069 63999 56224 64055
rect 56280 63999 56435 64055
rect 56491 63999 56646 64055
rect 56702 63999 56857 64055
rect 56913 63999 57068 64055
rect 57124 63999 57279 64055
rect 57335 63999 57371 64055
rect 55977 63960 57371 63999
rect 54758 63099 54853 63155
rect 54909 63099 55064 63155
rect 55120 63099 55276 63155
rect 55332 63099 55487 63155
rect 55543 63099 55638 63155
rect 54758 62253 55638 63099
rect 54758 62201 54855 62253
rect 54907 62201 55066 62253
rect 55118 62201 55278 62253
rect 55330 62201 55489 62253
rect 55541 62201 55638 62253
rect 54758 61355 55638 62201
rect 55977 62255 57371 62294
rect 55977 62199 56013 62255
rect 56069 62199 56224 62255
rect 56280 62199 56435 62255
rect 56491 62199 56646 62255
rect 56702 62199 56857 62255
rect 56913 62199 57068 62255
rect 57124 62199 57279 62255
rect 57335 62199 57371 62255
rect 55977 62160 57371 62199
rect 54758 61299 54853 61355
rect 54909 61299 55064 61355
rect 55120 61299 55276 61355
rect 55332 61299 55487 61355
rect 55543 61299 55638 61355
rect 54758 60453 55638 61299
rect 54758 60401 54855 60453
rect 54907 60401 55066 60453
rect 55118 60401 55278 60453
rect 55330 60401 55489 60453
rect 55541 60401 55638 60453
rect 54758 59555 55638 60401
rect 55977 60455 57371 60494
rect 55977 60399 56013 60455
rect 56069 60399 56224 60455
rect 56280 60399 56435 60455
rect 56491 60399 56646 60455
rect 56702 60399 56857 60455
rect 56913 60399 57068 60455
rect 57124 60399 57279 60455
rect 57335 60399 57371 60455
rect 55977 60360 57371 60399
rect 54758 59499 54853 59555
rect 54909 59499 55064 59555
rect 55120 59499 55276 59555
rect 55332 59499 55487 59555
rect 55543 59499 55638 59555
rect 54758 58653 55638 59499
rect 54758 58601 54855 58653
rect 54907 58601 55066 58653
rect 55118 58601 55278 58653
rect 55330 58601 55489 58653
rect 55541 58601 55638 58653
rect 54758 57755 55638 58601
rect 55977 58655 57371 58694
rect 55977 58599 56013 58655
rect 56069 58599 56224 58655
rect 56280 58599 56435 58655
rect 56491 58599 56646 58655
rect 56702 58599 56857 58655
rect 56913 58599 57068 58655
rect 57124 58599 57279 58655
rect 57335 58599 57371 58655
rect 55977 58560 57371 58599
rect 54758 57699 54853 57755
rect 54909 57699 55064 57755
rect 55120 57699 55276 57755
rect 55332 57699 55487 57755
rect 55543 57699 55638 57755
rect 54758 56853 55638 57699
rect 54758 56801 54855 56853
rect 54907 56801 55066 56853
rect 55118 56801 55278 56853
rect 55330 56801 55489 56853
rect 55541 56801 55638 56853
rect 54758 55955 55638 56801
rect 55977 56855 57371 56894
rect 55977 56799 56013 56855
rect 56069 56799 56224 56855
rect 56280 56799 56435 56855
rect 56491 56799 56646 56855
rect 56702 56799 56857 56855
rect 56913 56799 57068 56855
rect 57124 56799 57279 56855
rect 57335 56799 57371 56855
rect 55977 56760 57371 56799
rect 54758 55899 54853 55955
rect 54909 55899 55064 55955
rect 55120 55899 55276 55955
rect 55332 55899 55487 55955
rect 55543 55899 55638 55955
rect 54758 55053 55638 55899
rect 54758 55001 54855 55053
rect 54907 55001 55066 55053
rect 55118 55001 55278 55053
rect 55330 55001 55489 55053
rect 55541 55001 55638 55053
rect 54758 54155 55638 55001
rect 55977 55055 57371 55094
rect 55977 54999 56013 55055
rect 56069 54999 56224 55055
rect 56280 54999 56435 55055
rect 56491 54999 56646 55055
rect 56702 54999 56857 55055
rect 56913 54999 57068 55055
rect 57124 54999 57279 55055
rect 57335 54999 57371 55055
rect 55977 54960 57371 54999
rect 54758 54099 54853 54155
rect 54909 54099 55064 54155
rect 55120 54099 55276 54155
rect 55332 54099 55487 54155
rect 55543 54099 55638 54155
rect 54758 53253 55638 54099
rect 54758 53201 54855 53253
rect 54907 53201 55066 53253
rect 55118 53201 55278 53253
rect 55330 53201 55489 53253
rect 55541 53201 55638 53253
rect 54758 52355 55638 53201
rect 55977 53255 57371 53294
rect 55977 53199 56013 53255
rect 56069 53199 56224 53255
rect 56280 53199 56435 53255
rect 56491 53199 56646 53255
rect 56702 53199 56857 53255
rect 56913 53199 57068 53255
rect 57124 53199 57279 53255
rect 57335 53199 57371 53255
rect 55977 53160 57371 53199
rect 54758 52299 54853 52355
rect 54909 52299 55064 52355
rect 55120 52299 55276 52355
rect 55332 52299 55487 52355
rect 55543 52299 55638 52355
rect 54758 51453 55638 52299
rect 54758 51401 54855 51453
rect 54907 51401 55066 51453
rect 55118 51401 55278 51453
rect 55330 51401 55489 51453
rect 55541 51401 55638 51453
rect 54758 50555 55638 51401
rect 55977 51455 57371 51494
rect 55977 51399 56013 51455
rect 56069 51399 56224 51455
rect 56280 51399 56435 51455
rect 56491 51399 56646 51455
rect 56702 51399 56857 51455
rect 56913 51399 57068 51455
rect 57124 51399 57279 51455
rect 57335 51399 57371 51455
rect 55977 51360 57371 51399
rect 54758 50499 54853 50555
rect 54909 50499 55064 50555
rect 55120 50499 55276 50555
rect 55332 50499 55487 50555
rect 55543 50499 55638 50555
rect 54758 49653 55638 50499
rect 54758 49601 54855 49653
rect 54907 49601 55066 49653
rect 55118 49601 55278 49653
rect 55330 49601 55489 49653
rect 55541 49601 55638 49653
rect 54758 48755 55638 49601
rect 55977 49655 57371 49694
rect 55977 49599 56013 49655
rect 56069 49599 56224 49655
rect 56280 49599 56435 49655
rect 56491 49599 56646 49655
rect 56702 49599 56857 49655
rect 56913 49599 57068 49655
rect 57124 49599 57279 49655
rect 57335 49599 57371 49655
rect 55977 49560 57371 49599
rect 54758 48699 54853 48755
rect 54909 48699 55064 48755
rect 55120 48699 55276 48755
rect 55332 48699 55487 48755
rect 55543 48699 55638 48755
rect 54758 47853 55638 48699
rect 54758 47801 54855 47853
rect 54907 47801 55066 47853
rect 55118 47801 55278 47853
rect 55330 47801 55489 47853
rect 55541 47801 55638 47853
rect 54758 46955 55638 47801
rect 55977 47855 57371 47894
rect 55977 47799 56013 47855
rect 56069 47799 56224 47855
rect 56280 47799 56435 47855
rect 56491 47799 56646 47855
rect 56702 47799 56857 47855
rect 56913 47799 57068 47855
rect 57124 47799 57279 47855
rect 57335 47799 57371 47855
rect 55977 47760 57371 47799
rect 54758 46899 54853 46955
rect 54909 46899 55064 46955
rect 55120 46899 55276 46955
rect 55332 46899 55487 46955
rect 55543 46899 55638 46955
rect 54758 46053 55638 46899
rect 54758 46001 54855 46053
rect 54907 46001 55066 46053
rect 55118 46001 55278 46053
rect 55330 46001 55489 46053
rect 55541 46001 55638 46053
rect 54758 45155 55638 46001
rect 55977 46055 57371 46094
rect 55977 45999 56013 46055
rect 56069 45999 56224 46055
rect 56280 45999 56435 46055
rect 56491 45999 56646 46055
rect 56702 45999 56857 46055
rect 56913 45999 57068 46055
rect 57124 45999 57279 46055
rect 57335 45999 57371 46055
rect 55977 45960 57371 45999
rect 54758 45099 54853 45155
rect 54909 45099 55064 45155
rect 55120 45099 55276 45155
rect 55332 45099 55487 45155
rect 55543 45099 55638 45155
rect 54758 44253 55638 45099
rect 54758 44201 54855 44253
rect 54907 44201 55066 44253
rect 55118 44201 55278 44253
rect 55330 44201 55489 44253
rect 55541 44201 55638 44253
rect 54758 43355 55638 44201
rect 55977 44255 57371 44294
rect 55977 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 57371 44255
rect 55977 44160 57371 44199
rect 54758 43299 54853 43355
rect 54909 43299 55064 43355
rect 55120 43299 55276 43355
rect 55332 43299 55487 43355
rect 55543 43299 55638 43355
rect 54758 42453 55638 43299
rect 54758 42401 54855 42453
rect 54907 42401 55066 42453
rect 55118 42401 55278 42453
rect 55330 42401 55489 42453
rect 55541 42401 55638 42453
rect 54758 41555 55638 42401
rect 55977 42455 57371 42494
rect 55977 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 57371 42455
rect 55977 42360 57371 42399
rect 54758 41499 54853 41555
rect 54909 41499 55064 41555
rect 55120 41499 55276 41555
rect 55332 41499 55487 41555
rect 55543 41499 55638 41555
rect 54758 40653 55638 41499
rect 54758 40601 54855 40653
rect 54907 40601 55066 40653
rect 55118 40601 55278 40653
rect 55330 40601 55489 40653
rect 55541 40601 55638 40653
rect 54758 39755 55638 40601
rect 55977 40655 57371 40694
rect 55977 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 57371 40655
rect 55977 40560 57371 40599
rect 54758 39699 54853 39755
rect 54909 39699 55064 39755
rect 55120 39699 55276 39755
rect 55332 39699 55487 39755
rect 55543 39699 55638 39755
rect 54758 38853 55638 39699
rect 54758 38801 54855 38853
rect 54907 38801 55066 38853
rect 55118 38801 55278 38853
rect 55330 38801 55489 38853
rect 55541 38801 55638 38853
rect 54758 37955 55638 38801
rect 55977 38855 57371 38894
rect 55977 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 57371 38855
rect 55977 38760 57371 38799
rect 54758 37899 54853 37955
rect 54909 37899 55064 37955
rect 55120 37899 55276 37955
rect 55332 37899 55487 37955
rect 55543 37899 55638 37955
rect 54758 37053 55638 37899
rect 54758 37001 54855 37053
rect 54907 37001 55066 37053
rect 55118 37001 55278 37053
rect 55330 37001 55489 37053
rect 55541 37001 55638 37053
rect 54758 36155 55638 37001
rect 55977 37055 57371 37094
rect 55977 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 57371 37055
rect 55977 36960 57371 36999
rect 54758 36099 54853 36155
rect 54909 36099 55064 36155
rect 55120 36099 55276 36155
rect 55332 36099 55487 36155
rect 55543 36099 55638 36155
rect 54758 36027 55638 36099
rect 48157 35614 50120 35842
rect 47779 35278 49769 35507
rect 47402 34943 48486 35171
rect 47026 34607 48135 34836
rect 47913 33564 48135 34607
rect 48265 33576 48486 34943
rect 49547 33576 49769 35278
rect 49898 33576 50120 35614
rect 57909 34011 58351 66376
rect 57909 33955 57996 34011
rect 58052 33955 58208 34011
rect 58264 33955 58351 34011
rect 57909 33793 58351 33955
rect 57909 33737 57996 33793
rect 58052 33737 58208 33793
rect 58264 33737 58351 33793
rect 57909 33576 58351 33737
rect 57909 33520 57996 33576
rect 58052 33520 58208 33576
rect 58264 33520 58351 33576
rect 57295 33432 57736 33519
rect 57295 33380 57383 33432
rect 57435 33380 57595 33432
rect 57647 33380 57736 33432
rect 27387 33163 27476 33215
rect 27528 33163 27688 33215
rect 27740 33163 27828 33215
rect 27387 33141 27828 33163
rect 27387 33085 27474 33141
rect 27530 33085 27686 33141
rect 27742 33085 27828 33141
rect 27387 32997 27828 33085
rect 27387 32945 27476 32997
rect 27528 32945 27688 32997
rect 27740 32945 27828 32997
rect 27387 32923 27828 32945
rect 27387 32867 27474 32923
rect 27530 32867 27686 32923
rect 27742 32867 27828 32923
rect 27387 32779 27828 32867
rect 27387 32727 27476 32779
rect 27528 32727 27688 32779
rect 27740 32727 27828 32779
rect 27387 32705 27828 32727
rect 27387 32649 27474 32705
rect 27530 32649 27686 32705
rect 27742 32649 27828 32705
rect 27387 32562 27828 32649
rect 27387 32510 27476 32562
rect 27528 32510 27688 32562
rect 27740 32510 27828 32562
rect 27387 32487 27828 32510
rect 27387 32431 27474 32487
rect 27530 32431 27686 32487
rect 27742 32431 27828 32487
rect 27387 32344 27828 32431
rect 27387 32292 27476 32344
rect 27528 32292 27688 32344
rect 27740 32292 27828 32344
rect 27387 32127 27828 32292
rect 27387 32075 27476 32127
rect 27528 32075 27688 32127
rect 27740 32075 27828 32127
rect 27387 31909 27828 32075
rect 27387 31857 27476 31909
rect 27528 31857 27688 31909
rect 27740 31857 27828 31909
rect 27387 31691 27828 31857
rect 27387 31639 27476 31691
rect 27528 31639 27688 31691
rect 27740 31639 27828 31691
rect 27387 31474 27828 31639
rect 27387 31422 27476 31474
rect 27528 31422 27688 31474
rect 27740 31422 27828 31474
rect 27387 31256 27828 31422
rect 27387 31252 27476 31256
rect 27528 31252 27688 31256
rect 27740 31252 27828 31256
rect 27387 31196 27474 31252
rect 27530 31196 27686 31252
rect 27742 31196 27828 31252
rect 27387 31038 27828 31196
rect 27387 31034 27476 31038
rect 27528 31034 27688 31038
rect 27740 31034 27828 31038
rect 27387 30978 27474 31034
rect 27530 30978 27686 31034
rect 27742 30978 27828 31034
rect 27387 30821 27828 30978
rect 27387 30816 27476 30821
rect 27528 30816 27688 30821
rect 27740 30816 27828 30821
rect 27387 30760 27474 30816
rect 27530 30760 27686 30816
rect 27742 30760 27828 30816
rect 27387 30603 27828 30760
rect 27387 30598 27476 30603
rect 27528 30598 27688 30603
rect 27740 30598 27828 30603
rect 27387 30542 27474 30598
rect 27530 30542 27686 30598
rect 27742 30542 27828 30598
rect 27387 30386 27828 30542
rect 27387 30334 27476 30386
rect 27528 30334 27688 30386
rect 27740 30334 27828 30386
rect 27387 30168 27828 30334
rect 27387 30116 27476 30168
rect 27528 30116 27688 30168
rect 27740 30116 27828 30168
rect 27387 29950 27828 30116
rect 27387 29898 27476 29950
rect 27528 29898 27688 29950
rect 27740 29898 27828 29950
rect 27387 29733 27828 29898
rect 27387 29681 27476 29733
rect 27528 29681 27688 29733
rect 27740 29681 27828 29733
rect 27387 29515 27828 29681
rect 27387 29463 27476 29515
rect 27528 29463 27688 29515
rect 27740 29463 27828 29515
rect 27387 29297 27828 29463
rect 27387 29245 27476 29297
rect 27528 29245 27688 29297
rect 27740 29245 27828 29297
rect 27387 29080 27828 29245
rect 27387 29028 27476 29080
rect 27528 29028 27688 29080
rect 27740 29028 27828 29080
rect 27387 28862 27828 29028
rect 27387 28810 27476 28862
rect 27528 28810 27688 28862
rect 27740 28810 27828 28862
rect 27387 28644 27828 28810
rect 27387 28592 27476 28644
rect 27528 28592 27688 28644
rect 27740 28592 27828 28644
rect 27387 28427 27828 28592
rect 27387 28375 27476 28427
rect 27528 28375 27688 28427
rect 27740 28375 27828 28427
rect 27387 28209 27828 28375
rect 27387 28157 27476 28209
rect 27528 28157 27688 28209
rect 27740 28157 27828 28209
rect 27387 27992 27828 28157
rect 27387 27940 27476 27992
rect 27528 27940 27688 27992
rect 27740 27940 27828 27992
rect 27387 27774 27828 27940
rect 27387 27722 27476 27774
rect 27528 27722 27688 27774
rect 27740 27722 27828 27774
rect 27387 27556 27828 27722
rect 27387 27504 27476 27556
rect 27528 27504 27688 27556
rect 27740 27504 27828 27556
rect 25313 27267 25404 27323
rect 25460 27267 25528 27323
rect 25584 27267 25652 27323
rect 25708 27267 25776 27323
rect 25832 27267 25900 27323
rect 25956 27267 26039 27323
rect 25313 27199 26039 27267
rect 25313 27143 25404 27199
rect 25460 27143 25528 27199
rect 25584 27143 25652 27199
rect 25708 27143 25776 27199
rect 25832 27143 25900 27199
rect 25956 27143 26039 27199
rect 25313 27075 26039 27143
rect 25313 27019 25404 27075
rect 25460 27019 25528 27075
rect 25584 27019 25652 27075
rect 25708 27019 25776 27075
rect 25832 27019 25900 27075
rect 25956 27019 26039 27075
rect 25313 26951 26039 27019
rect 25313 26895 25404 26951
rect 25460 26895 25528 26951
rect 25584 26895 25652 26951
rect 25708 26895 25776 26951
rect 25832 26895 25900 26951
rect 25956 26895 26039 26951
rect 25313 26827 26039 26895
rect 25313 26771 25404 26827
rect 25460 26771 25528 26827
rect 25584 26771 25652 26827
rect 25708 26771 25776 26827
rect 25832 26771 25900 26827
rect 25956 26771 26039 26827
rect 25313 26703 26039 26771
rect 25313 26647 25404 26703
rect 25460 26647 25528 26703
rect 25584 26647 25652 26703
rect 25708 26647 25776 26703
rect 25832 26647 25900 26703
rect 25956 26647 26039 26703
rect 25313 26579 26039 26647
rect 25313 26523 25404 26579
rect 25460 26523 25528 26579
rect 25584 26523 25652 26579
rect 25708 26523 25776 26579
rect 25832 26523 25900 26579
rect 25956 26523 26039 26579
rect 25313 26433 26039 26523
rect 26823 27339 27163 27382
rect 26823 27287 26861 27339
rect 26913 27287 27073 27339
rect 27125 27287 27163 27339
rect 26823 27121 27163 27287
rect 26823 27069 26861 27121
rect 26913 27069 27073 27121
rect 27125 27069 27163 27121
rect 26823 26903 27163 27069
rect 26823 26851 26861 26903
rect 26913 26851 27073 26903
rect 27125 26851 27163 26903
rect 26823 26686 27163 26851
rect 26823 26634 26861 26686
rect 26913 26634 27073 26686
rect 27125 26634 27163 26686
rect 26823 26468 27163 26634
rect 26823 26416 26861 26468
rect 26913 26416 27073 26468
rect 27125 26416 27163 26468
rect 26435 26286 26643 26321
rect 26435 26126 26450 26286
rect 26610 26126 26643 26286
rect 26077 25967 26285 26002
rect 26077 25807 26092 25967
rect 26252 25807 26285 25967
rect 25741 25647 25949 25676
rect 25741 25487 25756 25647
rect 25916 25487 25949 25647
rect 25406 25328 25614 25357
rect 25406 25168 25421 25328
rect 25581 25168 25614 25328
rect 25066 24637 25274 24666
rect 25066 24477 25081 24637
rect 25241 24477 25274 24637
rect 24729 24316 24937 24345
rect 24729 24156 24744 24316
rect 24904 24156 24937 24316
rect 24401 23995 24609 24024
rect 24401 23835 24416 23995
rect 24576 23835 24609 23995
rect 24042 23673 24250 23702
rect 24042 23513 24057 23673
rect 24217 23513 24250 23673
rect 24042 17317 24250 23513
rect 24401 17656 24609 23835
rect 24729 17977 24937 24156
rect 25066 18350 25274 24477
rect 25406 18684 25614 25168
rect 25741 19027 25949 25487
rect 26077 19347 26285 25807
rect 26435 19692 26643 26126
rect 26435 19532 26465 19692
rect 26625 19532 26643 19692
rect 26435 19502 26643 19532
rect 26823 26250 27163 26416
rect 26823 26198 26861 26250
rect 26913 26198 27073 26250
rect 27125 26198 27163 26250
rect 26823 26033 27163 26198
rect 26823 25981 26861 26033
rect 26913 25981 27073 26033
rect 27125 25981 27163 26033
rect 26823 25815 27163 25981
rect 26823 25763 26861 25815
rect 26913 25763 27073 25815
rect 27125 25763 27163 25815
rect 26823 25598 27163 25763
rect 26823 25546 26861 25598
rect 26913 25546 27073 25598
rect 27125 25546 27163 25598
rect 26823 25380 27163 25546
rect 26823 25328 26861 25380
rect 26913 25328 27073 25380
rect 27125 25328 27163 25380
rect 26823 25162 27163 25328
rect 26823 25110 26861 25162
rect 26913 25110 27073 25162
rect 27125 25110 27163 25162
rect 26823 24945 27163 25110
rect 26823 24893 26861 24945
rect 26913 24893 27073 24945
rect 27125 24893 27163 24945
rect 26823 24727 27163 24893
rect 26823 24675 26861 24727
rect 26913 24675 27073 24727
rect 27125 24675 27163 24727
rect 26823 24509 27163 24675
rect 26823 24457 26861 24509
rect 26913 24457 27073 24509
rect 27125 24457 27163 24509
rect 26823 24292 27163 24457
rect 26823 24240 26861 24292
rect 26913 24240 27073 24292
rect 27125 24240 27163 24292
rect 26823 24075 27163 24240
rect 26823 23187 26858 24075
rect 27122 24074 27163 24075
rect 27125 24022 27163 24074
rect 27122 23857 27163 24022
rect 27125 23805 27163 23857
rect 27122 23639 27163 23805
rect 27125 23587 27163 23639
rect 27122 23421 27163 23587
rect 27125 23369 27163 23421
rect 27122 23204 27163 23369
rect 26823 23152 26861 23187
rect 26913 23152 27073 23187
rect 27125 23152 27163 23204
rect 26823 22986 27163 23152
rect 26823 22934 26861 22986
rect 26913 22934 27073 22986
rect 27125 22934 27163 22986
rect 26823 22768 27163 22934
rect 26823 22716 26861 22768
rect 26913 22716 27073 22768
rect 27125 22716 27163 22768
rect 26823 22551 27163 22716
rect 26823 22499 26861 22551
rect 26913 22499 27073 22551
rect 27125 22499 27163 22551
rect 26823 22333 27163 22499
rect 26823 22281 26861 22333
rect 26913 22281 27073 22333
rect 27125 22281 27163 22333
rect 26823 22115 27163 22281
rect 26823 22063 26861 22115
rect 26913 22063 27073 22115
rect 27125 22063 27163 22115
rect 26823 21898 27163 22063
rect 26823 21846 26861 21898
rect 26913 21846 27073 21898
rect 27125 21846 27163 21898
rect 26823 21680 27163 21846
rect 26823 21628 26861 21680
rect 26913 21628 27073 21680
rect 27125 21628 27163 21680
rect 26823 21463 27163 21628
rect 26823 21411 26861 21463
rect 26913 21411 27073 21463
rect 27125 21411 27163 21463
rect 26823 21245 27163 21411
rect 26823 21193 26861 21245
rect 26913 21193 27073 21245
rect 27125 21193 27163 21245
rect 26823 21027 27163 21193
rect 26823 20975 26861 21027
rect 26913 20975 27073 21027
rect 27125 20975 27163 21027
rect 26823 20810 27163 20975
rect 26823 20758 26861 20810
rect 26913 20758 27073 20810
rect 27125 20758 27163 20810
rect 26823 20592 27163 20758
rect 26823 20540 26861 20592
rect 26913 20570 27073 20592
rect 26913 20540 26924 20570
rect 27125 20540 27163 20592
rect 26823 20410 26924 20540
rect 27084 20410 27163 20540
rect 26823 20374 27163 20410
rect 26823 20322 26861 20374
rect 26913 20322 27073 20374
rect 27125 20322 27163 20374
rect 26823 20226 27163 20322
rect 26823 20157 26924 20226
rect 27084 20157 27163 20226
rect 26823 20105 26861 20157
rect 26913 20105 26924 20157
rect 27125 20105 27163 20157
rect 26823 20066 26924 20105
rect 27084 20066 27163 20105
rect 26823 19939 27163 20066
rect 26823 19887 26861 19939
rect 26913 19887 27073 19939
rect 27125 19887 27163 19939
rect 26823 19722 27163 19887
rect 26823 19670 26861 19722
rect 26913 19670 27073 19722
rect 27125 19670 27163 19722
rect 26823 19504 27163 19670
rect 26077 19187 26107 19347
rect 26267 19187 26285 19347
rect 26077 19162 26285 19187
rect 26823 19452 26861 19504
rect 26913 19452 27073 19504
rect 27125 19452 27163 19504
rect 26823 19286 27163 19452
rect 26823 19234 26861 19286
rect 26913 19234 27073 19286
rect 27125 19234 27163 19286
rect 25741 18867 25771 19027
rect 25931 18867 25949 19027
rect 25741 18822 25949 18867
rect 26823 19068 27163 19234
rect 26823 19016 26861 19068
rect 26913 19016 27073 19068
rect 27125 19016 27163 19068
rect 26823 18851 27163 19016
rect 25406 18524 25434 18684
rect 25594 18524 25614 18684
rect 25406 18482 25614 18524
rect 26823 18799 26861 18851
rect 26913 18799 27073 18851
rect 27125 18799 27163 18851
rect 26823 18633 27163 18799
rect 26823 18581 26861 18633
rect 26913 18581 27073 18633
rect 27125 18581 27163 18633
rect 25066 18190 25094 18350
rect 25254 18190 25274 18350
rect 25066 18142 25274 18190
rect 26823 18416 27163 18581
rect 26823 18364 26861 18416
rect 26913 18364 27073 18416
rect 27125 18364 27163 18416
rect 26823 18198 27163 18364
rect 26823 18146 26861 18198
rect 26913 18146 27073 18198
rect 27125 18146 27163 18198
rect 24729 17817 24757 17977
rect 24917 17817 24937 17977
rect 24729 17803 24937 17817
rect 26823 17980 27163 18146
rect 26823 17928 26861 17980
rect 26913 17928 27073 17980
rect 27125 17928 27163 17980
rect 24401 17496 24429 17656
rect 24589 17496 24609 17656
rect 24401 17462 24609 17496
rect 26823 17763 27163 17928
rect 26823 17711 26861 17763
rect 26913 17711 27073 17763
rect 27125 17711 27163 17763
rect 26823 17545 27163 17711
rect 26823 17493 26861 17545
rect 26913 17493 27073 17545
rect 27125 17493 27163 17545
rect 24042 17157 24069 17317
rect 24229 17157 24250 17317
rect 24042 17122 24250 17157
rect 26823 17327 27163 17493
rect 26823 17275 26861 17327
rect 26913 17275 27073 17327
rect 27125 17275 27163 17327
rect 26823 17110 27163 17275
rect 26823 17058 26861 17110
rect 26913 17058 27073 17110
rect 27125 17058 27163 17110
rect 26823 16892 27163 17058
rect 26823 16840 26861 16892
rect 26913 16840 27073 16892
rect 27125 16840 27163 16892
rect 26823 16675 27163 16840
rect 26823 16623 26861 16675
rect 26913 16623 27073 16675
rect 27125 16623 27163 16675
rect 26823 16457 27163 16623
rect 26823 16405 26861 16457
rect 26913 16405 27073 16457
rect 27125 16405 27163 16457
rect 26823 16239 27163 16405
rect 26823 16187 26861 16239
rect 26913 16187 27073 16239
rect 27125 16187 27163 16239
rect 26823 16022 27163 16187
rect 26823 15970 26861 16022
rect 26913 15970 27073 16022
rect 27125 15970 27163 16022
rect 26823 15804 27163 15970
rect 26823 15752 26861 15804
rect 26913 15752 27073 15804
rect 27125 15752 27163 15804
rect 26823 15586 27163 15752
rect 26823 15534 26861 15586
rect 26913 15534 27073 15586
rect 27125 15534 27163 15586
rect 26823 15369 27163 15534
rect 26823 15317 26861 15369
rect 26913 15317 27073 15369
rect 27125 15317 27163 15369
rect 26823 15151 27163 15317
rect 26823 15099 26861 15151
rect 26913 15099 27073 15151
rect 27125 15099 27163 15151
rect 26823 14933 27163 15099
rect 26823 14881 26861 14933
rect 26913 14881 27073 14933
rect 27125 14881 27163 14933
rect 26823 14716 27163 14881
rect 26823 14664 26861 14716
rect 26913 14664 27073 14716
rect 27125 14664 27163 14716
rect 26823 14498 27163 14664
rect 26823 14446 26861 14498
rect 26913 14446 27073 14498
rect 27125 14446 27163 14498
rect 26823 14281 27163 14446
rect 26823 14229 26861 14281
rect 26913 14229 27073 14281
rect 27125 14229 27163 14281
rect 26823 14119 27163 14229
rect 26823 14063 26859 14119
rect 26915 14063 27071 14119
rect 27127 14063 27163 14119
rect 26823 14011 26861 14063
rect 26913 14011 27073 14063
rect 27125 14011 27163 14063
rect 26823 13902 27163 14011
rect 26823 13846 26859 13902
rect 26915 13846 27071 13902
rect 27127 13846 27163 13902
rect 26823 13845 27163 13846
rect 26823 13793 26861 13845
rect 26913 13793 27073 13845
rect 27125 13793 27163 13845
rect 26823 13684 27163 13793
rect 26823 13628 26859 13684
rect 26915 13628 27071 13684
rect 27127 13628 27163 13684
rect 26823 13576 26861 13628
rect 26913 13576 27073 13628
rect 27125 13576 27163 13628
rect 26823 13467 27163 13576
rect 26823 13411 26859 13467
rect 26915 13411 27071 13467
rect 27127 13411 27163 13467
rect 26823 13410 27163 13411
rect 26823 13358 26861 13410
rect 26913 13358 27073 13410
rect 27125 13358 27163 13410
rect 26823 13249 27163 13358
rect 26823 13193 26859 13249
rect 26915 13193 27071 13249
rect 27127 13193 27163 13249
rect 26823 13192 27163 13193
rect 26823 13140 26861 13192
rect 26913 13140 27073 13192
rect 27125 13140 27163 13192
rect 26823 13031 27163 13140
rect 26823 12975 26859 13031
rect 26915 12975 27071 13031
rect 27127 12975 27163 13031
rect 26823 12923 26861 12975
rect 26913 12923 27073 12975
rect 27125 12923 27163 12975
rect 26823 12813 27163 12923
rect 26823 12757 26859 12813
rect 26915 12757 27071 12813
rect 27127 12757 27163 12813
rect 26823 12705 26861 12757
rect 26913 12705 27073 12757
rect 27125 12705 27163 12757
rect 26823 12596 27163 12705
rect 26823 12540 26859 12596
rect 26915 12540 27071 12596
rect 27127 12540 27163 12596
rect 26823 12488 26861 12540
rect 26913 12488 27073 12540
rect 27125 12488 27163 12540
rect 26823 12378 27163 12488
rect 26823 12322 26859 12378
rect 26915 12322 27071 12378
rect 27127 12322 27163 12378
rect 26823 12270 26861 12322
rect 26913 12270 27073 12322
rect 27125 12270 27163 12322
rect 26823 12161 27163 12270
rect 26823 12105 26859 12161
rect 26915 12105 27071 12161
rect 27127 12105 27163 12161
rect 26823 12104 27163 12105
rect 26823 12052 26861 12104
rect 26913 12052 27073 12104
rect 27125 12052 27163 12104
rect 26823 11887 27163 12052
rect 26823 11835 26861 11887
rect 26913 11835 27073 11887
rect 27125 11835 27163 11887
rect 26823 11669 27163 11835
rect 26823 11617 26861 11669
rect 26913 11617 27073 11669
rect 27125 11617 27163 11669
rect 26823 11451 27163 11617
rect 26823 11399 26861 11451
rect 26913 11399 27073 11451
rect 27125 11399 27163 11451
rect 26823 11234 27163 11399
rect 26823 11182 26861 11234
rect 26913 11182 27073 11234
rect 27125 11182 27163 11234
rect 26823 11016 27163 11182
rect 26823 10964 26861 11016
rect 26913 10964 27073 11016
rect 27125 10964 27163 11016
rect 26823 10798 27163 10964
rect 26823 10746 26861 10798
rect 26913 10746 27073 10798
rect 27125 10746 27163 10798
rect 26823 10581 27163 10746
rect 26823 10529 26861 10581
rect 26913 10529 27073 10581
rect 27125 10529 27163 10581
rect 26823 10363 27163 10529
rect 26823 10311 26861 10363
rect 26913 10311 27073 10363
rect 27125 10311 27163 10363
rect 26823 10146 27163 10311
rect 26823 10094 26861 10146
rect 26913 10094 27073 10146
rect 27125 10094 27163 10146
rect 26823 9928 27163 10094
rect 26823 9876 26861 9928
rect 26913 9876 27073 9928
rect 27125 9876 27163 9928
rect 26823 9710 27163 9876
rect 26823 9658 26861 9710
rect 26913 9658 27073 9710
rect 27125 9658 27163 9710
rect 26823 9493 27163 9658
rect 26823 9441 26861 9493
rect 26913 9441 27073 9493
rect 27125 9441 27163 9493
rect 26823 9407 27163 9441
rect 26823 9351 26859 9407
rect 26915 9351 27071 9407
rect 27127 9351 27163 9407
rect 26823 9275 27163 9351
rect 26823 9223 26861 9275
rect 26913 9223 27073 9275
rect 27125 9223 27163 9275
rect 26823 9190 27163 9223
rect 26823 9134 26859 9190
rect 26915 9134 27071 9190
rect 27127 9134 27163 9190
rect 26823 9057 27163 9134
rect 26823 9005 26861 9057
rect 26913 9005 27073 9057
rect 27125 9005 27163 9057
rect 26823 8972 27163 9005
rect 26823 8916 26859 8972
rect 26915 8916 27071 8972
rect 27127 8916 27163 8972
rect 26823 8840 27163 8916
rect 26823 8788 26861 8840
rect 26913 8788 27073 8840
rect 27125 8788 27163 8840
rect 26823 8754 27163 8788
rect 26823 8698 26859 8754
rect 26915 8698 27071 8754
rect 27127 8698 27163 8754
rect 26823 8622 27163 8698
rect 26823 8570 26861 8622
rect 26913 8570 27073 8622
rect 27125 8570 27163 8622
rect 26823 8536 27163 8570
rect 26823 8480 26859 8536
rect 26915 8480 27071 8536
rect 27127 8480 27163 8536
rect 26823 8404 27163 8480
rect 26823 8352 26861 8404
rect 26913 8352 27073 8404
rect 27125 8352 27163 8404
rect 26823 8319 27163 8352
rect 26823 8263 26859 8319
rect 26915 8263 27071 8319
rect 27127 8263 27163 8319
rect 26823 8187 27163 8263
rect 26823 8135 26861 8187
rect 26913 8135 27073 8187
rect 27125 8135 27163 8187
rect 26823 7969 27163 8135
rect 26823 7917 26861 7969
rect 26913 7917 27073 7969
rect 27125 7917 27163 7969
rect 26823 7752 27163 7917
rect 26823 7700 26861 7752
rect 26913 7700 27073 7752
rect 27125 7700 27163 7752
rect 26823 7534 27163 7700
rect 26823 7482 26861 7534
rect 26913 7482 27073 7534
rect 27125 7482 27163 7534
rect 26823 7316 27163 7482
rect 26823 7264 26861 7316
rect 26913 7264 27073 7316
rect 27125 7264 27163 7316
rect 26823 7099 27163 7264
rect 26823 7047 26861 7099
rect 26913 7047 27073 7099
rect 27125 7047 27163 7099
rect 26823 6881 27163 7047
rect 26823 6829 26861 6881
rect 26913 6829 27073 6881
rect 27125 6829 27163 6881
rect 26823 6663 27163 6829
rect 26823 6611 26861 6663
rect 26913 6611 27073 6663
rect 27125 6611 27163 6663
rect 26823 6446 27163 6611
rect 26823 6394 26861 6446
rect 26913 6394 27073 6446
rect 27125 6394 27163 6446
rect 26823 6228 27163 6394
rect 26823 6176 26861 6228
rect 26913 6176 27073 6228
rect 27125 6176 27163 6228
rect 26823 6011 27163 6176
rect 26823 5959 26861 6011
rect 26913 5959 27073 6011
rect 27125 5959 27163 6011
rect 26823 5793 27163 5959
rect 26823 5741 26861 5793
rect 26913 5741 27073 5793
rect 27125 5741 27163 5793
rect 26823 5575 27163 5741
rect 26823 5539 26861 5575
rect 26913 5539 27073 5575
rect 27125 5539 27163 5575
rect 26823 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27163 5539
rect 26823 5358 27163 5483
rect 26823 5321 26861 5358
rect 26913 5321 27073 5358
rect 27125 5321 27163 5358
rect 26823 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27163 5321
rect 26823 5226 27163 5265
rect 27387 27339 27828 27504
rect 27387 27287 27476 27339
rect 27528 27287 27688 27339
rect 27740 27287 27828 27339
rect 27387 27121 27828 27287
rect 27387 27069 27476 27121
rect 27528 27069 27688 27121
rect 27740 27069 27828 27121
rect 27387 26903 27828 27069
rect 27387 26851 27476 26903
rect 27528 26851 27688 26903
rect 27740 26851 27828 26903
rect 27387 26799 27828 26851
rect 27387 26743 27474 26799
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 27387 26686 27828 26743
rect 27387 26634 27476 26686
rect 27528 26634 27688 26686
rect 27740 26634 27828 26686
rect 27387 26581 27828 26634
rect 27387 26525 27474 26581
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 27387 26468 27828 26525
rect 27387 26416 27476 26468
rect 27528 26416 27688 26468
rect 27740 26416 27828 26468
rect 27387 26250 27828 26416
rect 27387 26198 27476 26250
rect 27528 26198 27688 26250
rect 27740 26198 27828 26250
rect 27387 26033 27828 26198
rect 27387 25981 27476 26033
rect 27528 25981 27688 26033
rect 27740 25981 27828 26033
rect 27387 25815 27828 25981
rect 27387 25763 27476 25815
rect 27528 25763 27688 25815
rect 27740 25763 27828 25815
rect 27387 25598 27828 25763
rect 27387 25546 27476 25598
rect 27528 25546 27688 25598
rect 27740 25546 27828 25598
rect 27387 25380 27828 25546
rect 27387 25328 27476 25380
rect 27528 25328 27688 25380
rect 27740 25328 27828 25380
rect 27387 25162 27828 25328
rect 27387 25110 27476 25162
rect 27528 25110 27688 25162
rect 27740 25110 27828 25162
rect 27387 25028 27828 25110
rect 27387 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 27828 25028
rect 27387 24945 27828 24972
rect 27387 24893 27476 24945
rect 27528 24893 27688 24945
rect 27740 24893 27828 24945
rect 27387 24810 27828 24893
rect 27387 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 27828 24810
rect 27387 24727 27828 24754
rect 27387 24675 27476 24727
rect 27528 24675 27688 24727
rect 27740 24675 27828 24727
rect 27387 24509 27828 24675
rect 27387 24457 27476 24509
rect 27528 24457 27688 24509
rect 27740 24457 27828 24509
rect 27387 24292 27828 24457
rect 27387 24240 27476 24292
rect 27528 24240 27688 24292
rect 27740 24240 27828 24292
rect 27387 24074 27828 24240
rect 27387 24022 27476 24074
rect 27528 24022 27688 24074
rect 27740 24022 27828 24074
rect 27387 23857 27828 24022
rect 27387 23805 27476 23857
rect 27528 23805 27688 23857
rect 27740 23805 27828 23857
rect 27387 23639 27828 23805
rect 27387 23587 27476 23639
rect 27528 23587 27688 23639
rect 27740 23587 27828 23639
rect 27387 23421 27828 23587
rect 27387 23369 27476 23421
rect 27528 23369 27688 23421
rect 27740 23369 27828 23421
rect 27387 23204 27828 23369
rect 27387 23152 27476 23204
rect 27528 23152 27688 23204
rect 27740 23152 27828 23204
rect 27387 22986 27828 23152
rect 27387 22936 27476 22986
rect 27528 22936 27688 22986
rect 27387 22048 27475 22936
rect 27740 22934 27828 22986
rect 27739 22768 27828 22934
rect 27740 22716 27828 22768
rect 27739 22551 27828 22716
rect 27740 22499 27828 22551
rect 27739 22333 27828 22499
rect 27740 22281 27828 22333
rect 27739 22115 27828 22281
rect 27740 22063 27828 22115
rect 27739 22048 27828 22063
rect 27387 21898 27828 22048
rect 27387 21846 27476 21898
rect 27528 21846 27688 21898
rect 27740 21846 27828 21898
rect 27387 21680 27828 21846
rect 27387 21628 27476 21680
rect 27528 21628 27688 21680
rect 27740 21628 27828 21680
rect 27387 21463 27828 21628
rect 27387 21411 27476 21463
rect 27528 21411 27688 21463
rect 27740 21411 27828 21463
rect 27387 21245 27828 21411
rect 27387 21193 27476 21245
rect 27528 21193 27688 21245
rect 27740 21193 27828 21245
rect 27387 21027 27828 21193
rect 27387 20975 27476 21027
rect 27528 20975 27688 21027
rect 27740 20975 27828 21027
rect 27387 20810 27828 20975
rect 27387 20758 27476 20810
rect 27528 20758 27688 20810
rect 27740 20758 27828 20810
rect 27387 20592 27828 20758
rect 27387 20540 27476 20592
rect 27528 20540 27688 20592
rect 27740 20540 27828 20592
rect 27387 20374 27828 20540
rect 27387 20322 27476 20374
rect 27528 20322 27688 20374
rect 27740 20322 27828 20374
rect 27387 20157 27828 20322
rect 27387 20105 27476 20157
rect 27528 20105 27688 20157
rect 27740 20105 27828 20157
rect 27387 19939 27828 20105
rect 27387 19887 27476 19939
rect 27528 19887 27688 19939
rect 27740 19887 27828 19939
rect 27387 19722 27828 19887
rect 27387 19670 27476 19722
rect 27528 19670 27688 19722
rect 27740 19670 27828 19722
rect 27387 19504 27828 19670
rect 27387 19452 27476 19504
rect 27528 19452 27688 19504
rect 27740 19452 27828 19504
rect 27387 19286 27828 19452
rect 27387 19234 27476 19286
rect 27528 19234 27688 19286
rect 27740 19234 27828 19286
rect 27387 19068 27828 19234
rect 27387 19016 27476 19068
rect 27528 19016 27688 19068
rect 27740 19016 27828 19068
rect 27387 18851 27828 19016
rect 27387 18799 27476 18851
rect 27528 18799 27688 18851
rect 27740 18799 27828 18851
rect 27387 18633 27828 18799
rect 27387 18581 27476 18633
rect 27528 18581 27688 18633
rect 27740 18581 27828 18633
rect 27387 18416 27828 18581
rect 27387 18364 27476 18416
rect 27528 18364 27688 18416
rect 27740 18364 27828 18416
rect 27387 18198 27828 18364
rect 27387 18146 27476 18198
rect 27528 18146 27688 18198
rect 27740 18146 27828 18198
rect 27387 17980 27828 18146
rect 27387 17928 27476 17980
rect 27528 17928 27688 17980
rect 27740 17928 27828 17980
rect 27387 17763 27828 17928
rect 27387 17711 27476 17763
rect 27528 17711 27688 17763
rect 27740 17711 27828 17763
rect 27387 17545 27828 17711
rect 27387 17493 27476 17545
rect 27528 17493 27688 17545
rect 27740 17493 27828 17545
rect 27387 17327 27828 17493
rect 27387 17275 27476 17327
rect 27528 17275 27688 17327
rect 27740 17275 27828 17327
rect 27387 17110 27828 17275
rect 27387 17058 27476 17110
rect 27528 17058 27688 17110
rect 27740 17058 27828 17110
rect 27387 16892 27828 17058
rect 27387 16840 27476 16892
rect 27528 16840 27688 16892
rect 27740 16840 27828 16892
rect 27387 16675 27828 16840
rect 27387 16623 27476 16675
rect 27528 16623 27688 16675
rect 27740 16623 27828 16675
rect 27387 16470 27828 16623
rect 27387 16414 27474 16470
rect 27530 16414 27686 16470
rect 27742 16414 27828 16470
rect 27387 16405 27476 16414
rect 27528 16405 27688 16414
rect 27740 16405 27828 16414
rect 27387 16253 27828 16405
rect 27387 16197 27474 16253
rect 27530 16197 27686 16253
rect 27742 16197 27828 16253
rect 27387 16187 27476 16197
rect 27528 16187 27688 16197
rect 27740 16187 27828 16197
rect 27387 16035 27828 16187
rect 27387 15979 27474 16035
rect 27530 15979 27686 16035
rect 27742 15979 27828 16035
rect 27387 15970 27476 15979
rect 27528 15970 27688 15979
rect 27740 15970 27828 15979
rect 27387 15818 27828 15970
rect 27387 15762 27474 15818
rect 27530 15762 27686 15818
rect 27742 15762 27828 15818
rect 27387 15752 27476 15762
rect 27528 15752 27688 15762
rect 27740 15752 27828 15762
rect 27387 15600 27828 15752
rect 27387 15544 27474 15600
rect 27530 15544 27686 15600
rect 27742 15544 27828 15600
rect 27387 15534 27476 15544
rect 27528 15534 27688 15544
rect 27740 15534 27828 15544
rect 27387 15382 27828 15534
rect 27387 15326 27474 15382
rect 27530 15326 27686 15382
rect 27742 15326 27828 15382
rect 27387 15317 27476 15326
rect 27528 15317 27688 15326
rect 27740 15317 27828 15326
rect 27387 15164 27828 15317
rect 27387 15108 27474 15164
rect 27530 15108 27686 15164
rect 27742 15108 27828 15164
rect 27387 15099 27476 15108
rect 27528 15099 27688 15108
rect 27740 15099 27828 15108
rect 27387 14947 27828 15099
rect 27387 14891 27474 14947
rect 27530 14891 27686 14947
rect 27742 14891 27828 14947
rect 27387 14881 27476 14891
rect 27528 14881 27688 14891
rect 27740 14881 27828 14891
rect 27387 14729 27828 14881
rect 27387 14673 27474 14729
rect 27530 14673 27686 14729
rect 27742 14673 27828 14729
rect 27387 14664 27476 14673
rect 27528 14664 27688 14673
rect 27740 14664 27828 14673
rect 27387 14512 27828 14664
rect 27387 14456 27474 14512
rect 27530 14456 27686 14512
rect 27742 14456 27828 14512
rect 27387 14446 27476 14456
rect 27528 14446 27688 14456
rect 27740 14446 27828 14456
rect 27387 14281 27828 14446
rect 27387 14231 27476 14281
rect 27528 14231 27688 14281
rect 27740 14231 27828 14281
rect 27387 14175 27474 14231
rect 27530 14175 27686 14231
rect 27742 14175 27828 14231
rect 27387 14063 27828 14175
rect 27387 14014 27476 14063
rect 27528 14014 27688 14063
rect 27740 14014 27828 14063
rect 27387 13958 27474 14014
rect 27530 13958 27686 14014
rect 27742 13958 27828 14014
rect 27387 13845 27828 13958
rect 27387 13796 27476 13845
rect 27528 13796 27688 13845
rect 27740 13796 27828 13845
rect 27387 13740 27474 13796
rect 27530 13740 27686 13796
rect 27742 13740 27828 13796
rect 27387 13628 27828 13740
rect 27387 13578 27476 13628
rect 27528 13578 27688 13628
rect 27740 13578 27828 13628
rect 27387 13522 27474 13578
rect 27530 13522 27686 13578
rect 27742 13522 27828 13578
rect 27387 13410 27828 13522
rect 27387 13361 27476 13410
rect 27528 13361 27688 13410
rect 27740 13361 27828 13410
rect 27387 13305 27474 13361
rect 27530 13305 27686 13361
rect 27742 13305 27828 13361
rect 27387 13192 27828 13305
rect 27387 13140 27476 13192
rect 27528 13140 27688 13192
rect 27740 13140 27828 13192
rect 27387 12975 27828 13140
rect 27387 12923 27476 12975
rect 27528 12923 27688 12975
rect 27740 12923 27828 12975
rect 27387 12757 27828 12923
rect 27387 12705 27476 12757
rect 27528 12705 27688 12757
rect 27740 12705 27828 12757
rect 27387 12540 27828 12705
rect 27387 12488 27476 12540
rect 27528 12488 27688 12540
rect 27740 12488 27828 12540
rect 27387 12322 27828 12488
rect 27387 12270 27476 12322
rect 27528 12270 27688 12322
rect 27740 12270 27828 12322
rect 27387 12104 27828 12270
rect 27387 12052 27476 12104
rect 27528 12052 27688 12104
rect 27740 12052 27828 12104
rect 27387 11887 27828 12052
rect 27387 11835 27476 11887
rect 27528 11835 27688 11887
rect 27740 11835 27828 11887
rect 27387 11669 27828 11835
rect 27387 11617 27476 11669
rect 27528 11617 27688 11669
rect 27740 11617 27828 11669
rect 27387 11451 27828 11617
rect 27387 11406 27476 11451
rect 27528 11406 27688 11451
rect 27740 11406 27828 11451
rect 27387 11350 27474 11406
rect 27530 11350 27686 11406
rect 27742 11350 27828 11406
rect 27387 11234 27828 11350
rect 27387 11189 27476 11234
rect 27528 11189 27688 11234
rect 27740 11189 27828 11234
rect 27387 11133 27474 11189
rect 27530 11133 27686 11189
rect 27742 11133 27828 11189
rect 27387 11016 27828 11133
rect 27387 10971 27476 11016
rect 27528 10971 27688 11016
rect 27740 10971 27828 11016
rect 27387 10915 27474 10971
rect 27530 10915 27686 10971
rect 27742 10915 27828 10971
rect 27387 10798 27828 10915
rect 27387 10753 27476 10798
rect 27528 10753 27688 10798
rect 27740 10753 27828 10798
rect 27387 10697 27474 10753
rect 27530 10697 27686 10753
rect 27742 10697 27828 10753
rect 27387 10581 27828 10697
rect 27387 10535 27476 10581
rect 27528 10535 27688 10581
rect 27740 10535 27828 10581
rect 27387 10479 27474 10535
rect 27530 10479 27686 10535
rect 27742 10479 27828 10535
rect 27387 10363 27828 10479
rect 27387 10318 27476 10363
rect 27528 10318 27688 10363
rect 27740 10318 27828 10363
rect 27387 10262 27474 10318
rect 27530 10262 27686 10318
rect 27742 10262 27828 10318
rect 27387 10146 27828 10262
rect 27387 10094 27476 10146
rect 27528 10094 27688 10146
rect 27740 10094 27828 10146
rect 27387 9928 27828 10094
rect 57295 33215 57736 33380
rect 57295 33163 57383 33215
rect 57435 33163 57595 33215
rect 57647 33163 57736 33215
rect 57295 33141 57736 33163
rect 57295 33085 57381 33141
rect 57437 33085 57593 33141
rect 57649 33085 57736 33141
rect 57295 32997 57736 33085
rect 57295 32945 57383 32997
rect 57435 32945 57595 32997
rect 57647 32945 57736 32997
rect 57295 32923 57736 32945
rect 57295 32867 57381 32923
rect 57437 32867 57593 32923
rect 57649 32867 57736 32923
rect 57295 32779 57736 32867
rect 57295 32727 57383 32779
rect 57435 32727 57595 32779
rect 57647 32727 57736 32779
rect 57295 32705 57736 32727
rect 57295 32649 57381 32705
rect 57437 32649 57593 32705
rect 57649 32649 57736 32705
rect 57295 32562 57736 32649
rect 57295 32510 57383 32562
rect 57435 32510 57595 32562
rect 57647 32510 57736 32562
rect 57295 32487 57736 32510
rect 57295 32431 57381 32487
rect 57437 32431 57593 32487
rect 57649 32431 57736 32487
rect 57295 32344 57736 32431
rect 57295 32292 57383 32344
rect 57435 32292 57595 32344
rect 57647 32292 57736 32344
rect 57295 32127 57736 32292
rect 57295 32075 57383 32127
rect 57435 32075 57595 32127
rect 57647 32075 57736 32127
rect 57295 31909 57736 32075
rect 57295 31857 57383 31909
rect 57435 31857 57595 31909
rect 57647 31857 57736 31909
rect 57295 31691 57736 31857
rect 57295 31639 57383 31691
rect 57435 31639 57595 31691
rect 57647 31639 57736 31691
rect 57295 31474 57736 31639
rect 57295 31422 57383 31474
rect 57435 31422 57595 31474
rect 57647 31422 57736 31474
rect 57295 31256 57736 31422
rect 57295 31252 57383 31256
rect 57435 31252 57595 31256
rect 57647 31252 57736 31256
rect 57295 31196 57381 31252
rect 57437 31196 57593 31252
rect 57649 31196 57736 31252
rect 57295 31038 57736 31196
rect 57295 31034 57383 31038
rect 57435 31034 57595 31038
rect 57647 31034 57736 31038
rect 57295 30978 57381 31034
rect 57437 30978 57593 31034
rect 57649 30978 57736 31034
rect 57295 30821 57736 30978
rect 57295 30816 57383 30821
rect 57435 30816 57595 30821
rect 57647 30816 57736 30821
rect 57295 30760 57381 30816
rect 57437 30760 57593 30816
rect 57649 30760 57736 30816
rect 57295 30603 57736 30760
rect 57295 30598 57383 30603
rect 57435 30598 57595 30603
rect 57647 30598 57736 30603
rect 57295 30542 57381 30598
rect 57437 30542 57593 30598
rect 57649 30542 57736 30598
rect 57295 30386 57736 30542
rect 57295 30334 57383 30386
rect 57435 30334 57595 30386
rect 57647 30334 57736 30386
rect 57295 30168 57736 30334
rect 57295 30116 57383 30168
rect 57435 30116 57595 30168
rect 57647 30116 57736 30168
rect 57295 29950 57736 30116
rect 57295 29898 57383 29950
rect 57435 29898 57595 29950
rect 57647 29898 57736 29950
rect 57295 29733 57736 29898
rect 57295 29681 57383 29733
rect 57435 29681 57595 29733
rect 57647 29681 57736 29733
rect 57295 29515 57736 29681
rect 57295 29463 57383 29515
rect 57435 29463 57595 29515
rect 57647 29463 57736 29515
rect 57295 29297 57736 29463
rect 57295 29245 57383 29297
rect 57435 29245 57595 29297
rect 57647 29245 57736 29297
rect 57295 29080 57736 29245
rect 57295 29028 57383 29080
rect 57435 29028 57595 29080
rect 57647 29028 57736 29080
rect 57295 28862 57736 29028
rect 57295 28810 57383 28862
rect 57435 28810 57595 28862
rect 57647 28810 57736 28862
rect 57295 28644 57736 28810
rect 57295 28592 57383 28644
rect 57435 28592 57595 28644
rect 57647 28592 57736 28644
rect 57295 28427 57736 28592
rect 57295 28375 57383 28427
rect 57435 28375 57595 28427
rect 57647 28375 57736 28427
rect 57295 28209 57736 28375
rect 57295 28157 57383 28209
rect 57435 28157 57595 28209
rect 57647 28157 57736 28209
rect 57295 27992 57736 28157
rect 57295 27940 57383 27992
rect 57435 27940 57595 27992
rect 57647 27940 57736 27992
rect 57295 27774 57736 27940
rect 57295 27722 57383 27774
rect 57435 27722 57595 27774
rect 57647 27722 57736 27774
rect 57295 27556 57736 27722
rect 57295 27504 57383 27556
rect 57435 27504 57595 27556
rect 57647 27504 57736 27556
rect 57295 27339 57736 27504
rect 57295 27287 57383 27339
rect 57435 27287 57595 27339
rect 57647 27287 57736 27339
rect 57295 27121 57736 27287
rect 57295 27069 57383 27121
rect 57435 27069 57595 27121
rect 57647 27069 57736 27121
rect 57295 26903 57736 27069
rect 57295 26851 57383 26903
rect 57435 26851 57595 26903
rect 57647 26851 57736 26903
rect 57295 26799 57736 26851
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26743 57736 26799
rect 57295 26686 57736 26743
rect 57295 26634 57383 26686
rect 57435 26634 57595 26686
rect 57647 26634 57736 26686
rect 57295 26581 57736 26634
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26525 57736 26581
rect 57295 26468 57736 26525
rect 57295 26416 57383 26468
rect 57435 26416 57595 26468
rect 57647 26416 57736 26468
rect 57295 26250 57736 26416
rect 57295 26198 57383 26250
rect 57435 26198 57595 26250
rect 57647 26198 57736 26250
rect 57295 26033 57736 26198
rect 57295 25981 57383 26033
rect 57435 25981 57595 26033
rect 57647 25981 57736 26033
rect 57295 25815 57736 25981
rect 57295 25763 57383 25815
rect 57435 25763 57595 25815
rect 57647 25763 57736 25815
rect 57295 25598 57736 25763
rect 57295 25546 57383 25598
rect 57435 25546 57595 25598
rect 57647 25546 57736 25598
rect 57295 25380 57736 25546
rect 57295 25328 57383 25380
rect 57435 25328 57595 25380
rect 57647 25328 57736 25380
rect 57295 25162 57736 25328
rect 57295 25110 57383 25162
rect 57435 25110 57595 25162
rect 57647 25110 57736 25162
rect 57295 24945 57736 25110
rect 57295 24893 57383 24945
rect 57435 24893 57595 24945
rect 57647 24893 57736 24945
rect 57295 24727 57736 24893
rect 57295 24675 57383 24727
rect 57435 24675 57595 24727
rect 57647 24675 57736 24727
rect 57295 24509 57736 24675
rect 57295 24457 57383 24509
rect 57435 24457 57595 24509
rect 57647 24457 57736 24509
rect 57295 24292 57736 24457
rect 57295 24240 57383 24292
rect 57435 24240 57595 24292
rect 57647 24240 57736 24292
rect 57295 24074 57736 24240
rect 57295 24022 57383 24074
rect 57435 24022 57595 24074
rect 57647 24022 57736 24074
rect 57295 23857 57736 24022
rect 57295 23805 57383 23857
rect 57435 23805 57595 23857
rect 57647 23805 57736 23857
rect 57295 23639 57736 23805
rect 57295 23587 57383 23639
rect 57435 23587 57595 23639
rect 57647 23587 57736 23639
rect 57295 23421 57736 23587
rect 57295 23369 57383 23421
rect 57435 23369 57595 23421
rect 57647 23369 57736 23421
rect 57295 23204 57736 23369
rect 57295 23152 57383 23204
rect 57435 23152 57595 23204
rect 57647 23152 57736 23204
rect 57295 22986 57736 23152
rect 57295 22934 57383 22986
rect 57435 22934 57595 22986
rect 57647 22934 57736 22986
rect 57295 22923 57736 22934
rect 57295 22035 57363 22923
rect 57627 22768 57736 22923
rect 57647 22716 57736 22768
rect 57627 22551 57736 22716
rect 57647 22499 57736 22551
rect 57627 22333 57736 22499
rect 57647 22281 57736 22333
rect 57627 22115 57736 22281
rect 57647 22063 57736 22115
rect 57627 22035 57736 22063
rect 57295 21898 57736 22035
rect 57295 21846 57383 21898
rect 57435 21846 57595 21898
rect 57647 21846 57736 21898
rect 57295 21680 57736 21846
rect 57295 21628 57383 21680
rect 57435 21628 57595 21680
rect 57647 21628 57736 21680
rect 57295 21463 57736 21628
rect 57295 21411 57383 21463
rect 57435 21411 57595 21463
rect 57647 21411 57736 21463
rect 57295 21245 57736 21411
rect 57295 21193 57383 21245
rect 57435 21193 57595 21245
rect 57647 21193 57736 21245
rect 57295 21027 57736 21193
rect 57295 20975 57383 21027
rect 57435 20975 57595 21027
rect 57647 20975 57736 21027
rect 57295 20810 57736 20975
rect 57295 20758 57383 20810
rect 57435 20758 57595 20810
rect 57647 20758 57736 20810
rect 57295 20592 57736 20758
rect 57295 20540 57383 20592
rect 57435 20540 57595 20592
rect 57647 20540 57736 20592
rect 57295 20374 57736 20540
rect 57295 20322 57383 20374
rect 57435 20322 57595 20374
rect 57647 20322 57736 20374
rect 57295 20157 57736 20322
rect 57295 20105 57383 20157
rect 57435 20105 57595 20157
rect 57647 20105 57736 20157
rect 57295 19939 57736 20105
rect 57295 19887 57383 19939
rect 57435 19887 57595 19939
rect 57647 19887 57736 19939
rect 57295 19722 57736 19887
rect 57295 19670 57383 19722
rect 57435 19670 57595 19722
rect 57647 19670 57736 19722
rect 57295 19504 57736 19670
rect 57295 19452 57383 19504
rect 57435 19452 57595 19504
rect 57647 19452 57736 19504
rect 57295 19286 57736 19452
rect 57295 19234 57383 19286
rect 57435 19234 57595 19286
rect 57647 19234 57736 19286
rect 57295 19068 57736 19234
rect 57295 19016 57383 19068
rect 57435 19016 57595 19068
rect 57647 19016 57736 19068
rect 57295 18851 57736 19016
rect 57295 18799 57383 18851
rect 57435 18799 57595 18851
rect 57647 18799 57736 18851
rect 57295 18633 57736 18799
rect 57295 18581 57383 18633
rect 57435 18581 57595 18633
rect 57647 18581 57736 18633
rect 57295 18416 57736 18581
rect 57295 18364 57383 18416
rect 57435 18364 57595 18416
rect 57647 18364 57736 18416
rect 57295 18198 57736 18364
rect 57295 18146 57383 18198
rect 57435 18146 57595 18198
rect 57647 18146 57736 18198
rect 57295 17980 57736 18146
rect 57295 17928 57383 17980
rect 57435 17928 57595 17980
rect 57647 17928 57736 17980
rect 57295 17763 57736 17928
rect 57295 17711 57383 17763
rect 57435 17711 57595 17763
rect 57647 17711 57736 17763
rect 57295 17545 57736 17711
rect 57295 17493 57383 17545
rect 57435 17493 57595 17545
rect 57647 17493 57736 17545
rect 57295 17327 57736 17493
rect 57295 17275 57383 17327
rect 57435 17275 57595 17327
rect 57647 17275 57736 17327
rect 57295 17110 57736 17275
rect 57295 17058 57383 17110
rect 57435 17058 57595 17110
rect 57647 17058 57736 17110
rect 57295 16892 57736 17058
rect 57295 16840 57383 16892
rect 57435 16840 57595 16892
rect 57647 16840 57736 16892
rect 57295 16678 57736 16840
rect 57295 16622 57381 16678
rect 57437 16622 57593 16678
rect 57649 16622 57736 16678
rect 57295 16461 57736 16622
rect 57295 16405 57381 16461
rect 57437 16405 57593 16461
rect 57649 16405 57736 16461
rect 57295 16243 57736 16405
rect 57295 16187 57381 16243
rect 57437 16187 57593 16243
rect 57649 16187 57736 16243
rect 57295 16026 57736 16187
rect 57295 15970 57381 16026
rect 57437 15970 57593 16026
rect 57649 15970 57736 16026
rect 57295 15808 57736 15970
rect 57295 15752 57381 15808
rect 57437 15752 57593 15808
rect 57649 15752 57736 15808
rect 57295 15590 57736 15752
rect 57295 15534 57381 15590
rect 57437 15534 57593 15590
rect 57649 15534 57736 15590
rect 57295 15372 57736 15534
rect 57295 15316 57381 15372
rect 57437 15316 57593 15372
rect 57649 15316 57736 15372
rect 57295 15155 57736 15316
rect 57295 15099 57381 15155
rect 57437 15099 57593 15155
rect 57649 15099 57736 15155
rect 57295 14937 57736 15099
rect 57295 14881 57381 14937
rect 57437 14881 57593 14937
rect 57649 14881 57736 14937
rect 57295 14720 57736 14881
rect 57295 14664 57381 14720
rect 57437 14664 57593 14720
rect 57649 14664 57736 14720
rect 57295 14498 57736 14664
rect 57295 14446 57383 14498
rect 57435 14446 57595 14498
rect 57647 14446 57736 14498
rect 57295 14281 57736 14446
rect 57295 14229 57383 14281
rect 57435 14229 57595 14281
rect 57647 14229 57736 14281
rect 57295 14063 57736 14229
rect 57295 14011 57383 14063
rect 57435 14011 57595 14063
rect 57647 14011 57736 14063
rect 57295 13845 57736 14011
rect 57295 13793 57383 13845
rect 57435 13793 57595 13845
rect 57647 13793 57736 13845
rect 57295 13628 57736 13793
rect 57295 13576 57383 13628
rect 57435 13576 57595 13628
rect 57647 13576 57736 13628
rect 57295 13410 57736 13576
rect 57295 13358 57383 13410
rect 57435 13358 57595 13410
rect 57647 13358 57736 13410
rect 57295 13192 57736 13358
rect 57295 13140 57383 13192
rect 57435 13140 57595 13192
rect 57647 13140 57736 13192
rect 57295 12975 57736 13140
rect 57295 12923 57383 12975
rect 57435 12923 57595 12975
rect 57647 12923 57736 12975
rect 57295 12757 57736 12923
rect 57295 12705 57383 12757
rect 57435 12705 57595 12757
rect 57647 12705 57736 12757
rect 57295 12540 57736 12705
rect 57295 12488 57383 12540
rect 57435 12488 57595 12540
rect 57647 12488 57736 12540
rect 57295 12322 57736 12488
rect 57295 12270 57383 12322
rect 57435 12270 57595 12322
rect 57647 12270 57736 12322
rect 57295 12104 57736 12270
rect 57295 12052 57383 12104
rect 57435 12052 57595 12104
rect 57647 12052 57736 12104
rect 57295 11887 57736 12052
rect 57295 11835 57383 11887
rect 57435 11835 57595 11887
rect 57647 11835 57736 11887
rect 57295 11669 57736 11835
rect 57295 11617 57383 11669
rect 57435 11617 57595 11669
rect 57647 11617 57736 11669
rect 57295 11451 57736 11617
rect 57295 11406 57383 11451
rect 57435 11406 57595 11451
rect 57647 11406 57736 11451
rect 57295 11350 57381 11406
rect 57437 11350 57593 11406
rect 57649 11350 57736 11406
rect 57295 11234 57736 11350
rect 57295 11189 57383 11234
rect 57435 11189 57595 11234
rect 57647 11189 57736 11234
rect 57295 11133 57381 11189
rect 57437 11133 57593 11189
rect 57649 11133 57736 11189
rect 57295 11016 57736 11133
rect 57295 10971 57383 11016
rect 57435 10971 57595 11016
rect 57647 10971 57736 11016
rect 57295 10915 57381 10971
rect 57437 10915 57593 10971
rect 57649 10915 57736 10971
rect 57295 10798 57736 10915
rect 57295 10753 57383 10798
rect 57435 10753 57595 10798
rect 57647 10753 57736 10798
rect 57295 10697 57381 10753
rect 57437 10697 57593 10753
rect 57649 10697 57736 10753
rect 57295 10581 57736 10697
rect 57295 10535 57383 10581
rect 57435 10535 57595 10581
rect 57647 10535 57736 10581
rect 57295 10479 57381 10535
rect 57437 10479 57593 10535
rect 57649 10479 57736 10535
rect 57295 10363 57736 10479
rect 57295 10318 57383 10363
rect 57435 10318 57595 10363
rect 57647 10318 57736 10363
rect 57295 10262 57381 10318
rect 57437 10262 57593 10318
rect 57649 10262 57736 10318
rect 57295 10146 57736 10262
rect 57295 10094 57383 10146
rect 57435 10094 57595 10146
rect 57647 10094 57736 10146
rect 27387 9876 27476 9928
rect 27528 9876 27688 9928
rect 27740 9876 27828 9928
rect 27387 9710 27828 9876
rect 51756 9971 51832 9981
rect 51756 9811 51766 9971
rect 51822 9811 51832 9971
rect 51756 9801 51832 9811
rect 57295 9928 57736 10094
rect 57295 9876 57383 9928
rect 57435 9876 57595 9928
rect 57647 9876 57736 9928
rect 27387 9658 27476 9710
rect 27528 9658 27688 9710
rect 27740 9658 27828 9710
rect 27387 9493 27828 9658
rect 27387 9441 27476 9493
rect 27528 9441 27688 9493
rect 27740 9441 27828 9493
rect 27387 9275 27828 9441
rect 27387 9223 27476 9275
rect 27528 9223 27688 9275
rect 27740 9223 27828 9275
rect 27387 9057 27828 9223
rect 27387 9005 27476 9057
rect 27528 9005 27688 9057
rect 27740 9005 27828 9057
rect 27387 8840 27828 9005
rect 49896 8953 50076 8963
rect 49896 8897 49906 8953
rect 50066 8897 50076 8953
rect 49896 8887 50076 8897
rect 27387 8788 27476 8840
rect 27528 8788 27688 8840
rect 27740 8788 27828 8840
rect 27387 8622 27828 8788
rect 27387 8570 27476 8622
rect 27528 8570 27688 8622
rect 27740 8570 27828 8622
rect 27387 8404 27828 8570
rect 27387 8352 27476 8404
rect 27528 8352 27688 8404
rect 27740 8352 27828 8404
rect 27387 8187 27828 8352
rect 27387 8135 27476 8187
rect 27528 8135 27688 8187
rect 27740 8135 27828 8187
rect 27387 7969 27828 8135
rect 27387 7917 27476 7969
rect 27528 7917 27688 7969
rect 27740 7917 27828 7969
rect 27387 7752 27828 7917
rect 27387 7700 27476 7752
rect 27528 7700 27688 7752
rect 27740 7700 27828 7752
rect 27387 7535 27828 7700
rect 27387 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 27387 7317 27828 7479
rect 27387 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 27387 7099 27828 7261
rect 27387 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 27387 6881 27828 7043
rect 27387 6829 27476 6881
rect 27528 6829 27688 6881
rect 27740 6829 27828 6881
rect 27387 6663 27828 6829
rect 27387 6611 27476 6663
rect 27528 6611 27688 6663
rect 27740 6611 27828 6663
rect 27387 6446 27828 6611
rect 27387 6394 27476 6446
rect 27528 6394 27688 6446
rect 27740 6394 27828 6446
rect 27387 6228 27828 6394
rect 28237 6836 28999 6874
rect 28237 6780 28273 6836
rect 28329 6780 28484 6836
rect 28540 6780 28696 6836
rect 28752 6780 28907 6836
rect 28963 6780 28999 6836
rect 28237 6618 28999 6780
rect 28237 6562 28273 6618
rect 28329 6562 28484 6618
rect 28540 6562 28696 6618
rect 28752 6562 28907 6618
rect 28963 6562 28999 6618
rect 28237 6400 28999 6562
rect 28237 6344 28273 6400
rect 28329 6344 28484 6400
rect 28540 6344 28696 6400
rect 28752 6344 28907 6400
rect 28963 6344 28999 6400
rect 49958 6361 50014 8887
rect 28237 6306 28999 6344
rect 49896 6349 50076 6361
rect 49896 6297 49908 6349
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 27387 6176 27476 6228
rect 27528 6176 27688 6228
rect 27740 6176 27828 6228
rect 27387 6120 27828 6176
rect 27387 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 27828 6120
rect 27387 6011 27828 6064
rect 27387 5959 27476 6011
rect 27528 5959 27688 6011
rect 27740 5959 27828 6011
rect 27387 5902 27828 5959
rect 27387 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 27828 5902
rect 27387 5793 27828 5846
rect 27387 5741 27476 5793
rect 27528 5741 27688 5793
rect 27740 5741 27828 5793
rect 27387 5575 27828 5741
rect 27387 5523 27476 5575
rect 27528 5523 27688 5575
rect 27740 5523 27828 5575
rect 27387 5358 27828 5523
rect 27387 5306 27476 5358
rect 27528 5306 27688 5358
rect 27740 5306 27828 5358
rect 1864 5024 2509 5135
rect 11727 5073 11783 5140
rect 1864 0 2088 5024
rect 3263 5001 3357 5062
rect 11617 5017 11783 5073
rect 3263 4880 3539 5001
rect 3445 1701 3539 4880
rect 11617 1701 11673 5017
rect 12575 4740 12631 5185
rect 12290 4684 12631 4740
rect 13253 4740 13309 5185
rect 14101 5073 14157 5140
rect 14101 5017 14267 5073
rect 13253 4684 13594 4740
rect 12290 1701 12346 4684
rect 13538 1701 13594 4684
rect 14211 1701 14267 5017
rect 22527 5001 22621 5062
rect 23375 5024 23953 5135
rect 22345 4880 22621 5001
rect 22345 1701 22439 4880
rect 23859 1701 23953 5024
rect 26823 4587 27163 4628
rect 26823 4535 26861 4587
rect 26913 4535 27073 4587
rect 27125 4535 27163 4587
rect 26823 4528 27163 4535
rect 26823 4472 26859 4528
rect 26915 4472 27071 4528
rect 27127 4472 27163 4528
rect 26823 4370 27163 4472
rect 26823 4318 26861 4370
rect 26913 4318 27073 4370
rect 27125 4318 27163 4370
rect 26823 4310 27163 4318
rect 26823 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 27163 4310
rect 26823 4152 27163 4254
rect 26823 4100 26861 4152
rect 26913 4100 27073 4152
rect 27125 4100 27163 4152
rect 26823 3934 27163 4100
rect 26823 3882 26861 3934
rect 26913 3882 27073 3934
rect 27125 3882 27163 3934
rect 26823 3717 27163 3882
rect 26823 3665 26861 3717
rect 26913 3665 27073 3717
rect 27125 3665 27163 3717
rect 26823 3624 27163 3665
rect 27387 4587 27828 5306
rect 27387 4535 27476 4587
rect 27528 4535 27688 4587
rect 27740 4535 27828 4587
rect 27387 4370 27828 4535
rect 27387 4318 27476 4370
rect 27528 4318 27688 4370
rect 27740 4318 27828 4370
rect 27387 4152 27828 4318
rect 27387 4100 27476 4152
rect 27528 4100 27688 4152
rect 27740 4100 27828 4152
rect 27387 3934 27828 4100
rect 27387 3882 27476 3934
rect 27528 3882 27688 3934
rect 27740 3882 27828 3934
rect 27387 3837 27828 3882
rect 27387 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 27828 3837
rect 27387 3717 27828 3781
rect 27387 3665 27476 3717
rect 27528 3665 27688 3717
rect 27740 3665 27828 3717
rect 27387 3619 27828 3665
rect 27387 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 27828 3619
rect 27387 3524 27828 3563
rect 28764 3837 28894 3876
rect 28764 3781 28801 3837
rect 28857 3781 28894 3837
rect 28764 3619 28894 3781
rect 28764 3563 28801 3619
rect 28857 3563 28894 3619
rect 28764 3525 28894 3563
rect 2539 1689 2763 1701
rect 2539 1637 2574 1689
rect 2730 1637 2763 1689
rect 2539 0 2763 1637
rect 3380 0 3604 1701
rect 11533 0 11757 1701
rect 12206 0 12430 1701
rect 12604 1689 12828 1701
rect 12604 1637 12639 1689
rect 12795 1637 12828 1689
rect 12604 0 12828 1637
rect 13054 1689 13278 1701
rect 13054 1637 13089 1689
rect 13245 1637 13278 1689
rect 13054 0 13278 1637
rect 13454 0 13678 1701
rect 14127 0 14351 1701
rect 22279 0 22503 1701
rect 23404 1689 23628 1701
rect 23404 1637 23439 1689
rect 23595 1637 23628 1689
rect 23404 0 23628 1637
rect 23795 0 24019 1701
rect 27936 0 28160 3418
rect 29006 2990 29135 3418
rect 29247 3243 29929 3418
rect 29006 917 29230 2990
rect 29006 657 29092 917
rect 29144 657 29230 917
rect 29006 0 29230 657
rect 29705 0 29929 3243
rect 30859 0 31083 6229
rect 32552 0 32776 6229
rect 34243 0 34467 6229
rect 40588 3282 40812 3294
rect 40588 3230 40623 3282
rect 40779 3230 40812 3282
rect 40588 0 40812 3230
rect 43790 3044 43970 3054
rect 43790 2988 43800 3044
rect 43960 2988 43970 3044
rect 43790 2978 43970 2988
rect 50342 0 50566 7745
rect 51766 5211 51822 9801
rect 57295 9710 57736 9876
rect 57295 9658 57383 9710
rect 57435 9658 57595 9710
rect 57647 9658 57736 9710
rect 57295 9493 57736 9658
rect 57295 9441 57383 9493
rect 57435 9441 57595 9493
rect 57647 9441 57736 9493
rect 57295 9275 57736 9441
rect 57295 9223 57383 9275
rect 57435 9223 57595 9275
rect 57647 9223 57736 9275
rect 57295 9057 57736 9223
rect 57295 9005 57383 9057
rect 57435 9005 57595 9057
rect 57647 9005 57736 9057
rect 57295 8854 57736 9005
rect 57295 8798 57381 8854
rect 57437 8798 57593 8854
rect 57649 8798 57736 8854
rect 57295 8788 57383 8798
rect 57435 8788 57595 8798
rect 57647 8788 57736 8798
rect 57295 8636 57736 8788
rect 57295 8580 57381 8636
rect 57437 8580 57593 8636
rect 57649 8580 57736 8636
rect 57295 8570 57383 8580
rect 57435 8570 57595 8580
rect 57647 8570 57736 8580
rect 57295 8419 57736 8570
rect 57295 8363 57381 8419
rect 57437 8363 57593 8419
rect 57649 8363 57736 8419
rect 57295 8352 57383 8363
rect 57435 8352 57595 8363
rect 57647 8352 57736 8363
rect 57295 8201 57736 8352
rect 57295 8145 57381 8201
rect 57437 8145 57593 8201
rect 57649 8145 57736 8201
rect 57295 8135 57383 8145
rect 57435 8135 57595 8145
rect 57647 8135 57736 8145
rect 57295 7983 57736 8135
rect 57295 7927 57381 7983
rect 57437 7927 57593 7983
rect 57649 7927 57736 7983
rect 57295 7917 57383 7927
rect 57435 7917 57595 7927
rect 57647 7917 57736 7927
rect 57295 7766 57736 7917
rect 57295 7710 57381 7766
rect 57437 7710 57593 7766
rect 57649 7710 57736 7766
rect 57295 7700 57383 7710
rect 57435 7700 57595 7710
rect 57647 7700 57736 7710
rect 57295 7548 57736 7700
rect 57295 7492 57381 7548
rect 57437 7492 57593 7548
rect 57649 7492 57736 7548
rect 57295 7482 57383 7492
rect 57435 7482 57595 7492
rect 57647 7482 57736 7492
rect 57295 7330 57736 7482
rect 57295 7274 57381 7330
rect 57437 7274 57593 7330
rect 57649 7274 57736 7330
rect 57295 7264 57383 7274
rect 57435 7264 57595 7274
rect 57647 7264 57736 7274
rect 57295 7113 57736 7264
rect 57295 7057 57381 7113
rect 57437 7057 57593 7113
rect 57649 7057 57736 7113
rect 57295 7047 57383 7057
rect 57435 7047 57595 7057
rect 57647 7047 57736 7057
rect 57295 6881 57736 7047
rect 56124 6836 56886 6874
rect 56124 6780 56160 6836
rect 56216 6780 56371 6836
rect 56427 6780 56583 6836
rect 56639 6780 56794 6836
rect 56850 6780 56886 6836
rect 56124 6618 56886 6780
rect 56124 6562 56160 6618
rect 56216 6562 56371 6618
rect 56427 6562 56583 6618
rect 56639 6562 56794 6618
rect 56850 6562 56886 6618
rect 56124 6400 56886 6562
rect 56124 6344 56160 6400
rect 56216 6344 56371 6400
rect 56427 6344 56583 6400
rect 56639 6344 56794 6400
rect 56850 6344 56886 6400
rect 56124 6306 56886 6344
rect 57295 6829 57383 6881
rect 57435 6829 57595 6881
rect 57647 6829 57736 6881
rect 57295 6663 57736 6829
rect 57295 6611 57383 6663
rect 57435 6611 57595 6663
rect 57647 6611 57736 6663
rect 57295 6446 57736 6611
rect 57295 6394 57383 6446
rect 57435 6394 57595 6446
rect 57647 6394 57736 6446
rect 51642 5199 51822 5211
rect 51642 5147 51654 5199
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 57295 6228 57736 6394
rect 57295 6176 57383 6228
rect 57435 6176 57595 6228
rect 57647 6176 57736 6228
rect 57295 6120 57736 6176
rect 57295 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 57736 6120
rect 57295 6011 57736 6064
rect 57295 5959 57383 6011
rect 57435 5959 57595 6011
rect 57647 5959 57736 6011
rect 57295 5902 57736 5959
rect 57295 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 57736 5902
rect 57295 5793 57736 5846
rect 57295 5741 57383 5793
rect 57435 5741 57595 5793
rect 57647 5741 57736 5793
rect 57295 5575 57736 5741
rect 57295 5523 57383 5575
rect 57435 5523 57595 5575
rect 57647 5523 57736 5575
rect 57295 5358 57736 5523
rect 57295 5306 57383 5358
rect 57435 5306 57595 5358
rect 57647 5306 57736 5358
rect 57295 4587 57736 5306
rect 57295 4535 57383 4587
rect 57435 4535 57595 4587
rect 57647 4535 57736 4587
rect 57295 4370 57736 4535
rect 57295 4318 57383 4370
rect 57435 4318 57595 4370
rect 57647 4318 57736 4370
rect 57295 4152 57736 4318
rect 57295 4100 57383 4152
rect 57435 4100 57595 4152
rect 57647 4100 57736 4152
rect 57295 3934 57736 4100
rect 55540 3309 55669 3891
rect 57295 3882 57383 3934
rect 57435 3882 57595 3934
rect 57647 3882 57736 3934
rect 57295 3837 57736 3882
rect 57295 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 57736 3837
rect 57295 3717 57736 3781
rect 57295 3665 57383 3717
rect 57435 3665 57595 3717
rect 57647 3665 57736 3717
rect 57295 3619 57736 3665
rect 57295 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 57736 3619
rect 57295 3524 57736 3563
rect 57909 33432 58351 33520
rect 57909 33380 57998 33432
rect 58050 33380 58210 33432
rect 58262 33380 58351 33432
rect 57909 33358 58351 33380
rect 57909 33302 57996 33358
rect 58052 33302 58208 33358
rect 58264 33302 58351 33358
rect 57909 33215 58351 33302
rect 57909 33163 57998 33215
rect 58050 33163 58210 33215
rect 58262 33163 58351 33215
rect 57909 33140 58351 33163
rect 57909 33084 57996 33140
rect 58052 33084 58208 33140
rect 58264 33084 58351 33140
rect 57909 32997 58351 33084
rect 57909 32945 57998 32997
rect 58050 32945 58210 32997
rect 58262 32945 58351 32997
rect 57909 32922 58351 32945
rect 57909 32866 57996 32922
rect 58052 32866 58208 32922
rect 58264 32866 58351 32922
rect 57909 32779 58351 32866
rect 57909 32727 57998 32779
rect 58050 32727 58210 32779
rect 58262 32727 58351 32779
rect 57909 32705 58351 32727
rect 57909 32649 57996 32705
rect 58052 32649 58208 32705
rect 58264 32649 58351 32705
rect 57909 32562 58351 32649
rect 57909 32510 57998 32562
rect 58050 32510 58210 32562
rect 58262 32510 58351 32562
rect 57909 32487 58351 32510
rect 57909 32431 57996 32487
rect 58052 32431 58208 32487
rect 58264 32431 58351 32487
rect 57909 32344 58351 32431
rect 57909 32292 57998 32344
rect 58050 32292 58210 32344
rect 58262 32292 58351 32344
rect 57909 32127 58351 32292
rect 57909 32088 57998 32127
rect 58050 32088 58210 32127
rect 58262 32088 58351 32127
rect 57909 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 57909 31909 58351 32032
rect 57909 31870 57998 31909
rect 58050 31870 58210 31909
rect 58262 31870 58351 31909
rect 57909 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 57909 31691 58351 31814
rect 57909 31652 57998 31691
rect 58050 31652 58210 31691
rect 58262 31652 58351 31691
rect 57909 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 57909 31474 58351 31596
rect 57909 31422 57998 31474
rect 58050 31422 58210 31474
rect 58262 31422 58351 31474
rect 57909 31256 58351 31422
rect 57909 31204 57998 31256
rect 58050 31204 58210 31256
rect 58262 31204 58351 31256
rect 57909 31038 58351 31204
rect 57909 30986 57998 31038
rect 58050 30986 58210 31038
rect 58262 30986 58351 31038
rect 57909 30821 58351 30986
rect 57909 30769 57998 30821
rect 58050 30769 58210 30821
rect 58262 30769 58351 30821
rect 57909 30603 58351 30769
rect 57909 30551 57998 30603
rect 58050 30551 58210 30603
rect 58262 30551 58351 30603
rect 57909 30386 58351 30551
rect 57909 30334 57998 30386
rect 58050 30334 58210 30386
rect 58262 30334 58351 30386
rect 57909 30168 58351 30334
rect 57909 30116 57998 30168
rect 58050 30116 58210 30168
rect 58262 30116 58351 30168
rect 57909 29968 58351 30116
rect 57909 29912 57996 29968
rect 58052 29912 58208 29968
rect 58264 29912 58351 29968
rect 57909 29898 57998 29912
rect 58050 29898 58210 29912
rect 58262 29898 58351 29912
rect 57909 29750 58351 29898
rect 57909 29694 57996 29750
rect 58052 29694 58208 29750
rect 58264 29694 58351 29750
rect 57909 29681 57998 29694
rect 58050 29681 58210 29694
rect 58262 29681 58351 29694
rect 57909 29533 58351 29681
rect 57909 29477 57996 29533
rect 58052 29477 58208 29533
rect 58264 29477 58351 29533
rect 57909 29463 57998 29477
rect 58050 29463 58210 29477
rect 58262 29463 58351 29477
rect 57909 29315 58351 29463
rect 57909 29259 57996 29315
rect 58052 29259 58208 29315
rect 58264 29259 58351 29315
rect 57909 29245 57998 29259
rect 58050 29245 58210 29259
rect 58262 29245 58351 29259
rect 57909 29098 58351 29245
rect 57909 29042 57996 29098
rect 58052 29042 58208 29098
rect 58264 29042 58351 29098
rect 57909 29028 57998 29042
rect 58050 29028 58210 29042
rect 58262 29028 58351 29042
rect 57909 28880 58351 29028
rect 57909 28824 57996 28880
rect 58052 28824 58208 28880
rect 58264 28824 58351 28880
rect 57909 28810 57998 28824
rect 58050 28810 58210 28824
rect 58262 28810 58351 28824
rect 57909 28662 58351 28810
rect 57909 28606 57996 28662
rect 58052 28606 58208 28662
rect 58264 28606 58351 28662
rect 57909 28592 57998 28606
rect 58050 28592 58210 28606
rect 58262 28592 58351 28606
rect 57909 28444 58351 28592
rect 57909 28388 57996 28444
rect 58052 28388 58208 28444
rect 58264 28388 58351 28444
rect 57909 28375 57998 28388
rect 58050 28375 58210 28388
rect 58262 28375 58351 28388
rect 57909 28227 58351 28375
rect 57909 28171 57996 28227
rect 58052 28171 58208 28227
rect 58264 28171 58351 28227
rect 57909 28157 57998 28171
rect 58050 28157 58210 28171
rect 58262 28157 58351 28171
rect 57909 28009 58351 28157
rect 57909 27953 57996 28009
rect 58052 27953 58208 28009
rect 58264 27953 58351 28009
rect 57909 27940 57998 27953
rect 58050 27940 58210 27953
rect 58262 27940 58351 27953
rect 57909 27792 58351 27940
rect 57909 27736 57996 27792
rect 58052 27736 58208 27792
rect 58264 27736 58351 27792
rect 57909 27722 57998 27736
rect 58050 27722 58210 27736
rect 58262 27722 58351 27736
rect 57909 27574 58351 27722
rect 57909 27518 57996 27574
rect 58052 27518 58208 27574
rect 58264 27518 58351 27574
rect 57909 27504 57998 27518
rect 58050 27504 58210 27518
rect 58262 27504 58351 27518
rect 57909 27339 58351 27504
rect 57909 27287 57998 27339
rect 58050 27287 58210 27339
rect 58262 27287 58351 27339
rect 57909 27121 58351 27287
rect 57909 27069 57998 27121
rect 58050 27069 58210 27121
rect 58262 27069 58351 27121
rect 57909 26903 58351 27069
rect 57909 26851 57998 26903
rect 58050 26851 58210 26903
rect 58262 26851 58351 26903
rect 57909 26686 58351 26851
rect 57909 26634 57998 26686
rect 58050 26634 58210 26686
rect 58262 26634 58351 26686
rect 57909 26468 58351 26634
rect 57909 26416 57998 26468
rect 58050 26416 58210 26468
rect 58262 26416 58351 26468
rect 58791 65916 59517 65955
rect 58791 65860 58856 65916
rect 58912 65860 58980 65916
rect 59036 65860 59104 65916
rect 59160 65860 59228 65916
rect 59284 65860 59352 65916
rect 59408 65860 59517 65916
rect 58791 65792 59517 65860
rect 58791 65736 58856 65792
rect 58912 65736 58980 65792
rect 59036 65736 59104 65792
rect 59160 65736 59228 65792
rect 59284 65736 59352 65792
rect 59408 65736 59517 65792
rect 58791 34981 59517 65736
rect 58791 34925 58822 34981
rect 58878 34925 58946 34981
rect 59002 34925 59070 34981
rect 59126 34925 59194 34981
rect 59250 34925 59318 34981
rect 59374 34925 59442 34981
rect 59498 34925 59517 34981
rect 58791 34857 59517 34925
rect 58791 34801 58822 34857
rect 58878 34801 58946 34857
rect 59002 34801 59070 34857
rect 59126 34801 59194 34857
rect 59250 34801 59318 34857
rect 59374 34801 59442 34857
rect 59498 34801 59517 34857
rect 58791 34733 59517 34801
rect 58791 34677 58822 34733
rect 58878 34677 58946 34733
rect 59002 34677 59070 34733
rect 59126 34677 59194 34733
rect 59250 34677 59318 34733
rect 59374 34677 59442 34733
rect 59498 34677 59517 34733
rect 58791 31298 59517 34677
rect 58791 31242 58873 31298
rect 58929 31242 58997 31298
rect 59053 31242 59121 31298
rect 59177 31242 59245 31298
rect 59301 31242 59369 31298
rect 59425 31242 59517 31298
rect 58791 31174 59517 31242
rect 58791 31118 58873 31174
rect 58929 31118 58997 31174
rect 59053 31118 59121 31174
rect 59177 31118 59245 31174
rect 59301 31118 59369 31174
rect 59425 31118 59517 31174
rect 58791 31050 59517 31118
rect 58791 30994 58873 31050
rect 58929 30994 58997 31050
rect 59053 30994 59121 31050
rect 59177 30994 59245 31050
rect 59301 30994 59369 31050
rect 59425 30994 59517 31050
rect 58791 30853 59517 30994
rect 58791 30797 58873 30853
rect 58929 30797 58997 30853
rect 59053 30797 59121 30853
rect 59177 30797 59245 30853
rect 59301 30797 59369 30853
rect 59425 30797 59517 30853
rect 58791 30729 59517 30797
rect 58791 30673 58873 30729
rect 58929 30673 58997 30729
rect 59053 30673 59121 30729
rect 59177 30673 59245 30729
rect 59301 30673 59369 30729
rect 59425 30673 59517 30729
rect 58791 30605 59517 30673
rect 58791 30549 58873 30605
rect 58929 30549 58997 30605
rect 59053 30549 59121 30605
rect 59177 30549 59245 30605
rect 59301 30549 59369 30605
rect 59425 30549 59517 30605
rect 58791 28321 59517 30549
rect 58791 28265 58859 28321
rect 58915 28265 58983 28321
rect 59039 28265 59107 28321
rect 59163 28265 59231 28321
rect 59287 28265 59355 28321
rect 59411 28265 59517 28321
rect 58791 28197 59517 28265
rect 58791 28141 58859 28197
rect 58915 28141 58983 28197
rect 59039 28141 59107 28197
rect 59163 28141 59231 28197
rect 59287 28141 59355 28197
rect 59411 28141 59517 28197
rect 58791 28073 59517 28141
rect 58791 28017 58859 28073
rect 58915 28017 58983 28073
rect 59039 28017 59107 28073
rect 59163 28017 59231 28073
rect 59287 28017 59355 28073
rect 59411 28017 59517 28073
rect 58791 27949 59517 28017
rect 58791 27893 58859 27949
rect 58915 27893 58983 27949
rect 59039 27893 59107 27949
rect 59163 27893 59231 27949
rect 59287 27893 59355 27949
rect 59411 27893 59517 27949
rect 58791 27825 59517 27893
rect 58791 27769 58859 27825
rect 58915 27769 58983 27825
rect 59039 27769 59107 27825
rect 59163 27769 59231 27825
rect 59287 27769 59355 27825
rect 59411 27769 59517 27825
rect 58791 27701 59517 27769
rect 58791 27645 58859 27701
rect 58915 27645 58983 27701
rect 59039 27645 59107 27701
rect 59163 27645 59231 27701
rect 59287 27645 59355 27701
rect 59411 27645 59517 27701
rect 58791 27577 59517 27645
rect 58791 27521 58859 27577
rect 58915 27521 58983 27577
rect 59039 27521 59107 27577
rect 59163 27521 59231 27577
rect 59287 27521 59355 27577
rect 59411 27521 59517 27577
rect 58791 27453 59517 27521
rect 58791 27397 58859 27453
rect 58915 27397 58983 27453
rect 59039 27397 59107 27453
rect 59163 27397 59231 27453
rect 59287 27397 59355 27453
rect 59411 27397 59517 27453
rect 58791 27329 59517 27397
rect 58791 27273 58859 27329
rect 58915 27273 58983 27329
rect 59039 27273 59107 27329
rect 59163 27273 59231 27329
rect 59287 27273 59355 27329
rect 59411 27273 59517 27329
rect 58791 27205 59517 27273
rect 58791 27149 58859 27205
rect 58915 27149 58983 27205
rect 59039 27149 59107 27205
rect 59163 27149 59231 27205
rect 59287 27149 59355 27205
rect 59411 27149 59517 27205
rect 58791 27081 59517 27149
rect 58791 27025 58859 27081
rect 58915 27025 58983 27081
rect 59039 27025 59107 27081
rect 59163 27025 59231 27081
rect 59287 27025 59355 27081
rect 59411 27025 59517 27081
rect 58791 26957 59517 27025
rect 58791 26901 58859 26957
rect 58915 26901 58983 26957
rect 59039 26901 59107 26957
rect 59163 26901 59231 26957
rect 59287 26901 59355 26957
rect 59411 26901 59517 26957
rect 58791 26833 59517 26901
rect 58791 26777 58859 26833
rect 58915 26777 58983 26833
rect 59039 26777 59107 26833
rect 59163 26777 59231 26833
rect 59287 26777 59355 26833
rect 59411 26777 59517 26833
rect 58791 26709 59517 26777
rect 58791 26653 58859 26709
rect 58915 26653 58983 26709
rect 59039 26653 59107 26709
rect 59163 26653 59231 26709
rect 59287 26653 59355 26709
rect 59411 26653 59517 26709
rect 58791 26585 59517 26653
rect 58791 26529 58859 26585
rect 58915 26529 58983 26585
rect 59039 26529 59107 26585
rect 59163 26529 59231 26585
rect 59287 26529 59355 26585
rect 59411 26529 59517 26585
rect 58791 26433 59517 26529
rect 57909 26250 58351 26416
rect 57909 26198 57998 26250
rect 58050 26198 58210 26250
rect 58262 26198 58351 26250
rect 57909 26033 58351 26198
rect 57909 25981 57998 26033
rect 58050 25981 58210 26033
rect 58262 25981 58351 26033
rect 57909 25815 58351 25981
rect 57909 25763 57998 25815
rect 58050 25763 58210 25815
rect 58262 25763 58351 25815
rect 57909 25598 58351 25763
rect 57909 25546 57998 25598
rect 58050 25546 58210 25598
rect 58262 25546 58351 25598
rect 57909 25380 58351 25546
rect 57909 25328 57998 25380
rect 58050 25328 58210 25380
rect 58262 25328 58351 25380
rect 57909 25162 58351 25328
rect 57909 25110 57998 25162
rect 58050 25110 58210 25162
rect 58262 25110 58351 25162
rect 57909 24945 58351 25110
rect 57909 24893 57998 24945
rect 58050 24893 58210 24945
rect 58262 24893 58351 24945
rect 57909 24727 58351 24893
rect 57909 24675 57998 24727
rect 58050 24675 58210 24727
rect 58262 24675 58351 24727
rect 57909 24509 58351 24675
rect 57909 24457 57998 24509
rect 58050 24457 58210 24509
rect 58262 24457 58351 24509
rect 57909 24292 58351 24457
rect 57909 24240 57998 24292
rect 58050 24240 58210 24292
rect 58262 24240 58351 24292
rect 57909 24075 58351 24240
rect 57909 23187 57994 24075
rect 58258 24074 58351 24075
rect 58262 24022 58351 24074
rect 58258 23857 58351 24022
rect 58262 23805 58351 23857
rect 58258 23639 58351 23805
rect 58262 23587 58351 23639
rect 58258 23421 58351 23587
rect 58262 23369 58351 23421
rect 58258 23204 58351 23369
rect 57909 23152 57998 23187
rect 58050 23152 58210 23187
rect 58262 23152 58351 23204
rect 57909 22986 58351 23152
rect 57909 22934 57998 22986
rect 58050 22934 58210 22986
rect 58262 22934 58351 22986
rect 57909 22768 58351 22934
rect 57909 22716 57998 22768
rect 58050 22716 58210 22768
rect 58262 22716 58351 22768
rect 57909 22551 58351 22716
rect 57909 22499 57998 22551
rect 58050 22499 58210 22551
rect 58262 22499 58351 22551
rect 57909 22333 58351 22499
rect 57909 22281 57998 22333
rect 58050 22281 58210 22333
rect 58262 22281 58351 22333
rect 57909 22115 58351 22281
rect 57909 22063 57998 22115
rect 58050 22063 58210 22115
rect 58262 22063 58351 22115
rect 57909 21898 58351 22063
rect 57909 21846 57998 21898
rect 58050 21846 58210 21898
rect 58262 21846 58351 21898
rect 57909 21680 58351 21846
rect 57909 21628 57998 21680
rect 58050 21628 58210 21680
rect 58262 21628 58351 21680
rect 57909 21463 58351 21628
rect 57909 21411 57998 21463
rect 58050 21411 58210 21463
rect 58262 21411 58351 21463
rect 57909 21245 58351 21411
rect 57909 21193 57998 21245
rect 58050 21193 58210 21245
rect 58262 21193 58351 21245
rect 57909 21027 58351 21193
rect 57909 20975 57998 21027
rect 58050 20975 58210 21027
rect 58262 20975 58351 21027
rect 57909 20810 58351 20975
rect 57909 20758 57998 20810
rect 58050 20758 58210 20810
rect 58262 20758 58351 20810
rect 57909 20592 58351 20758
rect 57909 20540 57998 20592
rect 58050 20570 58210 20592
rect 58208 20540 58210 20570
rect 58262 20540 58351 20592
rect 57909 20410 58048 20540
rect 58208 20410 58351 20540
rect 57909 20374 58351 20410
rect 57909 20322 57998 20374
rect 58050 20322 58210 20374
rect 58262 20322 58351 20374
rect 57909 20226 58351 20322
rect 57909 20157 58048 20226
rect 58208 20157 58351 20226
rect 57909 20105 57998 20157
rect 58208 20105 58210 20157
rect 58262 20105 58351 20157
rect 57909 20066 58048 20105
rect 58208 20066 58351 20105
rect 57909 19939 58351 20066
rect 57909 19887 57998 19939
rect 58050 19887 58210 19939
rect 58262 19887 58351 19939
rect 57909 19722 58351 19887
rect 57909 19670 57998 19722
rect 58050 19670 58210 19722
rect 58262 19670 58351 19722
rect 57909 19504 58351 19670
rect 57909 19452 57998 19504
rect 58050 19452 58210 19504
rect 58262 19452 58351 19504
rect 57909 19286 58351 19452
rect 57909 19234 57998 19286
rect 58050 19234 58210 19286
rect 58262 19234 58351 19286
rect 57909 19068 58351 19234
rect 57909 19016 57998 19068
rect 58050 19016 58210 19068
rect 58262 19016 58351 19068
rect 57909 18851 58351 19016
rect 57909 18799 57998 18851
rect 58050 18799 58210 18851
rect 58262 18799 58351 18851
rect 57909 18633 58351 18799
rect 57909 18581 57998 18633
rect 58050 18581 58210 18633
rect 58262 18581 58351 18633
rect 57909 18416 58351 18581
rect 57909 18364 57998 18416
rect 58050 18364 58210 18416
rect 58262 18364 58351 18416
rect 57909 18198 58351 18364
rect 57909 18146 57998 18198
rect 58050 18146 58210 18198
rect 58262 18146 58351 18198
rect 57909 17980 58351 18146
rect 57909 17928 57998 17980
rect 58050 17928 58210 17980
rect 58262 17928 58351 17980
rect 57909 17763 58351 17928
rect 57909 17711 57998 17763
rect 58050 17711 58210 17763
rect 58262 17711 58351 17763
rect 57909 17545 58351 17711
rect 57909 17493 57998 17545
rect 58050 17493 58210 17545
rect 58262 17493 58351 17545
rect 57909 17327 58351 17493
rect 57909 17275 57998 17327
rect 58050 17275 58210 17327
rect 58262 17275 58351 17327
rect 57909 17110 58351 17275
rect 57909 17058 57998 17110
rect 58050 17058 58210 17110
rect 58262 17058 58351 17110
rect 57909 16892 58351 17058
rect 57909 16840 57998 16892
rect 58050 16840 58210 16892
rect 58262 16840 58351 16892
rect 57909 16675 58351 16840
rect 57909 16623 57998 16675
rect 58050 16623 58210 16675
rect 58262 16623 58351 16675
rect 57909 16457 58351 16623
rect 57909 16405 57998 16457
rect 58050 16405 58210 16457
rect 58262 16405 58351 16457
rect 57909 16239 58351 16405
rect 57909 16187 57998 16239
rect 58050 16187 58210 16239
rect 58262 16187 58351 16239
rect 57909 16022 58351 16187
rect 57909 15970 57998 16022
rect 58050 15970 58210 16022
rect 58262 15970 58351 16022
rect 57909 15804 58351 15970
rect 57909 15752 57998 15804
rect 58050 15752 58210 15804
rect 58262 15752 58351 15804
rect 57909 15586 58351 15752
rect 57909 15534 57998 15586
rect 58050 15534 58210 15586
rect 58262 15534 58351 15586
rect 57909 15369 58351 15534
rect 57909 15317 57998 15369
rect 58050 15317 58210 15369
rect 58262 15317 58351 15369
rect 57909 15151 58351 15317
rect 57909 15099 57998 15151
rect 58050 15099 58210 15151
rect 58262 15099 58351 15151
rect 57909 14933 58351 15099
rect 57909 14881 57998 14933
rect 58050 14881 58210 14933
rect 58262 14881 58351 14933
rect 57909 14716 58351 14881
rect 57909 14664 57998 14716
rect 58050 14664 58210 14716
rect 58262 14664 58351 14716
rect 57909 14498 58351 14664
rect 57909 14446 57998 14498
rect 58050 14446 58210 14498
rect 58262 14446 58351 14498
rect 57909 14281 58351 14446
rect 57909 14229 57998 14281
rect 58050 14229 58210 14281
rect 58262 14229 58351 14281
rect 57909 14063 58351 14229
rect 57909 14011 57998 14063
rect 58050 14011 58210 14063
rect 58262 14011 58351 14063
rect 57909 13845 58351 14011
rect 57909 13793 57998 13845
rect 58050 13793 58210 13845
rect 58262 13793 58351 13845
rect 57909 13790 58351 13793
rect 57909 13734 57996 13790
rect 58052 13734 58208 13790
rect 58264 13734 58351 13790
rect 57909 13628 58351 13734
rect 57909 13576 57998 13628
rect 58050 13576 58210 13628
rect 58262 13576 58351 13628
rect 57909 13573 58351 13576
rect 57909 13517 57996 13573
rect 58052 13517 58208 13573
rect 58264 13517 58351 13573
rect 57909 13410 58351 13517
rect 57909 13358 57998 13410
rect 58050 13358 58210 13410
rect 58262 13358 58351 13410
rect 57909 13355 58351 13358
rect 57909 13299 57996 13355
rect 58052 13299 58208 13355
rect 58264 13299 58351 13355
rect 57909 13192 58351 13299
rect 57909 13140 57998 13192
rect 58050 13140 58210 13192
rect 58262 13140 58351 13192
rect 57909 13138 58351 13140
rect 57909 13082 57996 13138
rect 58052 13082 58208 13138
rect 58264 13082 58351 13138
rect 57909 12975 58351 13082
rect 57909 12923 57998 12975
rect 58050 12923 58210 12975
rect 58262 12923 58351 12975
rect 57909 12920 58351 12923
rect 57909 12864 57996 12920
rect 58052 12864 58208 12920
rect 58264 12864 58351 12920
rect 57909 12757 58351 12864
rect 57909 12705 57998 12757
rect 58050 12705 58210 12757
rect 58262 12705 58351 12757
rect 57909 12702 58351 12705
rect 57909 12646 57996 12702
rect 58052 12646 58208 12702
rect 58264 12646 58351 12702
rect 57909 12540 58351 12646
rect 57909 12488 57998 12540
rect 58050 12488 58210 12540
rect 58262 12488 58351 12540
rect 57909 12484 58351 12488
rect 57909 12428 57996 12484
rect 58052 12428 58208 12484
rect 58264 12428 58351 12484
rect 57909 12322 58351 12428
rect 57909 12270 57998 12322
rect 58050 12270 58210 12322
rect 58262 12270 58351 12322
rect 57909 12267 58351 12270
rect 57909 12211 57996 12267
rect 58052 12211 58208 12267
rect 58264 12211 58351 12267
rect 57909 12104 58351 12211
rect 57909 12052 57998 12104
rect 58050 12052 58210 12104
rect 58262 12052 58351 12104
rect 57909 12049 58351 12052
rect 57909 11993 57996 12049
rect 58052 11993 58208 12049
rect 58264 11993 58351 12049
rect 57909 11887 58351 11993
rect 57909 11835 57998 11887
rect 58050 11835 58210 11887
rect 58262 11835 58351 11887
rect 57909 11832 58351 11835
rect 57909 11776 57996 11832
rect 58052 11776 58208 11832
rect 58264 11776 58351 11832
rect 57909 11669 58351 11776
rect 57909 11617 57998 11669
rect 58050 11617 58210 11669
rect 58262 11617 58351 11669
rect 57909 11451 58351 11617
rect 57909 11399 57998 11451
rect 58050 11399 58210 11451
rect 58262 11399 58351 11451
rect 57909 11234 58351 11399
rect 57909 11182 57998 11234
rect 58050 11182 58210 11234
rect 58262 11182 58351 11234
rect 57909 11016 58351 11182
rect 57909 10964 57998 11016
rect 58050 10964 58210 11016
rect 58262 10964 58351 11016
rect 57909 10798 58351 10964
rect 57909 10746 57998 10798
rect 58050 10746 58210 10798
rect 58262 10746 58351 10798
rect 57909 10581 58351 10746
rect 57909 10529 57998 10581
rect 58050 10529 58210 10581
rect 58262 10529 58351 10581
rect 57909 10363 58351 10529
rect 57909 10311 57998 10363
rect 58050 10311 58210 10363
rect 58262 10311 58351 10363
rect 57909 10146 58351 10311
rect 57909 10094 57998 10146
rect 58050 10094 58210 10146
rect 58262 10094 58351 10146
rect 57909 9928 58351 10094
rect 57909 9876 57998 9928
rect 58050 9876 58210 9928
rect 58262 9876 58351 9928
rect 57909 9710 58351 9876
rect 57909 9658 57998 9710
rect 58050 9658 58210 9710
rect 58262 9658 58351 9710
rect 57909 9493 58351 9658
rect 57909 9441 57998 9493
rect 58050 9441 58210 9493
rect 58262 9441 58351 9493
rect 57909 9407 58351 9441
rect 57909 9351 57996 9407
rect 58052 9351 58208 9407
rect 58264 9351 58351 9407
rect 57909 9275 58351 9351
rect 57909 9223 57998 9275
rect 58050 9223 58210 9275
rect 58262 9223 58351 9275
rect 57909 9190 58351 9223
rect 57909 9134 57996 9190
rect 58052 9134 58208 9190
rect 58264 9134 58351 9190
rect 57909 9057 58351 9134
rect 57909 9005 57998 9057
rect 58050 9005 58210 9057
rect 58262 9005 58351 9057
rect 57909 8972 58351 9005
rect 57909 8916 57996 8972
rect 58052 8916 58208 8972
rect 58264 8916 58351 8972
rect 57909 8840 58351 8916
rect 57909 8788 57998 8840
rect 58050 8788 58210 8840
rect 58262 8788 58351 8840
rect 57909 8754 58351 8788
rect 57909 8698 57996 8754
rect 58052 8698 58208 8754
rect 58264 8698 58351 8754
rect 57909 8622 58351 8698
rect 57909 8570 57998 8622
rect 58050 8570 58210 8622
rect 58262 8570 58351 8622
rect 57909 8536 58351 8570
rect 57909 8480 57996 8536
rect 58052 8480 58208 8536
rect 58264 8480 58351 8536
rect 57909 8404 58351 8480
rect 57909 8352 57998 8404
rect 58050 8352 58210 8404
rect 58262 8352 58351 8404
rect 57909 8319 58351 8352
rect 57909 8263 57996 8319
rect 58052 8263 58208 8319
rect 58264 8263 58351 8319
rect 57909 8187 58351 8263
rect 57909 8135 57998 8187
rect 58050 8135 58210 8187
rect 58262 8135 58351 8187
rect 57909 7969 58351 8135
rect 57909 7917 57998 7969
rect 58050 7917 58210 7969
rect 58262 7917 58351 7969
rect 57909 7752 58351 7917
rect 57909 7700 57998 7752
rect 58050 7700 58210 7752
rect 58262 7700 58351 7752
rect 57909 7534 58351 7700
rect 57909 7482 57998 7534
rect 58050 7482 58210 7534
rect 58262 7482 58351 7534
rect 57909 7316 58351 7482
rect 57909 7264 57998 7316
rect 58050 7264 58210 7316
rect 58262 7264 58351 7316
rect 57909 7099 58351 7264
rect 57909 7047 57998 7099
rect 58050 7047 58210 7099
rect 58262 7047 58351 7099
rect 57909 6881 58351 7047
rect 57909 6829 57998 6881
rect 58050 6829 58210 6881
rect 58262 6829 58351 6881
rect 57909 6663 58351 6829
rect 57909 6611 57998 6663
rect 58050 6611 58210 6663
rect 58262 6611 58351 6663
rect 57909 6446 58351 6611
rect 57909 6394 57998 6446
rect 58050 6394 58210 6446
rect 58262 6394 58351 6446
rect 57909 6228 58351 6394
rect 57909 6176 57998 6228
rect 58050 6176 58210 6228
rect 58262 6176 58351 6228
rect 57909 6011 58351 6176
rect 57909 5959 57998 6011
rect 58050 5959 58210 6011
rect 58262 5959 58351 6011
rect 57909 5793 58351 5959
rect 57909 5741 57998 5793
rect 58050 5741 58210 5793
rect 58262 5741 58351 5793
rect 57909 5575 58351 5741
rect 57909 5539 57998 5575
rect 58050 5539 58210 5575
rect 58262 5539 58351 5575
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 58351 5539
rect 57909 5358 58351 5483
rect 57909 5321 57998 5358
rect 58050 5321 58210 5358
rect 58262 5321 58351 5358
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 58351 5321
rect 61277 5479 61457 5491
rect 61277 5462 61289 5479
rect 61445 5462 61457 5479
rect 61277 5302 61287 5462
rect 61447 5302 61457 5462
rect 61277 5292 61457 5302
rect 57909 4587 58351 5265
rect 57909 4535 57998 4587
rect 58050 4535 58210 4587
rect 58262 4535 58351 4587
rect 57909 4528 58351 4535
rect 57909 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4472 58351 4528
rect 57909 4370 58351 4472
rect 57909 4318 57998 4370
rect 58050 4318 58210 4370
rect 58262 4318 58351 4370
rect 57909 4310 58351 4318
rect 57909 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 58351 4310
rect 57909 4152 58351 4254
rect 57909 4100 57998 4152
rect 58050 4100 58210 4152
rect 58262 4100 58351 4152
rect 57909 3934 58351 4100
rect 57909 3882 57998 3934
rect 58050 3882 58210 3934
rect 58262 3882 58351 3934
rect 57909 3717 58351 3882
rect 57909 3665 57998 3717
rect 58050 3665 58210 3717
rect 58262 3665 58351 3717
rect 57909 3524 58351 3665
rect 61507 5024 62085 5135
rect 71303 5073 71359 5140
rect 53772 3096 55669 3309
rect 53772 0 53996 3096
rect 55781 2836 55911 3418
rect 54417 2623 55911 2836
rect 54417 0 54641 2623
rect 56023 2416 56153 3420
rect 55164 2203 56153 2416
rect 56265 2907 56394 3418
rect 55164 0 55388 2203
rect 56265 0 56489 2907
rect 61507 1701 61601 5024
rect 62839 5001 62933 5062
rect 71193 5017 71359 5073
rect 62839 4880 63115 5001
rect 63021 1701 63115 4880
rect 71193 1701 71249 5017
rect 72151 4740 72207 5185
rect 71866 4684 72207 4740
rect 72829 4740 72885 5185
rect 73677 5073 73733 5140
rect 82103 5073 82159 5140
rect 73677 5017 73843 5073
rect 72829 4684 73170 4740
rect 71866 1701 71922 4684
rect 73114 1701 73170 4684
rect 73787 1701 73843 5017
rect 81939 5017 82159 5073
rect 81939 1701 81995 5017
rect 82970 4740 83026 5185
rect 82970 4684 83512 4740
rect 83456 1701 83512 4684
rect 61447 0 61671 1701
rect 62115 1689 62339 1701
rect 62115 1637 62149 1689
rect 62305 1637 62339 1689
rect 62115 0 62339 1637
rect 62958 0 63182 1701
rect 71109 0 71333 1701
rect 71782 0 72006 1701
rect 72180 1689 72404 1701
rect 72180 1637 72215 1689
rect 72371 1637 72404 1689
rect 72180 0 72404 1637
rect 72630 1689 72854 1701
rect 72630 1637 72665 1689
rect 72821 1637 72854 1689
rect 72630 0 72854 1637
rect 73030 0 73254 1701
rect 73703 0 73927 1701
rect 81855 0 82079 1701
rect 82695 1689 82919 1701
rect 82695 1637 82730 1689
rect 82886 1637 82919 1689
rect 82695 0 82919 1637
rect 83372 0 83596 1701
<< via2 >>
rect 25378 65914 25434 65916
rect 25378 65862 25380 65914
rect 25380 65862 25432 65914
rect 25432 65862 25434 65914
rect 25378 65860 25434 65862
rect 25502 65914 25558 65916
rect 25502 65862 25504 65914
rect 25504 65862 25556 65914
rect 25556 65862 25558 65914
rect 25502 65860 25558 65862
rect 25626 65914 25682 65916
rect 25626 65862 25628 65914
rect 25628 65862 25680 65914
rect 25680 65862 25682 65914
rect 25626 65860 25682 65862
rect 25750 65914 25806 65916
rect 25750 65862 25752 65914
rect 25752 65862 25804 65914
rect 25804 65862 25806 65914
rect 25750 65860 25806 65862
rect 25874 65914 25930 65916
rect 25874 65862 25876 65914
rect 25876 65862 25928 65914
rect 25928 65862 25930 65914
rect 25874 65860 25930 65862
rect 25378 65790 25434 65792
rect 25378 65738 25380 65790
rect 25380 65738 25432 65790
rect 25432 65738 25434 65790
rect 25378 65736 25434 65738
rect 25502 65790 25558 65792
rect 25502 65738 25504 65790
rect 25504 65738 25556 65790
rect 25556 65738 25558 65790
rect 25502 65736 25558 65738
rect 25626 65790 25682 65792
rect 25626 65738 25628 65790
rect 25628 65738 25680 65790
rect 25680 65738 25682 65790
rect 25626 65736 25682 65738
rect 25750 65790 25806 65792
rect 25750 65738 25752 65790
rect 25752 65738 25804 65790
rect 25804 65738 25806 65790
rect 25750 65736 25806 65738
rect 25874 65790 25930 65792
rect 25874 65738 25876 65790
rect 25876 65738 25928 65790
rect 25928 65738 25930 65790
rect 25874 65736 25930 65738
rect 25344 34959 25400 34961
rect 25344 34907 25346 34959
rect 25346 34907 25398 34959
rect 25398 34907 25400 34959
rect 25344 34905 25400 34907
rect 25468 34959 25524 34961
rect 25468 34907 25470 34959
rect 25470 34907 25522 34959
rect 25522 34907 25524 34959
rect 25468 34905 25524 34907
rect 25592 34959 25648 34961
rect 25592 34907 25594 34959
rect 25594 34907 25646 34959
rect 25646 34907 25648 34959
rect 25592 34905 25648 34907
rect 25716 34959 25772 34961
rect 25716 34907 25718 34959
rect 25718 34907 25770 34959
rect 25770 34907 25772 34959
rect 25716 34905 25772 34907
rect 25840 34959 25896 34961
rect 25840 34907 25842 34959
rect 25842 34907 25894 34959
rect 25894 34907 25896 34959
rect 25840 34905 25896 34907
rect 25964 34959 26020 34961
rect 25964 34907 25966 34959
rect 25966 34907 26018 34959
rect 26018 34907 26020 34959
rect 25964 34905 26020 34907
rect 25344 34835 25400 34837
rect 25344 34783 25346 34835
rect 25346 34783 25398 34835
rect 25398 34783 25400 34835
rect 25344 34781 25400 34783
rect 25468 34835 25524 34837
rect 25468 34783 25470 34835
rect 25470 34783 25522 34835
rect 25522 34783 25524 34835
rect 25468 34781 25524 34783
rect 25592 34835 25648 34837
rect 25592 34783 25594 34835
rect 25594 34783 25646 34835
rect 25646 34783 25648 34835
rect 25592 34781 25648 34783
rect 25716 34835 25772 34837
rect 25716 34783 25718 34835
rect 25718 34783 25770 34835
rect 25770 34783 25772 34835
rect 25716 34781 25772 34783
rect 25840 34835 25896 34837
rect 25840 34783 25842 34835
rect 25842 34783 25894 34835
rect 25894 34783 25896 34835
rect 25840 34781 25896 34783
rect 25964 34835 26020 34837
rect 25964 34783 25966 34835
rect 25966 34783 26018 34835
rect 26018 34783 26020 34835
rect 25964 34781 26020 34783
rect 25344 34711 25400 34713
rect 25344 34659 25346 34711
rect 25346 34659 25398 34711
rect 25398 34659 25400 34711
rect 25344 34657 25400 34659
rect 25468 34711 25524 34713
rect 25468 34659 25470 34711
rect 25470 34659 25522 34711
rect 25522 34659 25524 34711
rect 25468 34657 25524 34659
rect 25592 34711 25648 34713
rect 25592 34659 25594 34711
rect 25594 34659 25646 34711
rect 25646 34659 25648 34711
rect 25592 34657 25648 34659
rect 25716 34711 25772 34713
rect 25716 34659 25718 34711
rect 25718 34659 25770 34711
rect 25770 34659 25772 34711
rect 25716 34657 25772 34659
rect 25840 34711 25896 34713
rect 25840 34659 25842 34711
rect 25842 34659 25894 34711
rect 25894 34659 25896 34711
rect 25840 34657 25896 34659
rect 25964 34711 26020 34713
rect 25964 34659 25966 34711
rect 25966 34659 26018 34711
rect 26018 34659 26020 34711
rect 25964 34657 26020 34659
rect 25398 31192 25454 31248
rect 25522 31192 25578 31248
rect 25646 31192 25702 31248
rect 25770 31192 25826 31248
rect 25894 31192 25950 31248
rect 25398 31068 25454 31124
rect 25522 31068 25578 31124
rect 25646 31068 25702 31124
rect 25770 31068 25826 31124
rect 25894 31068 25950 31124
rect 25398 30944 25454 31000
rect 25522 30944 25578 31000
rect 25646 30944 25702 31000
rect 25770 30944 25826 31000
rect 25894 30944 25950 31000
rect 25398 30737 25454 30793
rect 25522 30737 25578 30793
rect 25646 30737 25702 30793
rect 25770 30737 25826 30793
rect 25894 30737 25950 30793
rect 25398 30613 25454 30669
rect 25522 30613 25578 30669
rect 25646 30613 25702 30669
rect 25770 30613 25826 30669
rect 25894 30613 25950 30669
rect 25398 30489 25454 30545
rect 25522 30489 25578 30545
rect 25646 30489 25702 30545
rect 25770 30489 25826 30545
rect 25894 30489 25950 30545
rect 25404 28259 25460 28315
rect 25528 28259 25584 28315
rect 25652 28259 25708 28315
rect 25776 28259 25832 28315
rect 25900 28259 25956 28315
rect 25404 28135 25460 28191
rect 25528 28135 25584 28191
rect 25652 28135 25708 28191
rect 25776 28135 25832 28191
rect 25900 28135 25956 28191
rect 25404 28011 25460 28067
rect 25528 28011 25584 28067
rect 25652 28011 25708 28067
rect 25776 28011 25832 28067
rect 25900 28011 25956 28067
rect 25404 27887 25460 27943
rect 25528 27887 25584 27943
rect 25652 27887 25708 27943
rect 25776 27887 25832 27943
rect 25900 27887 25956 27943
rect 25404 27763 25460 27819
rect 25528 27763 25584 27819
rect 25652 27763 25708 27819
rect 25776 27763 25832 27819
rect 25900 27763 25956 27819
rect 25404 27639 25460 27695
rect 25528 27639 25584 27695
rect 25652 27639 25708 27695
rect 25776 27639 25832 27695
rect 25900 27639 25956 27695
rect 25404 27515 25460 27571
rect 25528 27515 25584 27571
rect 25652 27515 25708 27571
rect 25776 27515 25832 27571
rect 25900 27515 25956 27571
rect 25404 27391 25460 27447
rect 25528 27391 25584 27447
rect 25652 27391 25708 27447
rect 25776 27391 25832 27447
rect 25900 27391 25956 27447
rect 26859 33955 26915 34011
rect 27071 33955 27127 34011
rect 26859 33737 26915 33793
rect 27071 33737 27127 33793
rect 26859 33520 26915 33576
rect 27071 33520 27127 33576
rect 26859 33302 26915 33358
rect 27071 33302 27127 33358
rect 26859 33084 26915 33140
rect 27071 33084 27127 33140
rect 26859 32866 26915 32922
rect 27071 32866 27127 32922
rect 26859 32649 26915 32705
rect 27071 32649 27127 32705
rect 26859 32431 26915 32487
rect 27071 32431 27127 32487
rect 26859 32075 26861 32088
rect 26861 32075 26913 32088
rect 26913 32075 26915 32088
rect 26859 32032 26915 32075
rect 27071 32075 27073 32088
rect 27073 32075 27125 32088
rect 27125 32075 27127 32088
rect 27071 32032 27127 32075
rect 26859 31857 26861 31870
rect 26861 31857 26913 31870
rect 26913 31857 26915 31870
rect 26859 31814 26915 31857
rect 27071 31857 27073 31870
rect 27073 31857 27125 31870
rect 27125 31857 27127 31870
rect 27071 31814 27127 31857
rect 26859 31639 26861 31652
rect 26861 31639 26913 31652
rect 26913 31639 26915 31652
rect 26859 31596 26915 31639
rect 27071 31639 27073 31652
rect 27073 31639 27125 31652
rect 27125 31639 27127 31652
rect 27071 31596 27127 31639
rect 26859 29950 26915 29968
rect 26859 29912 26861 29950
rect 26861 29912 26913 29950
rect 26913 29912 26915 29950
rect 27071 29950 27127 29968
rect 27071 29912 27073 29950
rect 27073 29912 27125 29950
rect 27125 29912 27127 29950
rect 26859 29733 26915 29750
rect 26859 29694 26861 29733
rect 26861 29694 26913 29733
rect 26913 29694 26915 29733
rect 27071 29733 27127 29750
rect 27071 29694 27073 29733
rect 27073 29694 27125 29733
rect 27125 29694 27127 29733
rect 26859 29515 26915 29533
rect 26859 29477 26861 29515
rect 26861 29477 26913 29515
rect 26913 29477 26915 29515
rect 27071 29515 27127 29533
rect 27071 29477 27073 29515
rect 27073 29477 27125 29515
rect 27125 29477 27127 29515
rect 26859 29297 26915 29315
rect 26859 29259 26861 29297
rect 26861 29259 26913 29297
rect 26913 29259 26915 29297
rect 27071 29297 27127 29315
rect 27071 29259 27073 29297
rect 27073 29259 27125 29297
rect 27125 29259 27127 29297
rect 26859 29080 26915 29098
rect 26859 29042 26861 29080
rect 26861 29042 26913 29080
rect 26913 29042 26915 29080
rect 27071 29080 27127 29098
rect 27071 29042 27073 29080
rect 27073 29042 27125 29080
rect 27125 29042 27127 29080
rect 26859 28862 26915 28880
rect 26859 28824 26861 28862
rect 26861 28824 26913 28862
rect 26913 28824 26915 28862
rect 27071 28862 27127 28880
rect 27071 28824 27073 28862
rect 27073 28824 27125 28862
rect 27125 28824 27127 28862
rect 26859 28644 26915 28662
rect 26859 28606 26861 28644
rect 26861 28606 26913 28644
rect 26913 28606 26915 28644
rect 27071 28644 27127 28662
rect 27071 28606 27073 28644
rect 27073 28606 27125 28644
rect 27125 28606 27127 28644
rect 26859 28427 26915 28444
rect 26859 28388 26861 28427
rect 26861 28388 26913 28427
rect 26913 28388 26915 28427
rect 27071 28427 27127 28444
rect 27071 28388 27073 28427
rect 27073 28388 27125 28427
rect 27125 28388 27127 28427
rect 26859 28209 26915 28227
rect 26859 28171 26861 28209
rect 26861 28171 26913 28209
rect 26913 28171 26915 28209
rect 27071 28209 27127 28227
rect 27071 28171 27073 28209
rect 27073 28171 27125 28209
rect 27125 28171 27127 28209
rect 26859 27992 26915 28009
rect 26859 27953 26861 27992
rect 26861 27953 26913 27992
rect 26913 27953 26915 27992
rect 27071 27992 27127 28009
rect 27071 27953 27073 27992
rect 27073 27953 27125 27992
rect 27125 27953 27127 27992
rect 26859 27774 26915 27792
rect 26859 27736 26861 27774
rect 26861 27736 26913 27774
rect 26913 27736 26915 27774
rect 27071 27774 27127 27792
rect 27071 27736 27073 27774
rect 27073 27736 27125 27774
rect 27125 27736 27127 27774
rect 26859 27556 26915 27574
rect 26859 27518 26861 27556
rect 26861 27518 26913 27556
rect 26913 27518 26915 27556
rect 27071 27556 27127 27574
rect 27071 27518 27073 27556
rect 27073 27518 27125 27556
rect 27125 27518 27127 27556
rect 27788 65853 27844 65855
rect 27788 65801 27790 65853
rect 27790 65801 27842 65853
rect 27842 65801 27844 65853
rect 27788 65799 27844 65801
rect 27999 65853 28055 65855
rect 27999 65801 28001 65853
rect 28001 65801 28053 65853
rect 28053 65801 28055 65853
rect 27999 65799 28055 65801
rect 28210 65853 28266 65855
rect 28210 65801 28212 65853
rect 28212 65801 28264 65853
rect 28264 65801 28266 65853
rect 28210 65799 28266 65801
rect 28421 65853 28477 65855
rect 28421 65801 28423 65853
rect 28423 65801 28475 65853
rect 28475 65801 28477 65853
rect 28421 65799 28477 65801
rect 28632 65853 28688 65855
rect 28632 65801 28634 65853
rect 28634 65801 28686 65853
rect 28686 65801 28688 65853
rect 28632 65799 28688 65801
rect 28843 65853 28899 65855
rect 28843 65801 28845 65853
rect 28845 65801 28897 65853
rect 28897 65801 28899 65853
rect 28843 65799 28899 65801
rect 29054 65853 29110 65855
rect 29054 65801 29056 65853
rect 29056 65801 29108 65853
rect 29108 65801 29110 65853
rect 29054 65799 29110 65801
rect 29580 64953 29636 64955
rect 29580 64901 29582 64953
rect 29582 64901 29634 64953
rect 29634 64901 29636 64953
rect 29580 64899 29636 64901
rect 29791 64953 29847 64955
rect 29791 64901 29793 64953
rect 29793 64901 29845 64953
rect 29845 64901 29847 64953
rect 29791 64899 29847 64901
rect 30003 64953 30059 64955
rect 30003 64901 30005 64953
rect 30005 64901 30057 64953
rect 30057 64901 30059 64953
rect 30003 64899 30059 64901
rect 30214 64953 30270 64955
rect 30214 64901 30216 64953
rect 30216 64901 30268 64953
rect 30268 64901 30270 64953
rect 30214 64899 30270 64901
rect 34288 65853 34344 65855
rect 34288 65801 34290 65853
rect 34290 65801 34342 65853
rect 34342 65801 34344 65853
rect 34288 65799 34344 65801
rect 34499 65853 34555 65855
rect 34499 65801 34501 65853
rect 34501 65801 34553 65853
rect 34553 65801 34555 65853
rect 34499 65799 34555 65801
rect 34710 65853 34766 65855
rect 34710 65801 34712 65853
rect 34712 65801 34764 65853
rect 34764 65801 34766 65853
rect 34710 65799 34766 65801
rect 34921 65853 34977 65855
rect 34921 65801 34923 65853
rect 34923 65801 34975 65853
rect 34975 65801 34977 65853
rect 34921 65799 34977 65801
rect 33048 65372 33104 65374
rect 33048 65320 33050 65372
rect 33050 65320 33102 65372
rect 33102 65320 33104 65372
rect 33048 65318 33104 65320
rect 33259 65372 33315 65374
rect 33259 65320 33261 65372
rect 33261 65320 33313 65372
rect 33313 65320 33315 65372
rect 33259 65318 33315 65320
rect 33470 65372 33526 65374
rect 33470 65320 33472 65372
rect 33472 65320 33524 65372
rect 33524 65320 33526 65372
rect 33470 65318 33526 65320
rect 33681 65372 33737 65374
rect 33681 65320 33683 65372
rect 33683 65320 33735 65372
rect 33735 65320 33737 65372
rect 33681 65318 33737 65320
rect 33892 65372 33948 65374
rect 33892 65320 33894 65372
rect 33894 65320 33946 65372
rect 33946 65320 33948 65372
rect 33892 65318 33948 65320
rect 30852 64953 30908 64955
rect 27788 64053 27844 64055
rect 27788 64001 27790 64053
rect 27790 64001 27842 64053
rect 27842 64001 27844 64053
rect 27788 63999 27844 64001
rect 27999 64053 28055 64055
rect 27999 64001 28001 64053
rect 28001 64001 28053 64053
rect 28053 64001 28055 64053
rect 27999 63999 28055 64001
rect 28210 64053 28266 64055
rect 28210 64001 28212 64053
rect 28212 64001 28264 64053
rect 28264 64001 28266 64053
rect 28210 63999 28266 64001
rect 28421 64053 28477 64055
rect 28421 64001 28423 64053
rect 28423 64001 28475 64053
rect 28475 64001 28477 64053
rect 28421 63999 28477 64001
rect 28632 64053 28688 64055
rect 28632 64001 28634 64053
rect 28634 64001 28686 64053
rect 28686 64001 28688 64053
rect 28632 63999 28688 64001
rect 28843 64053 28899 64055
rect 28843 64001 28845 64053
rect 28845 64001 28897 64053
rect 28897 64001 28899 64053
rect 28843 63999 28899 64001
rect 29054 64053 29110 64055
rect 29054 64001 29056 64053
rect 29056 64001 29108 64053
rect 29108 64001 29110 64053
rect 29054 63999 29110 64001
rect 29580 63153 29636 63155
rect 29580 63101 29582 63153
rect 29582 63101 29634 63153
rect 29634 63101 29636 63153
rect 29580 63099 29636 63101
rect 29791 63153 29847 63155
rect 29791 63101 29793 63153
rect 29793 63101 29845 63153
rect 29845 63101 29847 63153
rect 29791 63099 29847 63101
rect 30003 63153 30059 63155
rect 30003 63101 30005 63153
rect 30005 63101 30057 63153
rect 30057 63101 30059 63153
rect 30003 63099 30059 63101
rect 30214 63153 30270 63155
rect 30214 63101 30216 63153
rect 30216 63101 30268 63153
rect 30268 63101 30270 63153
rect 30214 63099 30270 63101
rect 27788 62253 27844 62255
rect 27788 62201 27790 62253
rect 27790 62201 27842 62253
rect 27842 62201 27844 62253
rect 27788 62199 27844 62201
rect 27999 62253 28055 62255
rect 27999 62201 28001 62253
rect 28001 62201 28053 62253
rect 28053 62201 28055 62253
rect 27999 62199 28055 62201
rect 28210 62253 28266 62255
rect 28210 62201 28212 62253
rect 28212 62201 28264 62253
rect 28264 62201 28266 62253
rect 28210 62199 28266 62201
rect 28421 62253 28477 62255
rect 28421 62201 28423 62253
rect 28423 62201 28475 62253
rect 28475 62201 28477 62253
rect 28421 62199 28477 62201
rect 28632 62253 28688 62255
rect 28632 62201 28634 62253
rect 28634 62201 28686 62253
rect 28686 62201 28688 62253
rect 28632 62199 28688 62201
rect 28843 62253 28899 62255
rect 28843 62201 28845 62253
rect 28845 62201 28897 62253
rect 28897 62201 28899 62253
rect 28843 62199 28899 62201
rect 29054 62253 29110 62255
rect 29054 62201 29056 62253
rect 29056 62201 29108 62253
rect 29108 62201 29110 62253
rect 29054 62199 29110 62201
rect 29580 61353 29636 61355
rect 29580 61301 29582 61353
rect 29582 61301 29634 61353
rect 29634 61301 29636 61353
rect 29580 61299 29636 61301
rect 29791 61353 29847 61355
rect 29791 61301 29793 61353
rect 29793 61301 29845 61353
rect 29845 61301 29847 61353
rect 29791 61299 29847 61301
rect 30003 61353 30059 61355
rect 30003 61301 30005 61353
rect 30005 61301 30057 61353
rect 30057 61301 30059 61353
rect 30003 61299 30059 61301
rect 30214 61353 30270 61355
rect 30214 61301 30216 61353
rect 30216 61301 30268 61353
rect 30268 61301 30270 61353
rect 30214 61299 30270 61301
rect 27788 60453 27844 60455
rect 27788 60401 27790 60453
rect 27790 60401 27842 60453
rect 27842 60401 27844 60453
rect 27788 60399 27844 60401
rect 27999 60453 28055 60455
rect 27999 60401 28001 60453
rect 28001 60401 28053 60453
rect 28053 60401 28055 60453
rect 27999 60399 28055 60401
rect 28210 60453 28266 60455
rect 28210 60401 28212 60453
rect 28212 60401 28264 60453
rect 28264 60401 28266 60453
rect 28210 60399 28266 60401
rect 28421 60453 28477 60455
rect 28421 60401 28423 60453
rect 28423 60401 28475 60453
rect 28475 60401 28477 60453
rect 28421 60399 28477 60401
rect 28632 60453 28688 60455
rect 28632 60401 28634 60453
rect 28634 60401 28686 60453
rect 28686 60401 28688 60453
rect 28632 60399 28688 60401
rect 28843 60453 28899 60455
rect 28843 60401 28845 60453
rect 28845 60401 28897 60453
rect 28897 60401 28899 60453
rect 28843 60399 28899 60401
rect 29054 60453 29110 60455
rect 29054 60401 29056 60453
rect 29056 60401 29108 60453
rect 29108 60401 29110 60453
rect 29054 60399 29110 60401
rect 29580 59553 29636 59555
rect 29580 59501 29582 59553
rect 29582 59501 29634 59553
rect 29634 59501 29636 59553
rect 29580 59499 29636 59501
rect 29791 59553 29847 59555
rect 29791 59501 29793 59553
rect 29793 59501 29845 59553
rect 29845 59501 29847 59553
rect 29791 59499 29847 59501
rect 30003 59553 30059 59555
rect 30003 59501 30005 59553
rect 30005 59501 30057 59553
rect 30057 59501 30059 59553
rect 30003 59499 30059 59501
rect 30214 59553 30270 59555
rect 30214 59501 30216 59553
rect 30216 59501 30268 59553
rect 30268 59501 30270 59553
rect 30214 59499 30270 59501
rect 27788 58653 27844 58655
rect 27788 58601 27790 58653
rect 27790 58601 27842 58653
rect 27842 58601 27844 58653
rect 27788 58599 27844 58601
rect 27999 58653 28055 58655
rect 27999 58601 28001 58653
rect 28001 58601 28053 58653
rect 28053 58601 28055 58653
rect 27999 58599 28055 58601
rect 28210 58653 28266 58655
rect 28210 58601 28212 58653
rect 28212 58601 28264 58653
rect 28264 58601 28266 58653
rect 28210 58599 28266 58601
rect 28421 58653 28477 58655
rect 28421 58601 28423 58653
rect 28423 58601 28475 58653
rect 28475 58601 28477 58653
rect 28421 58599 28477 58601
rect 28632 58653 28688 58655
rect 28632 58601 28634 58653
rect 28634 58601 28686 58653
rect 28686 58601 28688 58653
rect 28632 58599 28688 58601
rect 28843 58653 28899 58655
rect 28843 58601 28845 58653
rect 28845 58601 28897 58653
rect 28897 58601 28899 58653
rect 28843 58599 28899 58601
rect 29054 58653 29110 58655
rect 29054 58601 29056 58653
rect 29056 58601 29108 58653
rect 29108 58601 29110 58653
rect 29054 58599 29110 58601
rect 29580 57753 29636 57755
rect 29580 57701 29582 57753
rect 29582 57701 29634 57753
rect 29634 57701 29636 57753
rect 29580 57699 29636 57701
rect 29791 57753 29847 57755
rect 29791 57701 29793 57753
rect 29793 57701 29845 57753
rect 29845 57701 29847 57753
rect 29791 57699 29847 57701
rect 30003 57753 30059 57755
rect 30003 57701 30005 57753
rect 30005 57701 30057 57753
rect 30057 57701 30059 57753
rect 30003 57699 30059 57701
rect 30214 57753 30270 57755
rect 30214 57701 30216 57753
rect 30216 57701 30268 57753
rect 30268 57701 30270 57753
rect 30214 57699 30270 57701
rect 27788 56853 27844 56855
rect 27788 56801 27790 56853
rect 27790 56801 27842 56853
rect 27842 56801 27844 56853
rect 27788 56799 27844 56801
rect 27999 56853 28055 56855
rect 27999 56801 28001 56853
rect 28001 56801 28053 56853
rect 28053 56801 28055 56853
rect 27999 56799 28055 56801
rect 28210 56853 28266 56855
rect 28210 56801 28212 56853
rect 28212 56801 28264 56853
rect 28264 56801 28266 56853
rect 28210 56799 28266 56801
rect 28421 56853 28477 56855
rect 28421 56801 28423 56853
rect 28423 56801 28475 56853
rect 28475 56801 28477 56853
rect 28421 56799 28477 56801
rect 28632 56853 28688 56855
rect 28632 56801 28634 56853
rect 28634 56801 28686 56853
rect 28686 56801 28688 56853
rect 28632 56799 28688 56801
rect 28843 56853 28899 56855
rect 28843 56801 28845 56853
rect 28845 56801 28897 56853
rect 28897 56801 28899 56853
rect 28843 56799 28899 56801
rect 29054 56853 29110 56855
rect 29054 56801 29056 56853
rect 29056 56801 29108 56853
rect 29108 56801 29110 56853
rect 29054 56799 29110 56801
rect 29580 55953 29636 55955
rect 29580 55901 29582 55953
rect 29582 55901 29634 55953
rect 29634 55901 29636 55953
rect 29580 55899 29636 55901
rect 29791 55953 29847 55955
rect 29791 55901 29793 55953
rect 29793 55901 29845 55953
rect 29845 55901 29847 55953
rect 29791 55899 29847 55901
rect 30003 55953 30059 55955
rect 30003 55901 30005 55953
rect 30005 55901 30057 55953
rect 30057 55901 30059 55953
rect 30003 55899 30059 55901
rect 30214 55953 30270 55955
rect 30214 55901 30216 55953
rect 30216 55901 30268 55953
rect 30268 55901 30270 55953
rect 30214 55899 30270 55901
rect 27788 55053 27844 55055
rect 27788 55001 27790 55053
rect 27790 55001 27842 55053
rect 27842 55001 27844 55053
rect 27788 54999 27844 55001
rect 27999 55053 28055 55055
rect 27999 55001 28001 55053
rect 28001 55001 28053 55053
rect 28053 55001 28055 55053
rect 27999 54999 28055 55001
rect 28210 55053 28266 55055
rect 28210 55001 28212 55053
rect 28212 55001 28264 55053
rect 28264 55001 28266 55053
rect 28210 54999 28266 55001
rect 28421 55053 28477 55055
rect 28421 55001 28423 55053
rect 28423 55001 28475 55053
rect 28475 55001 28477 55053
rect 28421 54999 28477 55001
rect 28632 55053 28688 55055
rect 28632 55001 28634 55053
rect 28634 55001 28686 55053
rect 28686 55001 28688 55053
rect 28632 54999 28688 55001
rect 28843 55053 28899 55055
rect 28843 55001 28845 55053
rect 28845 55001 28897 55053
rect 28897 55001 28899 55053
rect 28843 54999 28899 55001
rect 29054 55053 29110 55055
rect 29054 55001 29056 55053
rect 29056 55001 29108 55053
rect 29108 55001 29110 55053
rect 29054 54999 29110 55001
rect 29580 54153 29636 54155
rect 29580 54101 29582 54153
rect 29582 54101 29634 54153
rect 29634 54101 29636 54153
rect 29580 54099 29636 54101
rect 29791 54153 29847 54155
rect 29791 54101 29793 54153
rect 29793 54101 29845 54153
rect 29845 54101 29847 54153
rect 29791 54099 29847 54101
rect 30003 54153 30059 54155
rect 30003 54101 30005 54153
rect 30005 54101 30057 54153
rect 30057 54101 30059 54153
rect 30003 54099 30059 54101
rect 30214 54153 30270 54155
rect 30214 54101 30216 54153
rect 30216 54101 30268 54153
rect 30268 54101 30270 54153
rect 30214 54099 30270 54101
rect 27788 53253 27844 53255
rect 27788 53201 27790 53253
rect 27790 53201 27842 53253
rect 27842 53201 27844 53253
rect 27788 53199 27844 53201
rect 27999 53253 28055 53255
rect 27999 53201 28001 53253
rect 28001 53201 28053 53253
rect 28053 53201 28055 53253
rect 27999 53199 28055 53201
rect 28210 53253 28266 53255
rect 28210 53201 28212 53253
rect 28212 53201 28264 53253
rect 28264 53201 28266 53253
rect 28210 53199 28266 53201
rect 28421 53253 28477 53255
rect 28421 53201 28423 53253
rect 28423 53201 28475 53253
rect 28475 53201 28477 53253
rect 28421 53199 28477 53201
rect 28632 53253 28688 53255
rect 28632 53201 28634 53253
rect 28634 53201 28686 53253
rect 28686 53201 28688 53253
rect 28632 53199 28688 53201
rect 28843 53253 28899 53255
rect 28843 53201 28845 53253
rect 28845 53201 28897 53253
rect 28897 53201 28899 53253
rect 28843 53199 28899 53201
rect 29054 53253 29110 53255
rect 29054 53201 29056 53253
rect 29056 53201 29108 53253
rect 29108 53201 29110 53253
rect 29054 53199 29110 53201
rect 29580 52353 29636 52355
rect 29580 52301 29582 52353
rect 29582 52301 29634 52353
rect 29634 52301 29636 52353
rect 29580 52299 29636 52301
rect 29791 52353 29847 52355
rect 29791 52301 29793 52353
rect 29793 52301 29845 52353
rect 29845 52301 29847 52353
rect 29791 52299 29847 52301
rect 30003 52353 30059 52355
rect 30003 52301 30005 52353
rect 30005 52301 30057 52353
rect 30057 52301 30059 52353
rect 30003 52299 30059 52301
rect 30214 52353 30270 52355
rect 30214 52301 30216 52353
rect 30216 52301 30268 52353
rect 30268 52301 30270 52353
rect 30214 52299 30270 52301
rect 27788 51453 27844 51455
rect 27788 51401 27790 51453
rect 27790 51401 27842 51453
rect 27842 51401 27844 51453
rect 27788 51399 27844 51401
rect 27999 51453 28055 51455
rect 27999 51401 28001 51453
rect 28001 51401 28053 51453
rect 28053 51401 28055 51453
rect 27999 51399 28055 51401
rect 28210 51453 28266 51455
rect 28210 51401 28212 51453
rect 28212 51401 28264 51453
rect 28264 51401 28266 51453
rect 28210 51399 28266 51401
rect 28421 51453 28477 51455
rect 28421 51401 28423 51453
rect 28423 51401 28475 51453
rect 28475 51401 28477 51453
rect 28421 51399 28477 51401
rect 28632 51453 28688 51455
rect 28632 51401 28634 51453
rect 28634 51401 28686 51453
rect 28686 51401 28688 51453
rect 28632 51399 28688 51401
rect 28843 51453 28899 51455
rect 28843 51401 28845 51453
rect 28845 51401 28897 51453
rect 28897 51401 28899 51453
rect 28843 51399 28899 51401
rect 29054 51453 29110 51455
rect 29054 51401 29056 51453
rect 29056 51401 29108 51453
rect 29108 51401 29110 51453
rect 29054 51399 29110 51401
rect 29580 50553 29636 50555
rect 29580 50501 29582 50553
rect 29582 50501 29634 50553
rect 29634 50501 29636 50553
rect 29580 50499 29636 50501
rect 29791 50553 29847 50555
rect 29791 50501 29793 50553
rect 29793 50501 29845 50553
rect 29845 50501 29847 50553
rect 29791 50499 29847 50501
rect 30003 50553 30059 50555
rect 30003 50501 30005 50553
rect 30005 50501 30057 50553
rect 30057 50501 30059 50553
rect 30003 50499 30059 50501
rect 30214 50553 30270 50555
rect 30214 50501 30216 50553
rect 30216 50501 30268 50553
rect 30268 50501 30270 50553
rect 30214 50499 30270 50501
rect 27788 49653 27844 49655
rect 27788 49601 27790 49653
rect 27790 49601 27842 49653
rect 27842 49601 27844 49653
rect 27788 49599 27844 49601
rect 27999 49653 28055 49655
rect 27999 49601 28001 49653
rect 28001 49601 28053 49653
rect 28053 49601 28055 49653
rect 27999 49599 28055 49601
rect 28210 49653 28266 49655
rect 28210 49601 28212 49653
rect 28212 49601 28264 49653
rect 28264 49601 28266 49653
rect 28210 49599 28266 49601
rect 28421 49653 28477 49655
rect 28421 49601 28423 49653
rect 28423 49601 28475 49653
rect 28475 49601 28477 49653
rect 28421 49599 28477 49601
rect 28632 49653 28688 49655
rect 28632 49601 28634 49653
rect 28634 49601 28686 49653
rect 28686 49601 28688 49653
rect 28632 49599 28688 49601
rect 28843 49653 28899 49655
rect 28843 49601 28845 49653
rect 28845 49601 28897 49653
rect 28897 49601 28899 49653
rect 28843 49599 28899 49601
rect 29054 49653 29110 49655
rect 29054 49601 29056 49653
rect 29056 49601 29108 49653
rect 29108 49601 29110 49653
rect 29054 49599 29110 49601
rect 29580 48753 29636 48755
rect 29580 48701 29582 48753
rect 29582 48701 29634 48753
rect 29634 48701 29636 48753
rect 29580 48699 29636 48701
rect 29791 48753 29847 48755
rect 29791 48701 29793 48753
rect 29793 48701 29845 48753
rect 29845 48701 29847 48753
rect 29791 48699 29847 48701
rect 30003 48753 30059 48755
rect 30003 48701 30005 48753
rect 30005 48701 30057 48753
rect 30057 48701 30059 48753
rect 30003 48699 30059 48701
rect 30214 48753 30270 48755
rect 30214 48701 30216 48753
rect 30216 48701 30268 48753
rect 30268 48701 30270 48753
rect 30214 48699 30270 48701
rect 27788 47853 27844 47855
rect 27788 47801 27790 47853
rect 27790 47801 27842 47853
rect 27842 47801 27844 47853
rect 27788 47799 27844 47801
rect 27999 47853 28055 47855
rect 27999 47801 28001 47853
rect 28001 47801 28053 47853
rect 28053 47801 28055 47853
rect 27999 47799 28055 47801
rect 28210 47853 28266 47855
rect 28210 47801 28212 47853
rect 28212 47801 28264 47853
rect 28264 47801 28266 47853
rect 28210 47799 28266 47801
rect 28421 47853 28477 47855
rect 28421 47801 28423 47853
rect 28423 47801 28475 47853
rect 28475 47801 28477 47853
rect 28421 47799 28477 47801
rect 28632 47853 28688 47855
rect 28632 47801 28634 47853
rect 28634 47801 28686 47853
rect 28686 47801 28688 47853
rect 28632 47799 28688 47801
rect 28843 47853 28899 47855
rect 28843 47801 28845 47853
rect 28845 47801 28897 47853
rect 28897 47801 28899 47853
rect 28843 47799 28899 47801
rect 29054 47853 29110 47855
rect 29054 47801 29056 47853
rect 29056 47801 29108 47853
rect 29108 47801 29110 47853
rect 29054 47799 29110 47801
rect 29580 46953 29636 46955
rect 29580 46901 29582 46953
rect 29582 46901 29634 46953
rect 29634 46901 29636 46953
rect 29580 46899 29636 46901
rect 29791 46953 29847 46955
rect 29791 46901 29793 46953
rect 29793 46901 29845 46953
rect 29845 46901 29847 46953
rect 29791 46899 29847 46901
rect 30003 46953 30059 46955
rect 30003 46901 30005 46953
rect 30005 46901 30057 46953
rect 30057 46901 30059 46953
rect 30003 46899 30059 46901
rect 30214 46953 30270 46955
rect 30214 46901 30216 46953
rect 30216 46901 30268 46953
rect 30268 46901 30270 46953
rect 30214 46899 30270 46901
rect 27788 46053 27844 46055
rect 27788 46001 27790 46053
rect 27790 46001 27842 46053
rect 27842 46001 27844 46053
rect 27788 45999 27844 46001
rect 27999 46053 28055 46055
rect 27999 46001 28001 46053
rect 28001 46001 28053 46053
rect 28053 46001 28055 46053
rect 27999 45999 28055 46001
rect 28210 46053 28266 46055
rect 28210 46001 28212 46053
rect 28212 46001 28264 46053
rect 28264 46001 28266 46053
rect 28210 45999 28266 46001
rect 28421 46053 28477 46055
rect 28421 46001 28423 46053
rect 28423 46001 28475 46053
rect 28475 46001 28477 46053
rect 28421 45999 28477 46001
rect 28632 46053 28688 46055
rect 28632 46001 28634 46053
rect 28634 46001 28686 46053
rect 28686 46001 28688 46053
rect 28632 45999 28688 46001
rect 28843 46053 28899 46055
rect 28843 46001 28845 46053
rect 28845 46001 28897 46053
rect 28897 46001 28899 46053
rect 28843 45999 28899 46001
rect 29054 46053 29110 46055
rect 29054 46001 29056 46053
rect 29056 46001 29108 46053
rect 29108 46001 29110 46053
rect 29054 45999 29110 46001
rect 29580 45153 29636 45155
rect 29580 45101 29582 45153
rect 29582 45101 29634 45153
rect 29634 45101 29636 45153
rect 29580 45099 29636 45101
rect 29791 45153 29847 45155
rect 29791 45101 29793 45153
rect 29793 45101 29845 45153
rect 29845 45101 29847 45153
rect 29791 45099 29847 45101
rect 30003 45153 30059 45155
rect 30003 45101 30005 45153
rect 30005 45101 30057 45153
rect 30057 45101 30059 45153
rect 30003 45099 30059 45101
rect 30214 45153 30270 45155
rect 30214 45101 30216 45153
rect 30216 45101 30268 45153
rect 30268 45101 30270 45153
rect 30214 45099 30270 45101
rect 27788 44253 27844 44255
rect 27788 44201 27790 44253
rect 27790 44201 27842 44253
rect 27842 44201 27844 44253
rect 27788 44199 27844 44201
rect 27999 44253 28055 44255
rect 27999 44201 28001 44253
rect 28001 44201 28053 44253
rect 28053 44201 28055 44253
rect 27999 44199 28055 44201
rect 28210 44253 28266 44255
rect 28210 44201 28212 44253
rect 28212 44201 28264 44253
rect 28264 44201 28266 44253
rect 28210 44199 28266 44201
rect 28421 44253 28477 44255
rect 28421 44201 28423 44253
rect 28423 44201 28475 44253
rect 28475 44201 28477 44253
rect 28421 44199 28477 44201
rect 28632 44253 28688 44255
rect 28632 44201 28634 44253
rect 28634 44201 28686 44253
rect 28686 44201 28688 44253
rect 28632 44199 28688 44201
rect 28843 44253 28899 44255
rect 28843 44201 28845 44253
rect 28845 44201 28897 44253
rect 28897 44201 28899 44253
rect 28843 44199 28899 44201
rect 29054 44253 29110 44255
rect 29054 44201 29056 44253
rect 29056 44201 29108 44253
rect 29108 44201 29110 44253
rect 29054 44199 29110 44201
rect 29580 43353 29636 43355
rect 29580 43301 29582 43353
rect 29582 43301 29634 43353
rect 29634 43301 29636 43353
rect 29580 43299 29636 43301
rect 29791 43353 29847 43355
rect 29791 43301 29793 43353
rect 29793 43301 29845 43353
rect 29845 43301 29847 43353
rect 29791 43299 29847 43301
rect 30003 43353 30059 43355
rect 30003 43301 30005 43353
rect 30005 43301 30057 43353
rect 30057 43301 30059 43353
rect 30003 43299 30059 43301
rect 30214 43353 30270 43355
rect 30214 43301 30216 43353
rect 30216 43301 30268 43353
rect 30268 43301 30270 43353
rect 30214 43299 30270 43301
rect 27788 42453 27844 42455
rect 27788 42401 27790 42453
rect 27790 42401 27842 42453
rect 27842 42401 27844 42453
rect 27788 42399 27844 42401
rect 27999 42453 28055 42455
rect 27999 42401 28001 42453
rect 28001 42401 28053 42453
rect 28053 42401 28055 42453
rect 27999 42399 28055 42401
rect 28210 42453 28266 42455
rect 28210 42401 28212 42453
rect 28212 42401 28264 42453
rect 28264 42401 28266 42453
rect 28210 42399 28266 42401
rect 28421 42453 28477 42455
rect 28421 42401 28423 42453
rect 28423 42401 28475 42453
rect 28475 42401 28477 42453
rect 28421 42399 28477 42401
rect 28632 42453 28688 42455
rect 28632 42401 28634 42453
rect 28634 42401 28686 42453
rect 28686 42401 28688 42453
rect 28632 42399 28688 42401
rect 28843 42453 28899 42455
rect 28843 42401 28845 42453
rect 28845 42401 28897 42453
rect 28897 42401 28899 42453
rect 28843 42399 28899 42401
rect 29054 42453 29110 42455
rect 29054 42401 29056 42453
rect 29056 42401 29108 42453
rect 29108 42401 29110 42453
rect 29054 42399 29110 42401
rect 29580 41553 29636 41555
rect 29580 41501 29582 41553
rect 29582 41501 29634 41553
rect 29634 41501 29636 41553
rect 29580 41499 29636 41501
rect 29791 41553 29847 41555
rect 29791 41501 29793 41553
rect 29793 41501 29845 41553
rect 29845 41501 29847 41553
rect 29791 41499 29847 41501
rect 30003 41553 30059 41555
rect 30003 41501 30005 41553
rect 30005 41501 30057 41553
rect 30057 41501 30059 41553
rect 30003 41499 30059 41501
rect 30214 41553 30270 41555
rect 30214 41501 30216 41553
rect 30216 41501 30268 41553
rect 30268 41501 30270 41553
rect 30214 41499 30270 41501
rect 27788 40653 27844 40655
rect 27788 40601 27790 40653
rect 27790 40601 27842 40653
rect 27842 40601 27844 40653
rect 27788 40599 27844 40601
rect 27999 40653 28055 40655
rect 27999 40601 28001 40653
rect 28001 40601 28053 40653
rect 28053 40601 28055 40653
rect 27999 40599 28055 40601
rect 28210 40653 28266 40655
rect 28210 40601 28212 40653
rect 28212 40601 28264 40653
rect 28264 40601 28266 40653
rect 28210 40599 28266 40601
rect 28421 40653 28477 40655
rect 28421 40601 28423 40653
rect 28423 40601 28475 40653
rect 28475 40601 28477 40653
rect 28421 40599 28477 40601
rect 28632 40653 28688 40655
rect 28632 40601 28634 40653
rect 28634 40601 28686 40653
rect 28686 40601 28688 40653
rect 28632 40599 28688 40601
rect 28843 40653 28899 40655
rect 28843 40601 28845 40653
rect 28845 40601 28897 40653
rect 28897 40601 28899 40653
rect 28843 40599 28899 40601
rect 29054 40653 29110 40655
rect 29054 40601 29056 40653
rect 29056 40601 29108 40653
rect 29108 40601 29110 40653
rect 29054 40599 29110 40601
rect 29580 39753 29636 39755
rect 29580 39701 29582 39753
rect 29582 39701 29634 39753
rect 29634 39701 29636 39753
rect 29580 39699 29636 39701
rect 29791 39753 29847 39755
rect 29791 39701 29793 39753
rect 29793 39701 29845 39753
rect 29845 39701 29847 39753
rect 29791 39699 29847 39701
rect 30003 39753 30059 39755
rect 30003 39701 30005 39753
rect 30005 39701 30057 39753
rect 30057 39701 30059 39753
rect 30003 39699 30059 39701
rect 30214 39753 30270 39755
rect 30214 39701 30216 39753
rect 30216 39701 30268 39753
rect 30268 39701 30270 39753
rect 30214 39699 30270 39701
rect 27788 38853 27844 38855
rect 27788 38801 27790 38853
rect 27790 38801 27842 38853
rect 27842 38801 27844 38853
rect 27788 38799 27844 38801
rect 27999 38853 28055 38855
rect 27999 38801 28001 38853
rect 28001 38801 28053 38853
rect 28053 38801 28055 38853
rect 27999 38799 28055 38801
rect 28210 38853 28266 38855
rect 28210 38801 28212 38853
rect 28212 38801 28264 38853
rect 28264 38801 28266 38853
rect 28210 38799 28266 38801
rect 28421 38853 28477 38855
rect 28421 38801 28423 38853
rect 28423 38801 28475 38853
rect 28475 38801 28477 38853
rect 28421 38799 28477 38801
rect 28632 38853 28688 38855
rect 28632 38801 28634 38853
rect 28634 38801 28686 38853
rect 28686 38801 28688 38853
rect 28632 38799 28688 38801
rect 28843 38853 28899 38855
rect 28843 38801 28845 38853
rect 28845 38801 28897 38853
rect 28897 38801 28899 38853
rect 28843 38799 28899 38801
rect 29054 38853 29110 38855
rect 29054 38801 29056 38853
rect 29056 38801 29108 38853
rect 29108 38801 29110 38853
rect 29054 38799 29110 38801
rect 29580 37953 29636 37955
rect 29580 37901 29582 37953
rect 29582 37901 29634 37953
rect 29634 37901 29636 37953
rect 29580 37899 29636 37901
rect 29791 37953 29847 37955
rect 29791 37901 29793 37953
rect 29793 37901 29845 37953
rect 29845 37901 29847 37953
rect 29791 37899 29847 37901
rect 30003 37953 30059 37955
rect 30003 37901 30005 37953
rect 30005 37901 30057 37953
rect 30057 37901 30059 37953
rect 30003 37899 30059 37901
rect 30214 37953 30270 37955
rect 30214 37901 30216 37953
rect 30216 37901 30268 37953
rect 30268 37901 30270 37953
rect 30214 37899 30270 37901
rect 27788 37053 27844 37055
rect 27788 37001 27790 37053
rect 27790 37001 27842 37053
rect 27842 37001 27844 37053
rect 27788 36999 27844 37001
rect 27999 37053 28055 37055
rect 27999 37001 28001 37053
rect 28001 37001 28053 37053
rect 28053 37001 28055 37053
rect 27999 36999 28055 37001
rect 28210 37053 28266 37055
rect 28210 37001 28212 37053
rect 28212 37001 28264 37053
rect 28264 37001 28266 37053
rect 28210 36999 28266 37001
rect 28421 37053 28477 37055
rect 28421 37001 28423 37053
rect 28423 37001 28475 37053
rect 28475 37001 28477 37053
rect 28421 36999 28477 37001
rect 28632 37053 28688 37055
rect 28632 37001 28634 37053
rect 28634 37001 28686 37053
rect 28686 37001 28688 37053
rect 28632 36999 28688 37001
rect 28843 37053 28899 37055
rect 28843 37001 28845 37053
rect 28845 37001 28897 37053
rect 28897 37001 28899 37053
rect 28843 36999 28899 37001
rect 29054 37053 29110 37055
rect 29054 37001 29056 37053
rect 29056 37001 29108 37053
rect 29108 37001 29110 37053
rect 29054 36999 29110 37001
rect 29580 36153 29636 36155
rect 29580 36101 29582 36153
rect 29582 36101 29634 36153
rect 29634 36101 29636 36153
rect 29580 36099 29636 36101
rect 29791 36153 29847 36155
rect 29791 36101 29793 36153
rect 29793 36101 29845 36153
rect 29845 36101 29847 36153
rect 29791 36099 29847 36101
rect 30003 36153 30059 36155
rect 30003 36101 30005 36153
rect 30005 36101 30057 36153
rect 30057 36101 30059 36153
rect 30003 36099 30059 36101
rect 30214 36153 30270 36155
rect 30214 36101 30216 36153
rect 30216 36101 30268 36153
rect 30268 36101 30270 36153
rect 30214 36099 30270 36101
rect 30852 64901 30854 64953
rect 30854 64901 30906 64953
rect 30906 64901 30908 64953
rect 30852 64899 30908 64901
rect 31063 64953 31119 64955
rect 31063 64901 31065 64953
rect 31065 64901 31117 64953
rect 31117 64901 31119 64953
rect 31063 64899 31119 64901
rect 31274 64953 31330 64955
rect 31274 64901 31276 64953
rect 31276 64901 31328 64953
rect 31328 64901 31330 64953
rect 31274 64899 31330 64901
rect 31484 64953 31540 64955
rect 31484 64901 31486 64953
rect 31486 64901 31538 64953
rect 31538 64901 31540 64953
rect 31484 64899 31540 64901
rect 31695 64953 31751 64955
rect 31695 64901 31697 64953
rect 31697 64901 31749 64953
rect 31749 64901 31751 64953
rect 31695 64899 31751 64901
rect 31907 64953 31963 64955
rect 31907 64901 31909 64953
rect 31909 64901 31961 64953
rect 31961 64901 31963 64953
rect 31907 64899 31963 64901
rect 32118 64953 32174 64955
rect 32118 64901 32120 64953
rect 32120 64901 32172 64953
rect 32172 64901 32174 64953
rect 32118 64899 32174 64901
rect 32328 64953 32384 64955
rect 32328 64901 32330 64953
rect 32330 64901 32382 64953
rect 32382 64901 32384 64953
rect 32328 64899 32384 64901
rect 32539 64953 32595 64955
rect 32539 64901 32541 64953
rect 32541 64901 32593 64953
rect 32593 64901 32595 64953
rect 32539 64899 32595 64901
rect 32750 64953 32806 64955
rect 32750 64901 32752 64953
rect 32752 64901 32804 64953
rect 32804 64901 32806 64953
rect 32750 64899 32806 64901
rect 35218 64953 35274 64955
rect 33055 64466 33111 64522
rect 33235 64466 33291 64522
rect 33817 64459 33873 64515
rect 33997 64459 34053 64515
rect 34282 63999 34338 64055
rect 34493 63999 34549 64055
rect 34705 64053 34761 64055
rect 34916 64053 34972 64055
rect 34705 64001 34755 64053
rect 34755 64001 34761 64053
rect 34916 64001 34935 64053
rect 34935 64001 34972 64053
rect 34705 63999 34761 64001
rect 34916 63999 34972 64001
rect 33055 63532 33111 63588
rect 33235 63532 33291 63588
rect 33817 63539 33873 63595
rect 33997 63539 34053 63595
rect 30852 63153 30908 63155
rect 30852 63101 30854 63153
rect 30854 63101 30906 63153
rect 30906 63101 30908 63153
rect 30852 63099 30908 63101
rect 31063 63153 31119 63155
rect 31063 63101 31065 63153
rect 31065 63101 31117 63153
rect 31117 63101 31119 63153
rect 31063 63099 31119 63101
rect 31274 63153 31330 63155
rect 31274 63101 31276 63153
rect 31276 63101 31328 63153
rect 31328 63101 31330 63153
rect 31274 63099 31330 63101
rect 31484 63153 31540 63155
rect 31484 63101 31486 63153
rect 31486 63101 31538 63153
rect 31538 63101 31540 63153
rect 31484 63099 31540 63101
rect 31695 63153 31751 63155
rect 31695 63101 31697 63153
rect 31697 63101 31749 63153
rect 31749 63101 31751 63153
rect 31695 63099 31751 63101
rect 31907 63153 31963 63155
rect 31907 63101 31909 63153
rect 31909 63101 31961 63153
rect 31961 63101 31963 63153
rect 31907 63099 31963 63101
rect 32118 63153 32174 63155
rect 32118 63101 32120 63153
rect 32120 63101 32172 63153
rect 32172 63101 32174 63153
rect 32118 63099 32174 63101
rect 32328 63153 32384 63155
rect 32328 63101 32330 63153
rect 32330 63101 32382 63153
rect 32382 63101 32384 63153
rect 32328 63099 32384 63101
rect 32539 63153 32595 63155
rect 32539 63101 32541 63153
rect 32541 63101 32593 63153
rect 32593 63101 32595 63153
rect 32539 63099 32595 63101
rect 32750 63153 32806 63155
rect 32750 63101 32752 63153
rect 32752 63101 32804 63153
rect 32804 63101 32806 63153
rect 32750 63099 32806 63101
rect 33055 62666 33111 62722
rect 33235 62666 33291 62722
rect 33817 62659 33873 62715
rect 33997 62659 34053 62715
rect 34282 62199 34338 62255
rect 34493 62199 34549 62255
rect 34705 62253 34761 62255
rect 34916 62253 34972 62255
rect 34705 62201 34755 62253
rect 34755 62201 34761 62253
rect 34916 62201 34935 62253
rect 34935 62201 34972 62253
rect 34705 62199 34761 62201
rect 34916 62199 34972 62201
rect 33055 61732 33111 61788
rect 33235 61732 33291 61788
rect 33817 61739 33873 61795
rect 33997 61739 34053 61795
rect 30852 61353 30908 61355
rect 30852 61301 30854 61353
rect 30854 61301 30906 61353
rect 30906 61301 30908 61353
rect 30852 61299 30908 61301
rect 31063 61353 31119 61355
rect 31063 61301 31065 61353
rect 31065 61301 31117 61353
rect 31117 61301 31119 61353
rect 31063 61299 31119 61301
rect 31274 61353 31330 61355
rect 31274 61301 31276 61353
rect 31276 61301 31328 61353
rect 31328 61301 31330 61353
rect 31274 61299 31330 61301
rect 31484 61353 31540 61355
rect 31484 61301 31486 61353
rect 31486 61301 31538 61353
rect 31538 61301 31540 61353
rect 31484 61299 31540 61301
rect 31695 61353 31751 61355
rect 31695 61301 31697 61353
rect 31697 61301 31749 61353
rect 31749 61301 31751 61353
rect 31695 61299 31751 61301
rect 31907 61353 31963 61355
rect 31907 61301 31909 61353
rect 31909 61301 31961 61353
rect 31961 61301 31963 61353
rect 31907 61299 31963 61301
rect 32118 61353 32174 61355
rect 32118 61301 32120 61353
rect 32120 61301 32172 61353
rect 32172 61301 32174 61353
rect 32118 61299 32174 61301
rect 32328 61353 32384 61355
rect 32328 61301 32330 61353
rect 32330 61301 32382 61353
rect 32382 61301 32384 61353
rect 32328 61299 32384 61301
rect 32539 61353 32595 61355
rect 32539 61301 32541 61353
rect 32541 61301 32593 61353
rect 32593 61301 32595 61353
rect 32539 61299 32595 61301
rect 32750 61353 32806 61355
rect 32750 61301 32752 61353
rect 32752 61301 32804 61353
rect 32804 61301 32806 61353
rect 32750 61299 32806 61301
rect 33055 60866 33111 60922
rect 33235 60866 33291 60922
rect 33817 60859 33873 60915
rect 33997 60859 34053 60915
rect 34282 60399 34338 60455
rect 34493 60399 34549 60455
rect 34705 60453 34761 60455
rect 34916 60453 34972 60455
rect 34705 60401 34755 60453
rect 34755 60401 34761 60453
rect 34916 60401 34935 60453
rect 34935 60401 34972 60453
rect 34705 60399 34761 60401
rect 34916 60399 34972 60401
rect 33055 59932 33111 59988
rect 33235 59932 33291 59988
rect 33817 59939 33873 59995
rect 33997 59939 34053 59995
rect 30852 59553 30908 59555
rect 30852 59501 30854 59553
rect 30854 59501 30906 59553
rect 30906 59501 30908 59553
rect 30852 59499 30908 59501
rect 31063 59553 31119 59555
rect 31063 59501 31065 59553
rect 31065 59501 31117 59553
rect 31117 59501 31119 59553
rect 31063 59499 31119 59501
rect 31274 59553 31330 59555
rect 31274 59501 31276 59553
rect 31276 59501 31328 59553
rect 31328 59501 31330 59553
rect 31274 59499 31330 59501
rect 31484 59553 31540 59555
rect 31484 59501 31486 59553
rect 31486 59501 31538 59553
rect 31538 59501 31540 59553
rect 31484 59499 31540 59501
rect 31695 59553 31751 59555
rect 31695 59501 31697 59553
rect 31697 59501 31749 59553
rect 31749 59501 31751 59553
rect 31695 59499 31751 59501
rect 31907 59553 31963 59555
rect 31907 59501 31909 59553
rect 31909 59501 31961 59553
rect 31961 59501 31963 59553
rect 31907 59499 31963 59501
rect 32118 59553 32174 59555
rect 32118 59501 32120 59553
rect 32120 59501 32172 59553
rect 32172 59501 32174 59553
rect 32118 59499 32174 59501
rect 32328 59553 32384 59555
rect 32328 59501 32330 59553
rect 32330 59501 32382 59553
rect 32382 59501 32384 59553
rect 32328 59499 32384 59501
rect 32539 59553 32595 59555
rect 32539 59501 32541 59553
rect 32541 59501 32593 59553
rect 32593 59501 32595 59553
rect 32539 59499 32595 59501
rect 32750 59553 32806 59555
rect 32750 59501 32752 59553
rect 32752 59501 32804 59553
rect 32804 59501 32806 59553
rect 32750 59499 32806 59501
rect 33055 59066 33111 59122
rect 33235 59066 33291 59122
rect 33817 59059 33873 59115
rect 33997 59059 34053 59115
rect 34282 58599 34338 58655
rect 34493 58599 34549 58655
rect 34705 58653 34761 58655
rect 34916 58653 34972 58655
rect 34705 58601 34755 58653
rect 34755 58601 34761 58653
rect 34916 58601 34935 58653
rect 34935 58601 34972 58653
rect 34705 58599 34761 58601
rect 34916 58599 34972 58601
rect 33055 58132 33111 58188
rect 33235 58132 33291 58188
rect 33817 58139 33873 58195
rect 33997 58139 34053 58195
rect 30852 57753 30908 57755
rect 30852 57701 30854 57753
rect 30854 57701 30906 57753
rect 30906 57701 30908 57753
rect 30852 57699 30908 57701
rect 31063 57753 31119 57755
rect 31063 57701 31065 57753
rect 31065 57701 31117 57753
rect 31117 57701 31119 57753
rect 31063 57699 31119 57701
rect 31274 57753 31330 57755
rect 31274 57701 31276 57753
rect 31276 57701 31328 57753
rect 31328 57701 31330 57753
rect 31274 57699 31330 57701
rect 31484 57753 31540 57755
rect 31484 57701 31486 57753
rect 31486 57701 31538 57753
rect 31538 57701 31540 57753
rect 31484 57699 31540 57701
rect 31695 57753 31751 57755
rect 31695 57701 31697 57753
rect 31697 57701 31749 57753
rect 31749 57701 31751 57753
rect 31695 57699 31751 57701
rect 31907 57753 31963 57755
rect 31907 57701 31909 57753
rect 31909 57701 31961 57753
rect 31961 57701 31963 57753
rect 31907 57699 31963 57701
rect 32118 57753 32174 57755
rect 32118 57701 32120 57753
rect 32120 57701 32172 57753
rect 32172 57701 32174 57753
rect 32118 57699 32174 57701
rect 32328 57753 32384 57755
rect 32328 57701 32330 57753
rect 32330 57701 32382 57753
rect 32382 57701 32384 57753
rect 32328 57699 32384 57701
rect 32539 57753 32595 57755
rect 32539 57701 32541 57753
rect 32541 57701 32593 57753
rect 32593 57701 32595 57753
rect 32539 57699 32595 57701
rect 32750 57753 32806 57755
rect 32750 57701 32752 57753
rect 32752 57701 32804 57753
rect 32804 57701 32806 57753
rect 32750 57699 32806 57701
rect 33055 57266 33111 57322
rect 33235 57266 33291 57322
rect 33817 57259 33873 57315
rect 33997 57259 34053 57315
rect 34282 56799 34338 56855
rect 34493 56799 34549 56855
rect 34705 56853 34761 56855
rect 34916 56853 34972 56855
rect 34705 56801 34755 56853
rect 34755 56801 34761 56853
rect 34916 56801 34935 56853
rect 34935 56801 34972 56853
rect 34705 56799 34761 56801
rect 34916 56799 34972 56801
rect 33055 56332 33111 56388
rect 33235 56332 33291 56388
rect 33817 56339 33873 56395
rect 33997 56339 34053 56395
rect 30852 55953 30908 55955
rect 30852 55901 30854 55953
rect 30854 55901 30906 55953
rect 30906 55901 30908 55953
rect 30852 55899 30908 55901
rect 31063 55953 31119 55955
rect 31063 55901 31065 55953
rect 31065 55901 31117 55953
rect 31117 55901 31119 55953
rect 31063 55899 31119 55901
rect 31274 55953 31330 55955
rect 31274 55901 31276 55953
rect 31276 55901 31328 55953
rect 31328 55901 31330 55953
rect 31274 55899 31330 55901
rect 31484 55953 31540 55955
rect 31484 55901 31486 55953
rect 31486 55901 31538 55953
rect 31538 55901 31540 55953
rect 31484 55899 31540 55901
rect 31695 55953 31751 55955
rect 31695 55901 31697 55953
rect 31697 55901 31749 55953
rect 31749 55901 31751 55953
rect 31695 55899 31751 55901
rect 31907 55953 31963 55955
rect 31907 55901 31909 55953
rect 31909 55901 31961 55953
rect 31961 55901 31963 55953
rect 31907 55899 31963 55901
rect 32118 55953 32174 55955
rect 32118 55901 32120 55953
rect 32120 55901 32172 55953
rect 32172 55901 32174 55953
rect 32118 55899 32174 55901
rect 32328 55953 32384 55955
rect 32328 55901 32330 55953
rect 32330 55901 32382 55953
rect 32382 55901 32384 55953
rect 32328 55899 32384 55901
rect 32539 55953 32595 55955
rect 32539 55901 32541 55953
rect 32541 55901 32593 55953
rect 32593 55901 32595 55953
rect 32539 55899 32595 55901
rect 32750 55953 32806 55955
rect 32750 55901 32752 55953
rect 32752 55901 32804 55953
rect 32804 55901 32806 55953
rect 32750 55899 32806 55901
rect 33055 55466 33111 55522
rect 33235 55466 33291 55522
rect 33817 55459 33873 55515
rect 33997 55459 34053 55515
rect 34282 54999 34338 55055
rect 34493 54999 34549 55055
rect 34705 55053 34761 55055
rect 34916 55053 34972 55055
rect 34705 55001 34755 55053
rect 34755 55001 34761 55053
rect 34916 55001 34935 55053
rect 34935 55001 34972 55053
rect 34705 54999 34761 55001
rect 34916 54999 34972 55001
rect 33055 54532 33111 54588
rect 33235 54532 33291 54588
rect 33817 54539 33873 54595
rect 33997 54539 34053 54595
rect 30852 54153 30908 54155
rect 30852 54101 30854 54153
rect 30854 54101 30906 54153
rect 30906 54101 30908 54153
rect 30852 54099 30908 54101
rect 31063 54153 31119 54155
rect 31063 54101 31065 54153
rect 31065 54101 31117 54153
rect 31117 54101 31119 54153
rect 31063 54099 31119 54101
rect 31274 54153 31330 54155
rect 31274 54101 31276 54153
rect 31276 54101 31328 54153
rect 31328 54101 31330 54153
rect 31274 54099 31330 54101
rect 31484 54153 31540 54155
rect 31484 54101 31486 54153
rect 31486 54101 31538 54153
rect 31538 54101 31540 54153
rect 31484 54099 31540 54101
rect 31695 54153 31751 54155
rect 31695 54101 31697 54153
rect 31697 54101 31749 54153
rect 31749 54101 31751 54153
rect 31695 54099 31751 54101
rect 31907 54153 31963 54155
rect 31907 54101 31909 54153
rect 31909 54101 31961 54153
rect 31961 54101 31963 54153
rect 31907 54099 31963 54101
rect 32118 54153 32174 54155
rect 32118 54101 32120 54153
rect 32120 54101 32172 54153
rect 32172 54101 32174 54153
rect 32118 54099 32174 54101
rect 32328 54153 32384 54155
rect 32328 54101 32330 54153
rect 32330 54101 32382 54153
rect 32382 54101 32384 54153
rect 32328 54099 32384 54101
rect 32539 54153 32595 54155
rect 32539 54101 32541 54153
rect 32541 54101 32593 54153
rect 32593 54101 32595 54153
rect 32539 54099 32595 54101
rect 32750 54153 32806 54155
rect 32750 54101 32752 54153
rect 32752 54101 32804 54153
rect 32804 54101 32806 54153
rect 32750 54099 32806 54101
rect 33055 53666 33111 53722
rect 33235 53666 33291 53722
rect 33817 53659 33873 53715
rect 33997 53659 34053 53715
rect 34282 53199 34338 53255
rect 34493 53199 34549 53255
rect 34705 53253 34761 53255
rect 34916 53253 34972 53255
rect 34705 53201 34755 53253
rect 34755 53201 34761 53253
rect 34916 53201 34935 53253
rect 34935 53201 34972 53253
rect 34705 53199 34761 53201
rect 34916 53199 34972 53201
rect 33055 52732 33111 52788
rect 33235 52732 33291 52788
rect 33817 52739 33873 52795
rect 33997 52739 34053 52795
rect 30852 52353 30908 52355
rect 30852 52301 30854 52353
rect 30854 52301 30906 52353
rect 30906 52301 30908 52353
rect 30852 52299 30908 52301
rect 31063 52353 31119 52355
rect 31063 52301 31065 52353
rect 31065 52301 31117 52353
rect 31117 52301 31119 52353
rect 31063 52299 31119 52301
rect 31274 52353 31330 52355
rect 31274 52301 31276 52353
rect 31276 52301 31328 52353
rect 31328 52301 31330 52353
rect 31274 52299 31330 52301
rect 31484 52353 31540 52355
rect 31484 52301 31486 52353
rect 31486 52301 31538 52353
rect 31538 52301 31540 52353
rect 31484 52299 31540 52301
rect 31695 52353 31751 52355
rect 31695 52301 31697 52353
rect 31697 52301 31749 52353
rect 31749 52301 31751 52353
rect 31695 52299 31751 52301
rect 31907 52353 31963 52355
rect 31907 52301 31909 52353
rect 31909 52301 31961 52353
rect 31961 52301 31963 52353
rect 31907 52299 31963 52301
rect 32118 52353 32174 52355
rect 32118 52301 32120 52353
rect 32120 52301 32172 52353
rect 32172 52301 32174 52353
rect 32118 52299 32174 52301
rect 32328 52353 32384 52355
rect 32328 52301 32330 52353
rect 32330 52301 32382 52353
rect 32382 52301 32384 52353
rect 32328 52299 32384 52301
rect 32539 52353 32595 52355
rect 32539 52301 32541 52353
rect 32541 52301 32593 52353
rect 32593 52301 32595 52353
rect 32539 52299 32595 52301
rect 32750 52353 32806 52355
rect 32750 52301 32752 52353
rect 32752 52301 32804 52353
rect 32804 52301 32806 52353
rect 32750 52299 32806 52301
rect 33055 51866 33111 51922
rect 33235 51866 33291 51922
rect 33817 51859 33873 51915
rect 33997 51859 34053 51915
rect 34282 51399 34338 51455
rect 34493 51399 34549 51455
rect 34705 51453 34761 51455
rect 34916 51453 34972 51455
rect 34705 51401 34755 51453
rect 34755 51401 34761 51453
rect 34916 51401 34935 51453
rect 34935 51401 34972 51453
rect 34705 51399 34761 51401
rect 34916 51399 34972 51401
rect 33055 50932 33111 50988
rect 33235 50932 33291 50988
rect 33817 50939 33873 50995
rect 33997 50939 34053 50995
rect 30852 50553 30908 50555
rect 30852 50501 30854 50553
rect 30854 50501 30906 50553
rect 30906 50501 30908 50553
rect 30852 50499 30908 50501
rect 31063 50553 31119 50555
rect 31063 50501 31065 50553
rect 31065 50501 31117 50553
rect 31117 50501 31119 50553
rect 31063 50499 31119 50501
rect 31274 50553 31330 50555
rect 31274 50501 31276 50553
rect 31276 50501 31328 50553
rect 31328 50501 31330 50553
rect 31274 50499 31330 50501
rect 31484 50553 31540 50555
rect 31484 50501 31486 50553
rect 31486 50501 31538 50553
rect 31538 50501 31540 50553
rect 31484 50499 31540 50501
rect 31695 50553 31751 50555
rect 31695 50501 31697 50553
rect 31697 50501 31749 50553
rect 31749 50501 31751 50553
rect 31695 50499 31751 50501
rect 31907 50553 31963 50555
rect 31907 50501 31909 50553
rect 31909 50501 31961 50553
rect 31961 50501 31963 50553
rect 31907 50499 31963 50501
rect 32118 50553 32174 50555
rect 32118 50501 32120 50553
rect 32120 50501 32172 50553
rect 32172 50501 32174 50553
rect 32118 50499 32174 50501
rect 32328 50553 32384 50555
rect 32328 50501 32330 50553
rect 32330 50501 32382 50553
rect 32382 50501 32384 50553
rect 32328 50499 32384 50501
rect 32539 50553 32595 50555
rect 32539 50501 32541 50553
rect 32541 50501 32593 50553
rect 32593 50501 32595 50553
rect 32539 50499 32595 50501
rect 32750 50553 32806 50555
rect 32750 50501 32752 50553
rect 32752 50501 32804 50553
rect 32804 50501 32806 50553
rect 32750 50499 32806 50501
rect 33055 50066 33111 50122
rect 33235 50066 33291 50122
rect 33817 50059 33873 50115
rect 33997 50059 34053 50115
rect 34282 49599 34338 49655
rect 34493 49599 34549 49655
rect 34705 49653 34761 49655
rect 34916 49653 34972 49655
rect 34705 49601 34755 49653
rect 34755 49601 34761 49653
rect 34916 49601 34935 49653
rect 34935 49601 34972 49653
rect 34705 49599 34761 49601
rect 34916 49599 34972 49601
rect 33055 49132 33111 49188
rect 33235 49132 33291 49188
rect 33817 49139 33873 49195
rect 33997 49139 34053 49195
rect 30852 48753 30908 48755
rect 30852 48701 30854 48753
rect 30854 48701 30906 48753
rect 30906 48701 30908 48753
rect 30852 48699 30908 48701
rect 31063 48753 31119 48755
rect 31063 48701 31065 48753
rect 31065 48701 31117 48753
rect 31117 48701 31119 48753
rect 31063 48699 31119 48701
rect 31274 48753 31330 48755
rect 31274 48701 31276 48753
rect 31276 48701 31328 48753
rect 31328 48701 31330 48753
rect 31274 48699 31330 48701
rect 31484 48753 31540 48755
rect 31484 48701 31486 48753
rect 31486 48701 31538 48753
rect 31538 48701 31540 48753
rect 31484 48699 31540 48701
rect 31695 48753 31751 48755
rect 31695 48701 31697 48753
rect 31697 48701 31749 48753
rect 31749 48701 31751 48753
rect 31695 48699 31751 48701
rect 31907 48753 31963 48755
rect 31907 48701 31909 48753
rect 31909 48701 31961 48753
rect 31961 48701 31963 48753
rect 31907 48699 31963 48701
rect 32118 48753 32174 48755
rect 32118 48701 32120 48753
rect 32120 48701 32172 48753
rect 32172 48701 32174 48753
rect 32118 48699 32174 48701
rect 32328 48753 32384 48755
rect 32328 48701 32330 48753
rect 32330 48701 32382 48753
rect 32382 48701 32384 48753
rect 32328 48699 32384 48701
rect 32539 48753 32595 48755
rect 32539 48701 32541 48753
rect 32541 48701 32593 48753
rect 32593 48701 32595 48753
rect 32539 48699 32595 48701
rect 32750 48753 32806 48755
rect 32750 48701 32752 48753
rect 32752 48701 32804 48753
rect 32804 48701 32806 48753
rect 32750 48699 32806 48701
rect 33055 48266 33111 48322
rect 33235 48266 33291 48322
rect 33817 48259 33873 48315
rect 33997 48259 34053 48315
rect 34282 47799 34338 47855
rect 34493 47799 34549 47855
rect 34705 47853 34761 47855
rect 34916 47853 34972 47855
rect 34705 47801 34755 47853
rect 34755 47801 34761 47853
rect 34916 47801 34935 47853
rect 34935 47801 34972 47853
rect 34705 47799 34761 47801
rect 34916 47799 34972 47801
rect 33055 47332 33111 47388
rect 33235 47332 33291 47388
rect 33817 47339 33873 47395
rect 33997 47339 34053 47395
rect 30852 46953 30908 46955
rect 30852 46901 30854 46953
rect 30854 46901 30906 46953
rect 30906 46901 30908 46953
rect 30852 46899 30908 46901
rect 31063 46953 31119 46955
rect 31063 46901 31065 46953
rect 31065 46901 31117 46953
rect 31117 46901 31119 46953
rect 31063 46899 31119 46901
rect 31274 46953 31330 46955
rect 31274 46901 31276 46953
rect 31276 46901 31328 46953
rect 31328 46901 31330 46953
rect 31274 46899 31330 46901
rect 31484 46953 31540 46955
rect 31484 46901 31486 46953
rect 31486 46901 31538 46953
rect 31538 46901 31540 46953
rect 31484 46899 31540 46901
rect 31695 46953 31751 46955
rect 31695 46901 31697 46953
rect 31697 46901 31749 46953
rect 31749 46901 31751 46953
rect 31695 46899 31751 46901
rect 31907 46953 31963 46955
rect 31907 46901 31909 46953
rect 31909 46901 31961 46953
rect 31961 46901 31963 46953
rect 31907 46899 31963 46901
rect 32118 46953 32174 46955
rect 32118 46901 32120 46953
rect 32120 46901 32172 46953
rect 32172 46901 32174 46953
rect 32118 46899 32174 46901
rect 32328 46953 32384 46955
rect 32328 46901 32330 46953
rect 32330 46901 32382 46953
rect 32382 46901 32384 46953
rect 32328 46899 32384 46901
rect 32539 46953 32595 46955
rect 32539 46901 32541 46953
rect 32541 46901 32593 46953
rect 32593 46901 32595 46953
rect 32539 46899 32595 46901
rect 32750 46953 32806 46955
rect 32750 46901 32752 46953
rect 32752 46901 32804 46953
rect 32804 46901 32806 46953
rect 32750 46899 32806 46901
rect 33055 46466 33111 46522
rect 33235 46466 33291 46522
rect 33817 46459 33873 46515
rect 33997 46459 34053 46515
rect 34282 45999 34338 46055
rect 34493 45999 34549 46055
rect 34705 46053 34761 46055
rect 34916 46053 34972 46055
rect 34705 46001 34755 46053
rect 34755 46001 34761 46053
rect 34916 46001 34935 46053
rect 34935 46001 34972 46053
rect 34705 45999 34761 46001
rect 34916 45999 34972 46001
rect 33055 45532 33111 45588
rect 33235 45532 33291 45588
rect 33817 45539 33873 45595
rect 33997 45539 34053 45595
rect 30852 45153 30908 45155
rect 30852 45101 30854 45153
rect 30854 45101 30906 45153
rect 30906 45101 30908 45153
rect 30852 45099 30908 45101
rect 31063 45153 31119 45155
rect 31063 45101 31065 45153
rect 31065 45101 31117 45153
rect 31117 45101 31119 45153
rect 31063 45099 31119 45101
rect 31274 45153 31330 45155
rect 31274 45101 31276 45153
rect 31276 45101 31328 45153
rect 31328 45101 31330 45153
rect 31274 45099 31330 45101
rect 31484 45153 31540 45155
rect 31484 45101 31486 45153
rect 31486 45101 31538 45153
rect 31538 45101 31540 45153
rect 31484 45099 31540 45101
rect 31695 45153 31751 45155
rect 31695 45101 31697 45153
rect 31697 45101 31749 45153
rect 31749 45101 31751 45153
rect 31695 45099 31751 45101
rect 31907 45153 31963 45155
rect 31907 45101 31909 45153
rect 31909 45101 31961 45153
rect 31961 45101 31963 45153
rect 31907 45099 31963 45101
rect 32118 45153 32174 45155
rect 32118 45101 32120 45153
rect 32120 45101 32172 45153
rect 32172 45101 32174 45153
rect 32118 45099 32174 45101
rect 32328 45153 32384 45155
rect 32328 45101 32330 45153
rect 32330 45101 32382 45153
rect 32382 45101 32384 45153
rect 32328 45099 32384 45101
rect 32539 45153 32595 45155
rect 32539 45101 32541 45153
rect 32541 45101 32593 45153
rect 32593 45101 32595 45153
rect 32539 45099 32595 45101
rect 32750 45153 32806 45155
rect 32750 45101 32752 45153
rect 32752 45101 32804 45153
rect 32804 45101 32806 45153
rect 32750 45099 32806 45101
rect 33055 44666 33111 44722
rect 33235 44666 33291 44722
rect 33817 44659 33873 44715
rect 33997 44659 34053 44715
rect 34282 44199 34338 44255
rect 34493 44199 34549 44255
rect 34705 44253 34761 44255
rect 34916 44253 34972 44255
rect 34705 44201 34755 44253
rect 34755 44201 34761 44253
rect 34916 44201 34935 44253
rect 34935 44201 34972 44253
rect 34705 44199 34761 44201
rect 34916 44199 34972 44201
rect 33055 43732 33111 43788
rect 33235 43732 33291 43788
rect 33817 43739 33873 43795
rect 33997 43739 34053 43795
rect 30852 43353 30908 43355
rect 30852 43301 30854 43353
rect 30854 43301 30906 43353
rect 30906 43301 30908 43353
rect 30852 43299 30908 43301
rect 31063 43353 31119 43355
rect 31063 43301 31065 43353
rect 31065 43301 31117 43353
rect 31117 43301 31119 43353
rect 31063 43299 31119 43301
rect 31274 43353 31330 43355
rect 31274 43301 31276 43353
rect 31276 43301 31328 43353
rect 31328 43301 31330 43353
rect 31274 43299 31330 43301
rect 31484 43353 31540 43355
rect 31484 43301 31486 43353
rect 31486 43301 31538 43353
rect 31538 43301 31540 43353
rect 31484 43299 31540 43301
rect 31695 43353 31751 43355
rect 31695 43301 31697 43353
rect 31697 43301 31749 43353
rect 31749 43301 31751 43353
rect 31695 43299 31751 43301
rect 31907 43353 31963 43355
rect 31907 43301 31909 43353
rect 31909 43301 31961 43353
rect 31961 43301 31963 43353
rect 31907 43299 31963 43301
rect 32118 43353 32174 43355
rect 32118 43301 32120 43353
rect 32120 43301 32172 43353
rect 32172 43301 32174 43353
rect 32118 43299 32174 43301
rect 32328 43353 32384 43355
rect 32328 43301 32330 43353
rect 32330 43301 32382 43353
rect 32382 43301 32384 43353
rect 32328 43299 32384 43301
rect 32539 43353 32595 43355
rect 32539 43301 32541 43353
rect 32541 43301 32593 43353
rect 32593 43301 32595 43353
rect 32539 43299 32595 43301
rect 32750 43353 32806 43355
rect 32750 43301 32752 43353
rect 32752 43301 32804 43353
rect 32804 43301 32806 43353
rect 32750 43299 32806 43301
rect 33055 42866 33111 42922
rect 33235 42866 33291 42922
rect 33817 42859 33873 42915
rect 33997 42859 34053 42915
rect 34282 42399 34338 42455
rect 34493 42399 34549 42455
rect 34705 42453 34761 42455
rect 34916 42453 34972 42455
rect 34705 42401 34755 42453
rect 34755 42401 34761 42453
rect 34916 42401 34935 42453
rect 34935 42401 34972 42453
rect 34705 42399 34761 42401
rect 34916 42399 34972 42401
rect 33055 41932 33111 41988
rect 33235 41932 33291 41988
rect 33817 41939 33873 41995
rect 33997 41939 34053 41995
rect 30852 41553 30908 41555
rect 30852 41501 30854 41553
rect 30854 41501 30906 41553
rect 30906 41501 30908 41553
rect 30852 41499 30908 41501
rect 31063 41553 31119 41555
rect 31063 41501 31065 41553
rect 31065 41501 31117 41553
rect 31117 41501 31119 41553
rect 31063 41499 31119 41501
rect 31274 41553 31330 41555
rect 31274 41501 31276 41553
rect 31276 41501 31328 41553
rect 31328 41501 31330 41553
rect 31274 41499 31330 41501
rect 31484 41553 31540 41555
rect 31484 41501 31486 41553
rect 31486 41501 31538 41553
rect 31538 41501 31540 41553
rect 31484 41499 31540 41501
rect 31695 41553 31751 41555
rect 31695 41501 31697 41553
rect 31697 41501 31749 41553
rect 31749 41501 31751 41553
rect 31695 41499 31751 41501
rect 31907 41553 31963 41555
rect 31907 41501 31909 41553
rect 31909 41501 31961 41553
rect 31961 41501 31963 41553
rect 31907 41499 31963 41501
rect 32118 41553 32174 41555
rect 32118 41501 32120 41553
rect 32120 41501 32172 41553
rect 32172 41501 32174 41553
rect 32118 41499 32174 41501
rect 32328 41553 32384 41555
rect 32328 41501 32330 41553
rect 32330 41501 32382 41553
rect 32382 41501 32384 41553
rect 32328 41499 32384 41501
rect 32539 41553 32595 41555
rect 32539 41501 32541 41553
rect 32541 41501 32593 41553
rect 32593 41501 32595 41553
rect 32539 41499 32595 41501
rect 32750 41553 32806 41555
rect 32750 41501 32752 41553
rect 32752 41501 32804 41553
rect 32804 41501 32806 41553
rect 32750 41499 32806 41501
rect 33055 41066 33111 41122
rect 33235 41066 33291 41122
rect 33817 41059 33873 41115
rect 33997 41059 34053 41115
rect 34282 40599 34338 40655
rect 34493 40599 34549 40655
rect 34705 40653 34761 40655
rect 34916 40653 34972 40655
rect 34705 40601 34755 40653
rect 34755 40601 34761 40653
rect 34916 40601 34935 40653
rect 34935 40601 34972 40653
rect 34705 40599 34761 40601
rect 34916 40599 34972 40601
rect 33055 40132 33111 40188
rect 33235 40132 33291 40188
rect 33817 40139 33873 40195
rect 33997 40139 34053 40195
rect 30852 39753 30908 39755
rect 30852 39701 30854 39753
rect 30854 39701 30906 39753
rect 30906 39701 30908 39753
rect 30852 39699 30908 39701
rect 31063 39753 31119 39755
rect 31063 39701 31065 39753
rect 31065 39701 31117 39753
rect 31117 39701 31119 39753
rect 31063 39699 31119 39701
rect 31274 39753 31330 39755
rect 31274 39701 31276 39753
rect 31276 39701 31328 39753
rect 31328 39701 31330 39753
rect 31274 39699 31330 39701
rect 31484 39753 31540 39755
rect 31484 39701 31486 39753
rect 31486 39701 31538 39753
rect 31538 39701 31540 39753
rect 31484 39699 31540 39701
rect 31695 39753 31751 39755
rect 31695 39701 31697 39753
rect 31697 39701 31749 39753
rect 31749 39701 31751 39753
rect 31695 39699 31751 39701
rect 31907 39753 31963 39755
rect 31907 39701 31909 39753
rect 31909 39701 31961 39753
rect 31961 39701 31963 39753
rect 31907 39699 31963 39701
rect 32118 39753 32174 39755
rect 32118 39701 32120 39753
rect 32120 39701 32172 39753
rect 32172 39701 32174 39753
rect 32118 39699 32174 39701
rect 32328 39753 32384 39755
rect 32328 39701 32330 39753
rect 32330 39701 32382 39753
rect 32382 39701 32384 39753
rect 32328 39699 32384 39701
rect 32539 39753 32595 39755
rect 32539 39701 32541 39753
rect 32541 39701 32593 39753
rect 32593 39701 32595 39753
rect 32539 39699 32595 39701
rect 32750 39753 32806 39755
rect 32750 39701 32752 39753
rect 32752 39701 32804 39753
rect 32804 39701 32806 39753
rect 32750 39699 32806 39701
rect 33055 39266 33111 39322
rect 33235 39266 33291 39322
rect 33817 39259 33873 39315
rect 33997 39259 34053 39315
rect 34282 38799 34338 38855
rect 34493 38799 34549 38855
rect 34705 38853 34761 38855
rect 34916 38853 34972 38855
rect 34705 38801 34755 38853
rect 34755 38801 34761 38853
rect 34916 38801 34935 38853
rect 34935 38801 34972 38853
rect 34705 38799 34761 38801
rect 34916 38799 34972 38801
rect 33055 38332 33111 38388
rect 33235 38332 33291 38388
rect 33817 38339 33873 38395
rect 33997 38339 34053 38395
rect 30852 37953 30908 37955
rect 30852 37901 30854 37953
rect 30854 37901 30906 37953
rect 30906 37901 30908 37953
rect 30852 37899 30908 37901
rect 31063 37953 31119 37955
rect 31063 37901 31065 37953
rect 31065 37901 31117 37953
rect 31117 37901 31119 37953
rect 31063 37899 31119 37901
rect 31274 37953 31330 37955
rect 31274 37901 31276 37953
rect 31276 37901 31328 37953
rect 31328 37901 31330 37953
rect 31274 37899 31330 37901
rect 31484 37953 31540 37955
rect 31484 37901 31486 37953
rect 31486 37901 31538 37953
rect 31538 37901 31540 37953
rect 31484 37899 31540 37901
rect 31695 37953 31751 37955
rect 31695 37901 31697 37953
rect 31697 37901 31749 37953
rect 31749 37901 31751 37953
rect 31695 37899 31751 37901
rect 31907 37953 31963 37955
rect 31907 37901 31909 37953
rect 31909 37901 31961 37953
rect 31961 37901 31963 37953
rect 31907 37899 31963 37901
rect 32118 37953 32174 37955
rect 32118 37901 32120 37953
rect 32120 37901 32172 37953
rect 32172 37901 32174 37953
rect 32118 37899 32174 37901
rect 32328 37953 32384 37955
rect 32328 37901 32330 37953
rect 32330 37901 32382 37953
rect 32382 37901 32384 37953
rect 32328 37899 32384 37901
rect 32539 37953 32595 37955
rect 32539 37901 32541 37953
rect 32541 37901 32593 37953
rect 32593 37901 32595 37953
rect 32539 37899 32595 37901
rect 32750 37953 32806 37955
rect 32750 37901 32752 37953
rect 32752 37901 32804 37953
rect 32804 37901 32806 37953
rect 32750 37899 32806 37901
rect 33055 37466 33111 37522
rect 33235 37466 33291 37522
rect 33817 37459 33873 37515
rect 33997 37459 34053 37515
rect 34282 36999 34338 37055
rect 34493 36999 34549 37055
rect 34705 37053 34761 37055
rect 34916 37053 34972 37055
rect 34705 37001 34755 37053
rect 34755 37001 34761 37053
rect 34916 37001 34935 37053
rect 34935 37001 34972 37053
rect 34705 36999 34761 37001
rect 34916 36999 34972 37001
rect 33055 36532 33111 36588
rect 33235 36532 33291 36588
rect 33817 36539 33873 36595
rect 33997 36539 34053 36595
rect 30852 36153 30908 36155
rect 30852 36101 30854 36153
rect 30854 36101 30906 36153
rect 30906 36101 30908 36153
rect 30852 36099 30908 36101
rect 31063 36153 31119 36155
rect 31063 36101 31065 36153
rect 31065 36101 31117 36153
rect 31117 36101 31119 36153
rect 31063 36099 31119 36101
rect 31274 36153 31330 36155
rect 31274 36101 31276 36153
rect 31276 36101 31328 36153
rect 31328 36101 31330 36153
rect 31274 36099 31330 36101
rect 31484 36153 31540 36155
rect 31484 36101 31486 36153
rect 31486 36101 31538 36153
rect 31538 36101 31540 36153
rect 31484 36099 31540 36101
rect 31695 36153 31751 36155
rect 31695 36101 31697 36153
rect 31697 36101 31749 36153
rect 31749 36101 31751 36153
rect 31695 36099 31751 36101
rect 31907 36153 31963 36155
rect 31907 36101 31909 36153
rect 31909 36101 31961 36153
rect 31961 36101 31963 36153
rect 31907 36099 31963 36101
rect 32118 36153 32174 36155
rect 32118 36101 32120 36153
rect 32120 36101 32172 36153
rect 32172 36101 32174 36153
rect 32118 36099 32174 36101
rect 32328 36153 32384 36155
rect 32328 36101 32330 36153
rect 32330 36101 32382 36153
rect 32382 36101 32384 36153
rect 32328 36099 32384 36101
rect 32539 36153 32595 36155
rect 32539 36101 32541 36153
rect 32541 36101 32593 36153
rect 32593 36101 32595 36153
rect 32539 36099 32595 36101
rect 32750 36153 32806 36155
rect 32750 36101 32752 36153
rect 32752 36101 32804 36153
rect 32804 36101 32806 36153
rect 32750 36099 32806 36101
rect 35218 64901 35220 64953
rect 35220 64901 35272 64953
rect 35272 64901 35274 64953
rect 35218 64899 35274 64901
rect 35428 64953 35484 64955
rect 35428 64901 35430 64953
rect 35430 64901 35482 64953
rect 35482 64901 35484 64953
rect 35428 64899 35484 64901
rect 35639 64953 35695 64955
rect 35639 64901 35641 64953
rect 35641 64901 35693 64953
rect 35693 64901 35695 64953
rect 35639 64899 35695 64901
rect 35851 64953 35907 64955
rect 35851 64901 35853 64953
rect 35853 64901 35905 64953
rect 35905 64901 35907 64953
rect 35851 64899 35907 64901
rect 36062 64953 36118 64955
rect 36062 64901 36064 64953
rect 36064 64901 36116 64953
rect 36116 64901 36118 64953
rect 36062 64899 36118 64901
rect 36272 64953 36328 64955
rect 36272 64901 36274 64953
rect 36274 64901 36326 64953
rect 36326 64901 36328 64953
rect 36272 64899 36328 64901
rect 36899 65316 36955 65372
rect 37110 65316 37166 65372
rect 37321 65316 37377 65372
rect 37532 65316 37588 65372
rect 40250 65806 40252 65855
rect 40252 65806 40304 65855
rect 40304 65806 40306 65855
rect 40250 65799 40306 65806
rect 40430 65806 40432 65855
rect 40432 65806 40484 65855
rect 40484 65806 40486 65855
rect 40430 65799 40486 65806
rect 41008 65370 41064 65372
rect 41008 65318 41010 65370
rect 41010 65318 41062 65370
rect 41062 65318 41064 65370
rect 41008 65316 41064 65318
rect 41219 65370 41275 65372
rect 41219 65318 41221 65370
rect 41221 65318 41273 65370
rect 41273 65318 41275 65370
rect 41219 65316 41275 65318
rect 41430 65370 41486 65372
rect 41430 65318 41432 65370
rect 41432 65318 41484 65370
rect 41484 65318 41486 65370
rect 41430 65316 41486 65318
rect 41641 65370 41697 65372
rect 41641 65318 41643 65370
rect 41643 65318 41695 65370
rect 41695 65318 41697 65370
rect 41641 65316 41697 65318
rect 41852 65370 41908 65372
rect 41852 65318 41854 65370
rect 41854 65318 41906 65370
rect 41906 65318 41908 65370
rect 41852 65316 41908 65318
rect 42062 65370 42118 65372
rect 42062 65318 42064 65370
rect 42064 65318 42116 65370
rect 42116 65318 42118 65370
rect 42062 65316 42118 65318
rect 42708 65309 42764 65365
rect 42919 65309 42975 65365
rect 43130 65309 43186 65365
rect 36676 64507 36732 64563
rect 39050 64953 39106 64955
rect 36676 63491 36732 63547
rect 37889 64276 37945 64332
rect 38069 64276 38125 64332
rect 38328 63999 38384 64055
rect 38539 63999 38595 64055
rect 38750 63999 38806 64055
rect 35218 63153 35274 63155
rect 35218 63101 35220 63153
rect 35220 63101 35272 63153
rect 35272 63101 35274 63153
rect 35218 63099 35274 63101
rect 35428 63153 35484 63155
rect 35428 63101 35430 63153
rect 35430 63101 35482 63153
rect 35482 63101 35484 63153
rect 35428 63099 35484 63101
rect 35639 63153 35695 63155
rect 35639 63101 35641 63153
rect 35641 63101 35693 63153
rect 35693 63101 35695 63153
rect 35639 63099 35695 63101
rect 35851 63153 35907 63155
rect 35851 63101 35853 63153
rect 35853 63101 35905 63153
rect 35905 63101 35907 63153
rect 35851 63099 35907 63101
rect 36062 63153 36118 63155
rect 36062 63101 36064 63153
rect 36064 63101 36116 63153
rect 36116 63101 36118 63153
rect 36062 63099 36118 63101
rect 36272 63153 36328 63155
rect 36272 63101 36274 63153
rect 36274 63101 36326 63153
rect 36326 63101 36328 63153
rect 36272 63099 36328 63101
rect 36676 62707 36732 62763
rect 37889 63722 37945 63778
rect 38069 63722 38125 63778
rect 36676 61691 36732 61747
rect 37889 62476 37945 62532
rect 38069 62476 38125 62532
rect 38328 62199 38384 62255
rect 38539 62199 38595 62255
rect 38750 62199 38806 62255
rect 35218 61353 35274 61355
rect 35218 61301 35220 61353
rect 35220 61301 35272 61353
rect 35272 61301 35274 61353
rect 35218 61299 35274 61301
rect 35428 61353 35484 61355
rect 35428 61301 35430 61353
rect 35430 61301 35482 61353
rect 35482 61301 35484 61353
rect 35428 61299 35484 61301
rect 35639 61353 35695 61355
rect 35639 61301 35641 61353
rect 35641 61301 35693 61353
rect 35693 61301 35695 61353
rect 35639 61299 35695 61301
rect 35851 61353 35907 61355
rect 35851 61301 35853 61353
rect 35853 61301 35905 61353
rect 35905 61301 35907 61353
rect 35851 61299 35907 61301
rect 36062 61353 36118 61355
rect 36062 61301 36064 61353
rect 36064 61301 36116 61353
rect 36116 61301 36118 61353
rect 36062 61299 36118 61301
rect 36272 61353 36328 61355
rect 36272 61301 36274 61353
rect 36274 61301 36326 61353
rect 36326 61301 36328 61353
rect 36272 61299 36328 61301
rect 36676 60907 36732 60963
rect 37889 61922 37945 61978
rect 38069 61922 38125 61978
rect 36676 59891 36732 59947
rect 37889 60676 37945 60732
rect 38069 60676 38125 60732
rect 38328 60399 38384 60455
rect 38539 60399 38595 60455
rect 38750 60399 38806 60455
rect 35218 59553 35274 59555
rect 35218 59501 35220 59553
rect 35220 59501 35272 59553
rect 35272 59501 35274 59553
rect 35218 59499 35274 59501
rect 35428 59553 35484 59555
rect 35428 59501 35430 59553
rect 35430 59501 35482 59553
rect 35482 59501 35484 59553
rect 35428 59499 35484 59501
rect 35639 59553 35695 59555
rect 35639 59501 35641 59553
rect 35641 59501 35693 59553
rect 35693 59501 35695 59553
rect 35639 59499 35695 59501
rect 35851 59553 35907 59555
rect 35851 59501 35853 59553
rect 35853 59501 35905 59553
rect 35905 59501 35907 59553
rect 35851 59499 35907 59501
rect 36062 59553 36118 59555
rect 36062 59501 36064 59553
rect 36064 59501 36116 59553
rect 36116 59501 36118 59553
rect 36062 59499 36118 59501
rect 36272 59553 36328 59555
rect 36272 59501 36274 59553
rect 36274 59501 36326 59553
rect 36326 59501 36328 59553
rect 36272 59499 36328 59501
rect 36676 59107 36732 59163
rect 37889 60122 37945 60178
rect 38069 60122 38125 60178
rect 36676 58091 36732 58147
rect 37889 58876 37945 58932
rect 38069 58876 38125 58932
rect 38328 58599 38384 58655
rect 38539 58599 38595 58655
rect 38750 58599 38806 58655
rect 35218 57753 35274 57755
rect 35218 57701 35220 57753
rect 35220 57701 35272 57753
rect 35272 57701 35274 57753
rect 35218 57699 35274 57701
rect 35428 57753 35484 57755
rect 35428 57701 35430 57753
rect 35430 57701 35482 57753
rect 35482 57701 35484 57753
rect 35428 57699 35484 57701
rect 35639 57753 35695 57755
rect 35639 57701 35641 57753
rect 35641 57701 35693 57753
rect 35693 57701 35695 57753
rect 35639 57699 35695 57701
rect 35851 57753 35907 57755
rect 35851 57701 35853 57753
rect 35853 57701 35905 57753
rect 35905 57701 35907 57753
rect 35851 57699 35907 57701
rect 36062 57753 36118 57755
rect 36062 57701 36064 57753
rect 36064 57701 36116 57753
rect 36116 57701 36118 57753
rect 36062 57699 36118 57701
rect 36272 57753 36328 57755
rect 36272 57701 36274 57753
rect 36274 57701 36326 57753
rect 36326 57701 36328 57753
rect 36272 57699 36328 57701
rect 36676 57307 36732 57363
rect 37889 58322 37945 58378
rect 38069 58322 38125 58378
rect 36676 56291 36732 56347
rect 37889 57076 37945 57132
rect 38069 57076 38125 57132
rect 38328 56799 38384 56855
rect 38539 56799 38595 56855
rect 38750 56799 38806 56855
rect 35218 55953 35274 55955
rect 35218 55901 35220 55953
rect 35220 55901 35272 55953
rect 35272 55901 35274 55953
rect 35218 55899 35274 55901
rect 35428 55953 35484 55955
rect 35428 55901 35430 55953
rect 35430 55901 35482 55953
rect 35482 55901 35484 55953
rect 35428 55899 35484 55901
rect 35639 55953 35695 55955
rect 35639 55901 35641 55953
rect 35641 55901 35693 55953
rect 35693 55901 35695 55953
rect 35639 55899 35695 55901
rect 35851 55953 35907 55955
rect 35851 55901 35853 55953
rect 35853 55901 35905 55953
rect 35905 55901 35907 55953
rect 35851 55899 35907 55901
rect 36062 55953 36118 55955
rect 36062 55901 36064 55953
rect 36064 55901 36116 55953
rect 36116 55901 36118 55953
rect 36062 55899 36118 55901
rect 36272 55953 36328 55955
rect 36272 55901 36274 55953
rect 36274 55901 36326 55953
rect 36326 55901 36328 55953
rect 36272 55899 36328 55901
rect 36676 55507 36732 55563
rect 37889 56522 37945 56578
rect 38069 56522 38125 56578
rect 36676 54491 36732 54547
rect 37889 55276 37945 55332
rect 38069 55276 38125 55332
rect 38328 54999 38384 55055
rect 38539 54999 38595 55055
rect 38750 54999 38806 55055
rect 35218 54153 35274 54155
rect 35218 54101 35220 54153
rect 35220 54101 35272 54153
rect 35272 54101 35274 54153
rect 35218 54099 35274 54101
rect 35428 54153 35484 54155
rect 35428 54101 35430 54153
rect 35430 54101 35482 54153
rect 35482 54101 35484 54153
rect 35428 54099 35484 54101
rect 35639 54153 35695 54155
rect 35639 54101 35641 54153
rect 35641 54101 35693 54153
rect 35693 54101 35695 54153
rect 35639 54099 35695 54101
rect 35851 54153 35907 54155
rect 35851 54101 35853 54153
rect 35853 54101 35905 54153
rect 35905 54101 35907 54153
rect 35851 54099 35907 54101
rect 36062 54153 36118 54155
rect 36062 54101 36064 54153
rect 36064 54101 36116 54153
rect 36116 54101 36118 54153
rect 36062 54099 36118 54101
rect 36272 54153 36328 54155
rect 36272 54101 36274 54153
rect 36274 54101 36326 54153
rect 36326 54101 36328 54153
rect 36272 54099 36328 54101
rect 36676 53707 36732 53763
rect 37889 54722 37945 54778
rect 38069 54722 38125 54778
rect 36676 52691 36732 52747
rect 37889 53476 37945 53532
rect 38069 53476 38125 53532
rect 38328 53199 38384 53255
rect 38539 53199 38595 53255
rect 38750 53199 38806 53255
rect 35218 52353 35274 52355
rect 35218 52301 35220 52353
rect 35220 52301 35272 52353
rect 35272 52301 35274 52353
rect 35218 52299 35274 52301
rect 35428 52353 35484 52355
rect 35428 52301 35430 52353
rect 35430 52301 35482 52353
rect 35482 52301 35484 52353
rect 35428 52299 35484 52301
rect 35639 52353 35695 52355
rect 35639 52301 35641 52353
rect 35641 52301 35693 52353
rect 35693 52301 35695 52353
rect 35639 52299 35695 52301
rect 35851 52353 35907 52355
rect 35851 52301 35853 52353
rect 35853 52301 35905 52353
rect 35905 52301 35907 52353
rect 35851 52299 35907 52301
rect 36062 52353 36118 52355
rect 36062 52301 36064 52353
rect 36064 52301 36116 52353
rect 36116 52301 36118 52353
rect 36062 52299 36118 52301
rect 36272 52353 36328 52355
rect 36272 52301 36274 52353
rect 36274 52301 36326 52353
rect 36326 52301 36328 52353
rect 36272 52299 36328 52301
rect 36676 51907 36732 51963
rect 37889 52922 37945 52978
rect 38069 52922 38125 52978
rect 36676 50891 36732 50947
rect 37889 51676 37945 51732
rect 38069 51676 38125 51732
rect 38328 51399 38384 51455
rect 38539 51399 38595 51455
rect 38750 51399 38806 51455
rect 35218 50553 35274 50555
rect 35218 50501 35220 50553
rect 35220 50501 35272 50553
rect 35272 50501 35274 50553
rect 35218 50499 35274 50501
rect 35428 50553 35484 50555
rect 35428 50501 35430 50553
rect 35430 50501 35482 50553
rect 35482 50501 35484 50553
rect 35428 50499 35484 50501
rect 35639 50553 35695 50555
rect 35639 50501 35641 50553
rect 35641 50501 35693 50553
rect 35693 50501 35695 50553
rect 35639 50499 35695 50501
rect 35851 50553 35907 50555
rect 35851 50501 35853 50553
rect 35853 50501 35905 50553
rect 35905 50501 35907 50553
rect 35851 50499 35907 50501
rect 36062 50553 36118 50555
rect 36062 50501 36064 50553
rect 36064 50501 36116 50553
rect 36116 50501 36118 50553
rect 36062 50499 36118 50501
rect 36272 50553 36328 50555
rect 36272 50501 36274 50553
rect 36274 50501 36326 50553
rect 36326 50501 36328 50553
rect 36272 50499 36328 50501
rect 36676 50107 36732 50163
rect 37889 51122 37945 51178
rect 38069 51122 38125 51178
rect 36676 49091 36732 49147
rect 37889 49876 37945 49932
rect 38069 49876 38125 49932
rect 38328 49599 38384 49655
rect 38539 49599 38595 49655
rect 38750 49599 38806 49655
rect 35218 48753 35274 48755
rect 35218 48701 35220 48753
rect 35220 48701 35272 48753
rect 35272 48701 35274 48753
rect 35218 48699 35274 48701
rect 35428 48753 35484 48755
rect 35428 48701 35430 48753
rect 35430 48701 35482 48753
rect 35482 48701 35484 48753
rect 35428 48699 35484 48701
rect 35639 48753 35695 48755
rect 35639 48701 35641 48753
rect 35641 48701 35693 48753
rect 35693 48701 35695 48753
rect 35639 48699 35695 48701
rect 35851 48753 35907 48755
rect 35851 48701 35853 48753
rect 35853 48701 35905 48753
rect 35905 48701 35907 48753
rect 35851 48699 35907 48701
rect 36062 48753 36118 48755
rect 36062 48701 36064 48753
rect 36064 48701 36116 48753
rect 36116 48701 36118 48753
rect 36062 48699 36118 48701
rect 36272 48753 36328 48755
rect 36272 48701 36274 48753
rect 36274 48701 36326 48753
rect 36326 48701 36328 48753
rect 36272 48699 36328 48701
rect 36676 48307 36732 48363
rect 37889 49322 37945 49378
rect 38069 49322 38125 49378
rect 36676 47291 36732 47347
rect 37889 48076 37945 48132
rect 38069 48076 38125 48132
rect 38328 47799 38384 47855
rect 38539 47799 38595 47855
rect 38750 47799 38806 47855
rect 35218 46953 35274 46955
rect 35218 46901 35220 46953
rect 35220 46901 35272 46953
rect 35272 46901 35274 46953
rect 35218 46899 35274 46901
rect 35428 46953 35484 46955
rect 35428 46901 35430 46953
rect 35430 46901 35482 46953
rect 35482 46901 35484 46953
rect 35428 46899 35484 46901
rect 35639 46953 35695 46955
rect 35639 46901 35641 46953
rect 35641 46901 35693 46953
rect 35693 46901 35695 46953
rect 35639 46899 35695 46901
rect 35851 46953 35907 46955
rect 35851 46901 35853 46953
rect 35853 46901 35905 46953
rect 35905 46901 35907 46953
rect 35851 46899 35907 46901
rect 36062 46953 36118 46955
rect 36062 46901 36064 46953
rect 36064 46901 36116 46953
rect 36116 46901 36118 46953
rect 36062 46899 36118 46901
rect 36272 46953 36328 46955
rect 36272 46901 36274 46953
rect 36274 46901 36326 46953
rect 36326 46901 36328 46953
rect 36272 46899 36328 46901
rect 36676 46507 36732 46563
rect 37889 47522 37945 47578
rect 38069 47522 38125 47578
rect 36676 45491 36732 45547
rect 37889 46276 37945 46332
rect 38069 46276 38125 46332
rect 38328 45999 38384 46055
rect 38539 45999 38595 46055
rect 38750 45999 38806 46055
rect 35218 45153 35274 45155
rect 35218 45101 35220 45153
rect 35220 45101 35272 45153
rect 35272 45101 35274 45153
rect 35218 45099 35274 45101
rect 35428 45153 35484 45155
rect 35428 45101 35430 45153
rect 35430 45101 35482 45153
rect 35482 45101 35484 45153
rect 35428 45099 35484 45101
rect 35639 45153 35695 45155
rect 35639 45101 35641 45153
rect 35641 45101 35693 45153
rect 35693 45101 35695 45153
rect 35639 45099 35695 45101
rect 35851 45153 35907 45155
rect 35851 45101 35853 45153
rect 35853 45101 35905 45153
rect 35905 45101 35907 45153
rect 35851 45099 35907 45101
rect 36062 45153 36118 45155
rect 36062 45101 36064 45153
rect 36064 45101 36116 45153
rect 36116 45101 36118 45153
rect 36062 45099 36118 45101
rect 36272 45153 36328 45155
rect 36272 45101 36274 45153
rect 36274 45101 36326 45153
rect 36326 45101 36328 45153
rect 36272 45099 36328 45101
rect 36676 44707 36732 44763
rect 37889 45722 37945 45778
rect 38069 45722 38125 45778
rect 36676 43691 36732 43747
rect 37889 44476 37945 44532
rect 38069 44476 38125 44532
rect 38328 44199 38384 44255
rect 38539 44199 38595 44255
rect 38750 44199 38806 44255
rect 35218 43353 35274 43355
rect 35218 43301 35220 43353
rect 35220 43301 35272 43353
rect 35272 43301 35274 43353
rect 35218 43299 35274 43301
rect 35428 43353 35484 43355
rect 35428 43301 35430 43353
rect 35430 43301 35482 43353
rect 35482 43301 35484 43353
rect 35428 43299 35484 43301
rect 35639 43353 35695 43355
rect 35639 43301 35641 43353
rect 35641 43301 35693 43353
rect 35693 43301 35695 43353
rect 35639 43299 35695 43301
rect 35851 43353 35907 43355
rect 35851 43301 35853 43353
rect 35853 43301 35905 43353
rect 35905 43301 35907 43353
rect 35851 43299 35907 43301
rect 36062 43353 36118 43355
rect 36062 43301 36064 43353
rect 36064 43301 36116 43353
rect 36116 43301 36118 43353
rect 36062 43299 36118 43301
rect 36272 43353 36328 43355
rect 36272 43301 36274 43353
rect 36274 43301 36326 43353
rect 36326 43301 36328 43353
rect 36272 43299 36328 43301
rect 36676 42907 36732 42963
rect 37889 43922 37945 43978
rect 38069 43922 38125 43978
rect 36676 41891 36732 41947
rect 37889 42676 37945 42732
rect 38069 42676 38125 42732
rect 38328 42399 38384 42455
rect 38539 42399 38595 42455
rect 38750 42399 38806 42455
rect 35218 41553 35274 41555
rect 35218 41501 35220 41553
rect 35220 41501 35272 41553
rect 35272 41501 35274 41553
rect 35218 41499 35274 41501
rect 35428 41553 35484 41555
rect 35428 41501 35430 41553
rect 35430 41501 35482 41553
rect 35482 41501 35484 41553
rect 35428 41499 35484 41501
rect 35639 41553 35695 41555
rect 35639 41501 35641 41553
rect 35641 41501 35693 41553
rect 35693 41501 35695 41553
rect 35639 41499 35695 41501
rect 35851 41553 35907 41555
rect 35851 41501 35853 41553
rect 35853 41501 35905 41553
rect 35905 41501 35907 41553
rect 35851 41499 35907 41501
rect 36062 41553 36118 41555
rect 36062 41501 36064 41553
rect 36064 41501 36116 41553
rect 36116 41501 36118 41553
rect 36062 41499 36118 41501
rect 36272 41553 36328 41555
rect 36272 41501 36274 41553
rect 36274 41501 36326 41553
rect 36326 41501 36328 41553
rect 36272 41499 36328 41501
rect 36676 41107 36732 41163
rect 37889 42122 37945 42178
rect 38069 42122 38125 42178
rect 36676 40091 36732 40147
rect 37889 40876 37945 40932
rect 38069 40876 38125 40932
rect 38328 40599 38384 40655
rect 38539 40599 38595 40655
rect 38750 40599 38806 40655
rect 35218 39753 35274 39755
rect 35218 39701 35220 39753
rect 35220 39701 35272 39753
rect 35272 39701 35274 39753
rect 35218 39699 35274 39701
rect 35428 39753 35484 39755
rect 35428 39701 35430 39753
rect 35430 39701 35482 39753
rect 35482 39701 35484 39753
rect 35428 39699 35484 39701
rect 35639 39753 35695 39755
rect 35639 39701 35641 39753
rect 35641 39701 35693 39753
rect 35693 39701 35695 39753
rect 35639 39699 35695 39701
rect 35851 39753 35907 39755
rect 35851 39701 35853 39753
rect 35853 39701 35905 39753
rect 35905 39701 35907 39753
rect 35851 39699 35907 39701
rect 36062 39753 36118 39755
rect 36062 39701 36064 39753
rect 36064 39701 36116 39753
rect 36116 39701 36118 39753
rect 36062 39699 36118 39701
rect 36272 39753 36328 39755
rect 36272 39701 36274 39753
rect 36274 39701 36326 39753
rect 36326 39701 36328 39753
rect 36272 39699 36328 39701
rect 36676 39307 36732 39363
rect 37889 40322 37945 40378
rect 38069 40322 38125 40378
rect 36676 38291 36732 38347
rect 37889 39076 37945 39132
rect 38069 39076 38125 39132
rect 38328 38799 38384 38855
rect 38539 38799 38595 38855
rect 38750 38799 38806 38855
rect 35218 37953 35274 37955
rect 35218 37901 35220 37953
rect 35220 37901 35272 37953
rect 35272 37901 35274 37953
rect 35218 37899 35274 37901
rect 35428 37953 35484 37955
rect 35428 37901 35430 37953
rect 35430 37901 35482 37953
rect 35482 37901 35484 37953
rect 35428 37899 35484 37901
rect 35639 37953 35695 37955
rect 35639 37901 35641 37953
rect 35641 37901 35693 37953
rect 35693 37901 35695 37953
rect 35639 37899 35695 37901
rect 35851 37953 35907 37955
rect 35851 37901 35853 37953
rect 35853 37901 35905 37953
rect 35905 37901 35907 37953
rect 35851 37899 35907 37901
rect 36062 37953 36118 37955
rect 36062 37901 36064 37953
rect 36064 37901 36116 37953
rect 36116 37901 36118 37953
rect 36062 37899 36118 37901
rect 36272 37953 36328 37955
rect 36272 37901 36274 37953
rect 36274 37901 36326 37953
rect 36326 37901 36328 37953
rect 36272 37899 36328 37901
rect 36676 37507 36732 37563
rect 37889 38522 37945 38578
rect 38069 38522 38125 38578
rect 37889 37276 37945 37332
rect 38069 37276 38125 37332
rect 38328 36999 38384 37055
rect 38539 36999 38595 37055
rect 38750 36999 38806 37055
rect 36676 36491 36732 36547
rect 35218 36153 35274 36155
rect 35218 36101 35220 36153
rect 35220 36101 35272 36153
rect 35272 36101 35274 36153
rect 35218 36099 35274 36101
rect 35428 36153 35484 36155
rect 35428 36101 35430 36153
rect 35430 36101 35482 36153
rect 35482 36101 35484 36153
rect 35428 36099 35484 36101
rect 35639 36153 35695 36155
rect 35639 36101 35641 36153
rect 35641 36101 35693 36153
rect 35693 36101 35695 36153
rect 35639 36099 35695 36101
rect 35851 36153 35907 36155
rect 35851 36101 35853 36153
rect 35853 36101 35905 36153
rect 35905 36101 35907 36153
rect 35851 36099 35907 36101
rect 36062 36153 36118 36155
rect 36062 36101 36064 36153
rect 36064 36101 36116 36153
rect 36116 36101 36118 36153
rect 36062 36099 36118 36101
rect 36272 36153 36328 36155
rect 36272 36101 36274 36153
rect 36274 36101 36326 36153
rect 36326 36101 36328 36153
rect 36272 36099 36328 36101
rect 37889 36722 37945 36778
rect 38069 36722 38125 36778
rect 39050 64901 39052 64953
rect 39052 64901 39104 64953
rect 39104 64901 39106 64953
rect 39050 64899 39106 64901
rect 39230 64953 39286 64955
rect 39230 64901 39232 64953
rect 39232 64901 39284 64953
rect 39284 64901 39286 64953
rect 39230 64899 39286 64901
rect 39773 64276 39829 64332
rect 39992 64507 40048 64563
rect 40777 64899 40833 64955
rect 40988 64899 41044 64955
rect 41199 64899 41255 64955
rect 40251 63999 40307 64055
rect 40431 63999 40487 64055
rect 39773 63722 39829 63778
rect 39992 63491 40048 63547
rect 39050 63153 39106 63155
rect 39050 63101 39052 63153
rect 39052 63101 39104 63153
rect 39104 63101 39106 63153
rect 39050 63099 39106 63101
rect 39230 63153 39286 63155
rect 39230 63101 39232 63153
rect 39232 63101 39284 63153
rect 39284 63101 39286 63153
rect 39230 63099 39286 63101
rect 39773 62476 39829 62532
rect 39992 62707 40048 62763
rect 40251 62199 40307 62255
rect 40431 62199 40487 62255
rect 39773 61922 39829 61978
rect 39992 61691 40048 61747
rect 39050 61353 39106 61355
rect 39050 61301 39052 61353
rect 39052 61301 39104 61353
rect 39104 61301 39106 61353
rect 39050 61299 39106 61301
rect 39230 61353 39286 61355
rect 39230 61301 39232 61353
rect 39232 61301 39284 61353
rect 39284 61301 39286 61353
rect 39230 61299 39286 61301
rect 39773 60676 39829 60732
rect 39992 60907 40048 60963
rect 40251 60399 40307 60455
rect 40431 60399 40487 60455
rect 39773 60122 39829 60178
rect 39992 59891 40048 59947
rect 39050 59553 39106 59555
rect 39050 59501 39052 59553
rect 39052 59501 39104 59553
rect 39104 59501 39106 59553
rect 39050 59499 39106 59501
rect 39230 59553 39286 59555
rect 39230 59501 39232 59553
rect 39232 59501 39284 59553
rect 39284 59501 39286 59553
rect 39230 59499 39286 59501
rect 39773 58876 39829 58932
rect 39992 59107 40048 59163
rect 40251 58599 40307 58655
rect 40431 58599 40487 58655
rect 39773 58322 39829 58378
rect 39992 58091 40048 58147
rect 39050 57753 39106 57755
rect 39050 57701 39052 57753
rect 39052 57701 39104 57753
rect 39104 57701 39106 57753
rect 39050 57699 39106 57701
rect 39230 57753 39286 57755
rect 39230 57701 39232 57753
rect 39232 57701 39284 57753
rect 39284 57701 39286 57753
rect 39230 57699 39286 57701
rect 39773 57076 39829 57132
rect 39992 57307 40048 57363
rect 40251 56799 40307 56855
rect 40431 56799 40487 56855
rect 39773 56522 39829 56578
rect 39992 56291 40048 56347
rect 39050 55953 39106 55955
rect 39050 55901 39052 55953
rect 39052 55901 39104 55953
rect 39104 55901 39106 55953
rect 39050 55899 39106 55901
rect 39230 55953 39286 55955
rect 39230 55901 39232 55953
rect 39232 55901 39284 55953
rect 39284 55901 39286 55953
rect 39230 55899 39286 55901
rect 39773 55276 39829 55332
rect 39992 55507 40048 55563
rect 40251 54999 40307 55055
rect 40431 54999 40487 55055
rect 39773 54722 39829 54778
rect 39992 54491 40048 54547
rect 39050 54153 39106 54155
rect 39050 54101 39052 54153
rect 39052 54101 39104 54153
rect 39104 54101 39106 54153
rect 39050 54099 39106 54101
rect 39230 54153 39286 54155
rect 39230 54101 39232 54153
rect 39232 54101 39284 54153
rect 39284 54101 39286 54153
rect 39230 54099 39286 54101
rect 39773 53476 39829 53532
rect 39992 53707 40048 53763
rect 40251 53199 40307 53255
rect 40431 53199 40487 53255
rect 39773 52922 39829 52978
rect 39992 52691 40048 52747
rect 39050 52353 39106 52355
rect 39050 52301 39052 52353
rect 39052 52301 39104 52353
rect 39104 52301 39106 52353
rect 39050 52299 39106 52301
rect 39230 52353 39286 52355
rect 39230 52301 39232 52353
rect 39232 52301 39284 52353
rect 39284 52301 39286 52353
rect 39230 52299 39286 52301
rect 39773 51676 39829 51732
rect 39992 51907 40048 51963
rect 40251 51399 40307 51455
rect 40431 51399 40487 51455
rect 39773 51122 39829 51178
rect 39992 50891 40048 50947
rect 39050 50553 39106 50555
rect 39050 50501 39052 50553
rect 39052 50501 39104 50553
rect 39104 50501 39106 50553
rect 39050 50499 39106 50501
rect 39230 50553 39286 50555
rect 39230 50501 39232 50553
rect 39232 50501 39284 50553
rect 39284 50501 39286 50553
rect 39230 50499 39286 50501
rect 39773 49876 39829 49932
rect 39992 50107 40048 50163
rect 40251 49599 40307 49655
rect 40431 49599 40487 49655
rect 39773 49322 39829 49378
rect 39992 49091 40048 49147
rect 39050 48753 39106 48755
rect 39050 48701 39052 48753
rect 39052 48701 39104 48753
rect 39104 48701 39106 48753
rect 39050 48699 39106 48701
rect 39230 48753 39286 48755
rect 39230 48701 39232 48753
rect 39232 48701 39284 48753
rect 39284 48701 39286 48753
rect 39230 48699 39286 48701
rect 39773 48076 39829 48132
rect 39992 48307 40048 48363
rect 40251 47799 40307 47855
rect 40431 47799 40487 47855
rect 39773 47522 39829 47578
rect 39992 47291 40048 47347
rect 39050 46953 39106 46955
rect 39050 46901 39052 46953
rect 39052 46901 39104 46953
rect 39104 46901 39106 46953
rect 39050 46899 39106 46901
rect 39230 46953 39286 46955
rect 39230 46901 39232 46953
rect 39232 46901 39284 46953
rect 39284 46901 39286 46953
rect 39230 46899 39286 46901
rect 39773 46276 39829 46332
rect 39992 46507 40048 46563
rect 40251 45999 40307 46055
rect 40431 45999 40487 46055
rect 39773 45722 39829 45778
rect 39992 45491 40048 45547
rect 39050 45153 39106 45155
rect 39050 45101 39052 45153
rect 39052 45101 39104 45153
rect 39104 45101 39106 45153
rect 39050 45099 39106 45101
rect 39230 45153 39286 45155
rect 39230 45101 39232 45153
rect 39232 45101 39284 45153
rect 39284 45101 39286 45153
rect 39230 45099 39286 45101
rect 39773 44476 39829 44532
rect 39992 44707 40048 44763
rect 40251 44199 40307 44255
rect 40431 44199 40487 44255
rect 39773 43922 39829 43978
rect 39992 43691 40048 43747
rect 39050 43353 39106 43355
rect 39050 43301 39052 43353
rect 39052 43301 39104 43353
rect 39104 43301 39106 43353
rect 39050 43299 39106 43301
rect 39230 43353 39286 43355
rect 39230 43301 39232 43353
rect 39232 43301 39284 43353
rect 39284 43301 39286 43353
rect 39230 43299 39286 43301
rect 39773 42676 39829 42732
rect 39992 42907 40048 42963
rect 40251 42399 40307 42455
rect 40431 42399 40487 42455
rect 39773 42122 39829 42178
rect 39992 41891 40048 41947
rect 39050 41553 39106 41555
rect 39050 41501 39052 41553
rect 39052 41501 39104 41553
rect 39104 41501 39106 41553
rect 39050 41499 39106 41501
rect 39230 41553 39286 41555
rect 39230 41501 39232 41553
rect 39232 41501 39284 41553
rect 39284 41501 39286 41553
rect 39230 41499 39286 41501
rect 39773 40876 39829 40932
rect 39992 41107 40048 41163
rect 40251 40599 40307 40655
rect 40431 40599 40487 40655
rect 39773 40322 39829 40378
rect 39992 40091 40048 40147
rect 39050 39753 39106 39755
rect 39050 39701 39052 39753
rect 39052 39701 39104 39753
rect 39104 39701 39106 39753
rect 39050 39699 39106 39701
rect 39230 39753 39286 39755
rect 39230 39701 39232 39753
rect 39232 39701 39284 39753
rect 39284 39701 39286 39753
rect 39230 39699 39286 39701
rect 39773 39076 39829 39132
rect 39992 39307 40048 39363
rect 40251 38799 40307 38855
rect 40431 38799 40487 38855
rect 39773 38522 39829 38578
rect 39992 38291 40048 38347
rect 39050 37953 39106 37955
rect 39050 37901 39052 37953
rect 39052 37901 39104 37953
rect 39104 37901 39106 37953
rect 39050 37899 39106 37901
rect 39230 37953 39286 37955
rect 39230 37901 39232 37953
rect 39232 37901 39284 37953
rect 39284 37901 39286 37953
rect 39230 37899 39286 37901
rect 39773 37276 39829 37332
rect 39992 37507 40048 37563
rect 40251 36999 40307 37055
rect 40431 36999 40487 37055
rect 39773 36722 39829 36778
rect 39992 36491 40048 36547
rect 39050 36153 39106 36155
rect 39050 36101 39052 36153
rect 39052 36101 39104 36153
rect 39104 36101 39106 36153
rect 39050 36099 39106 36101
rect 39230 36153 39286 36155
rect 39230 36101 39232 36153
rect 39232 36101 39284 36153
rect 39284 36101 39286 36153
rect 39230 36099 39286 36101
rect 41881 64898 42041 64954
rect 36958 35825 37014 35881
rect 37169 35825 37225 35881
rect 37381 35825 37437 35881
rect 37592 35825 37648 35881
rect 27478 34968 27534 35024
rect 27690 34968 27746 35024
rect 27478 34750 27534 34806
rect 27690 34750 27729 34806
rect 27729 34750 27746 34806
rect 27478 34532 27534 34588
rect 27690 34532 27746 34588
rect 43788 63999 43844 64055
rect 43999 63999 44055 64055
rect 44211 63999 44267 64055
rect 44422 63999 44478 64055
rect 43788 62199 43844 62255
rect 43999 62199 44055 62255
rect 44211 62199 44267 62255
rect 44422 62199 44478 62255
rect 43788 60399 43844 60455
rect 43999 60399 44055 60455
rect 44211 60399 44267 60455
rect 44422 60399 44478 60455
rect 43788 58599 43844 58655
rect 43999 58599 44055 58655
rect 44211 58599 44267 58655
rect 44422 58599 44478 58655
rect 43788 56799 43844 56855
rect 43999 56799 44055 56855
rect 44211 56799 44267 56855
rect 44422 56799 44478 56855
rect 43788 54999 43844 55055
rect 43999 54999 44055 55055
rect 44211 54999 44267 55055
rect 44422 54999 44478 55055
rect 43788 53199 43844 53255
rect 43999 53199 44055 53255
rect 44211 53199 44267 53255
rect 44422 53199 44478 53255
rect 43788 51399 43844 51455
rect 43999 51399 44055 51455
rect 44211 51399 44267 51455
rect 44422 51399 44478 51455
rect 43788 49599 43844 49655
rect 43999 49599 44055 49655
rect 44211 49599 44267 49655
rect 44422 49599 44478 49655
rect 43788 47799 43844 47855
rect 43999 47799 44055 47855
rect 44211 47799 44267 47855
rect 44422 47799 44478 47855
rect 43788 45999 43844 46055
rect 43999 45999 44055 46055
rect 44211 45999 44267 46055
rect 44422 45999 44478 46055
rect 43788 44199 43844 44255
rect 43999 44199 44055 44255
rect 44211 44199 44267 44255
rect 44422 44199 44478 44255
rect 43788 42399 43844 42455
rect 43999 42399 44055 42455
rect 44211 42399 44267 42455
rect 44422 42399 44478 42455
rect 43788 40599 43844 40655
rect 43999 40599 44055 40655
rect 44211 40599 44267 40655
rect 44422 40599 44478 40655
rect 43788 38799 43844 38855
rect 43999 38799 44055 38855
rect 44211 38799 44267 38855
rect 44422 38799 44478 38855
rect 43788 36999 43844 37055
rect 43999 36999 44055 37055
rect 44211 36999 44267 37055
rect 44422 36999 44478 37055
rect 44832 64953 44888 64955
rect 44832 64901 44834 64953
rect 44834 64901 44886 64953
rect 44886 64901 44888 64953
rect 44832 64899 44888 64901
rect 45043 64953 45099 64955
rect 45043 64901 45045 64953
rect 45045 64901 45097 64953
rect 45097 64901 45099 64953
rect 45043 64899 45099 64901
rect 45254 64953 45310 64955
rect 45254 64901 45256 64953
rect 45256 64901 45308 64953
rect 45308 64901 45310 64953
rect 45254 64899 45310 64901
rect 44832 63153 44888 63155
rect 44832 63101 44834 63153
rect 44834 63101 44886 63153
rect 44886 63101 44888 63153
rect 44832 63099 44888 63101
rect 45043 63153 45099 63155
rect 45043 63101 45045 63153
rect 45045 63101 45097 63153
rect 45097 63101 45099 63153
rect 45043 63099 45099 63101
rect 45254 63153 45310 63155
rect 45254 63101 45256 63153
rect 45256 63101 45308 63153
rect 45308 63101 45310 63153
rect 45254 63099 45310 63101
rect 44832 61353 44888 61355
rect 44832 61301 44834 61353
rect 44834 61301 44886 61353
rect 44886 61301 44888 61353
rect 44832 61299 44888 61301
rect 45043 61353 45099 61355
rect 45043 61301 45045 61353
rect 45045 61301 45097 61353
rect 45097 61301 45099 61353
rect 45043 61299 45099 61301
rect 45254 61353 45310 61355
rect 45254 61301 45256 61353
rect 45256 61301 45308 61353
rect 45308 61301 45310 61353
rect 45254 61299 45310 61301
rect 44832 59553 44888 59555
rect 44832 59501 44834 59553
rect 44834 59501 44886 59553
rect 44886 59501 44888 59553
rect 44832 59499 44888 59501
rect 45043 59553 45099 59555
rect 45043 59501 45045 59553
rect 45045 59501 45097 59553
rect 45097 59501 45099 59553
rect 45043 59499 45099 59501
rect 45254 59553 45310 59555
rect 45254 59501 45256 59553
rect 45256 59501 45308 59553
rect 45308 59501 45310 59553
rect 45254 59499 45310 59501
rect 44832 57753 44888 57755
rect 44832 57701 44834 57753
rect 44834 57701 44886 57753
rect 44886 57701 44888 57753
rect 44832 57699 44888 57701
rect 45043 57753 45099 57755
rect 45043 57701 45045 57753
rect 45045 57701 45097 57753
rect 45097 57701 45099 57753
rect 45043 57699 45099 57701
rect 45254 57753 45310 57755
rect 45254 57701 45256 57753
rect 45256 57701 45308 57753
rect 45308 57701 45310 57753
rect 45254 57699 45310 57701
rect 44832 55953 44888 55955
rect 44832 55901 44834 55953
rect 44834 55901 44886 55953
rect 44886 55901 44888 55953
rect 44832 55899 44888 55901
rect 45043 55953 45099 55955
rect 45043 55901 45045 55953
rect 45045 55901 45097 55953
rect 45097 55901 45099 55953
rect 45043 55899 45099 55901
rect 45254 55953 45310 55955
rect 45254 55901 45256 55953
rect 45256 55901 45308 55953
rect 45308 55901 45310 55953
rect 45254 55899 45310 55901
rect 44832 54153 44888 54155
rect 44832 54101 44834 54153
rect 44834 54101 44886 54153
rect 44886 54101 44888 54153
rect 44832 54099 44888 54101
rect 45043 54153 45099 54155
rect 45043 54101 45045 54153
rect 45045 54101 45097 54153
rect 45097 54101 45099 54153
rect 45043 54099 45099 54101
rect 45254 54153 45310 54155
rect 45254 54101 45256 54153
rect 45256 54101 45308 54153
rect 45308 54101 45310 54153
rect 45254 54099 45310 54101
rect 44832 52353 44888 52355
rect 44832 52301 44834 52353
rect 44834 52301 44886 52353
rect 44886 52301 44888 52353
rect 44832 52299 44888 52301
rect 45043 52353 45099 52355
rect 45043 52301 45045 52353
rect 45045 52301 45097 52353
rect 45097 52301 45099 52353
rect 45043 52299 45099 52301
rect 45254 52353 45310 52355
rect 45254 52301 45256 52353
rect 45256 52301 45308 52353
rect 45308 52301 45310 52353
rect 45254 52299 45310 52301
rect 44832 50553 44888 50555
rect 44832 50501 44834 50553
rect 44834 50501 44886 50553
rect 44886 50501 44888 50553
rect 44832 50499 44888 50501
rect 45043 50553 45099 50555
rect 45043 50501 45045 50553
rect 45045 50501 45097 50553
rect 45097 50501 45099 50553
rect 45043 50499 45099 50501
rect 45254 50553 45310 50555
rect 45254 50501 45256 50553
rect 45256 50501 45308 50553
rect 45308 50501 45310 50553
rect 45254 50499 45310 50501
rect 44832 48753 44888 48755
rect 44832 48701 44834 48753
rect 44834 48701 44886 48753
rect 44886 48701 44888 48753
rect 44832 48699 44888 48701
rect 45043 48753 45099 48755
rect 45043 48701 45045 48753
rect 45045 48701 45097 48753
rect 45097 48701 45099 48753
rect 45043 48699 45099 48701
rect 45254 48753 45310 48755
rect 45254 48701 45256 48753
rect 45256 48701 45308 48753
rect 45308 48701 45310 48753
rect 45254 48699 45310 48701
rect 44832 46953 44888 46955
rect 44832 46901 44834 46953
rect 44834 46901 44886 46953
rect 44886 46901 44888 46953
rect 44832 46899 44888 46901
rect 45043 46953 45099 46955
rect 45043 46901 45045 46953
rect 45045 46901 45097 46953
rect 45097 46901 45099 46953
rect 45043 46899 45099 46901
rect 45254 46953 45310 46955
rect 45254 46901 45256 46953
rect 45256 46901 45308 46953
rect 45308 46901 45310 46953
rect 45254 46899 45310 46901
rect 44832 45153 44888 45155
rect 44832 45101 44834 45153
rect 44834 45101 44886 45153
rect 44886 45101 44888 45153
rect 44832 45099 44888 45101
rect 45043 45153 45099 45155
rect 45043 45101 45045 45153
rect 45045 45101 45097 45153
rect 45097 45101 45099 45153
rect 45043 45099 45099 45101
rect 45254 45153 45310 45155
rect 45254 45101 45256 45153
rect 45256 45101 45308 45153
rect 45308 45101 45310 45153
rect 45254 45099 45310 45101
rect 44832 43353 44888 43355
rect 44832 43301 44834 43353
rect 44834 43301 44886 43353
rect 44886 43301 44888 43353
rect 44832 43299 44888 43301
rect 45043 43353 45099 43355
rect 45043 43301 45045 43353
rect 45045 43301 45097 43353
rect 45097 43301 45099 43353
rect 45043 43299 45099 43301
rect 45254 43353 45310 43355
rect 45254 43301 45256 43353
rect 45256 43301 45308 43353
rect 45308 43301 45310 43353
rect 45254 43299 45310 43301
rect 44832 41553 44888 41555
rect 44832 41501 44834 41553
rect 44834 41501 44886 41553
rect 44886 41501 44888 41553
rect 44832 41499 44888 41501
rect 45043 41553 45099 41555
rect 45043 41501 45045 41553
rect 45045 41501 45097 41553
rect 45097 41501 45099 41553
rect 45043 41499 45099 41501
rect 45254 41553 45310 41555
rect 45254 41501 45256 41553
rect 45256 41501 45308 41553
rect 45308 41501 45310 41553
rect 45254 41499 45310 41501
rect 44832 39753 44888 39755
rect 44832 39701 44834 39753
rect 44834 39701 44886 39753
rect 44886 39701 44888 39753
rect 44832 39699 44888 39701
rect 45043 39753 45099 39755
rect 45043 39701 45045 39753
rect 45045 39701 45097 39753
rect 45097 39701 45099 39753
rect 45043 39699 45099 39701
rect 45254 39753 45310 39755
rect 45254 39701 45256 39753
rect 45256 39701 45308 39753
rect 45308 39701 45310 39753
rect 45254 39699 45310 39701
rect 44832 37953 44888 37955
rect 44832 37901 44834 37953
rect 44834 37901 44886 37953
rect 44886 37901 44888 37953
rect 44832 37899 44888 37901
rect 45043 37953 45099 37955
rect 45043 37901 45045 37953
rect 45045 37901 45097 37953
rect 45097 37901 45099 37953
rect 45043 37899 45099 37901
rect 45254 37953 45310 37955
rect 45254 37901 45256 37953
rect 45256 37901 45308 37953
rect 45308 37901 45310 37953
rect 45254 37899 45310 37901
rect 44832 36153 44888 36155
rect 44832 36101 44834 36153
rect 44834 36101 44886 36153
rect 44886 36101 44888 36153
rect 44832 36099 44888 36101
rect 45043 36153 45099 36155
rect 45043 36101 45045 36153
rect 45045 36101 45097 36153
rect 45097 36101 45099 36153
rect 45043 36099 45099 36101
rect 45254 36153 45310 36155
rect 45254 36101 45256 36153
rect 45256 36101 45308 36153
rect 45308 36101 45310 36153
rect 45254 36099 45310 36101
rect 50135 65853 50191 65855
rect 50135 65801 50137 65853
rect 50137 65801 50189 65853
rect 50189 65801 50191 65853
rect 50135 65799 50191 65801
rect 50346 65853 50402 65855
rect 50346 65801 50348 65853
rect 50348 65801 50400 65853
rect 50400 65801 50402 65853
rect 50346 65799 50402 65801
rect 50557 65853 50613 65855
rect 50557 65801 50559 65853
rect 50559 65801 50611 65853
rect 50611 65801 50613 65853
rect 50557 65799 50613 65801
rect 50768 65853 50824 65855
rect 50768 65801 50770 65853
rect 50770 65801 50822 65853
rect 50822 65801 50824 65853
rect 50768 65799 50824 65801
rect 48836 64953 48892 64955
rect 48836 64901 48838 64953
rect 48838 64901 48890 64953
rect 48890 64901 48892 64953
rect 48836 64899 48892 64901
rect 49046 64953 49102 64955
rect 49046 64901 49048 64953
rect 49048 64901 49100 64953
rect 49100 64901 49102 64953
rect 49046 64899 49102 64901
rect 49257 64953 49313 64955
rect 49257 64901 49259 64953
rect 49259 64901 49311 64953
rect 49311 64901 49313 64953
rect 49257 64899 49313 64901
rect 49469 64953 49525 64955
rect 49469 64901 49471 64953
rect 49471 64901 49523 64953
rect 49523 64901 49525 64953
rect 49469 64899 49525 64901
rect 49680 64953 49736 64955
rect 49680 64901 49682 64953
rect 49682 64901 49734 64953
rect 49734 64901 49736 64953
rect 49680 64899 49736 64901
rect 49890 64953 49946 64955
rect 49890 64901 49892 64953
rect 49892 64901 49944 64953
rect 49944 64901 49946 64953
rect 49890 64899 49946 64901
rect 51079 65370 51135 65372
rect 51079 65318 51081 65370
rect 51081 65318 51133 65370
rect 51133 65318 51135 65370
rect 51079 65316 51135 65318
rect 51290 65370 51346 65372
rect 51290 65318 51292 65370
rect 51292 65318 51344 65370
rect 51344 65318 51346 65370
rect 51290 65316 51346 65318
rect 51501 65370 51557 65372
rect 51501 65318 51503 65370
rect 51503 65318 51555 65370
rect 51555 65318 51557 65370
rect 51501 65316 51557 65318
rect 51712 65370 51768 65372
rect 51712 65318 51714 65370
rect 51714 65318 51766 65370
rect 51766 65318 51768 65370
rect 51712 65316 51768 65318
rect 51923 65370 51979 65372
rect 51923 65318 51925 65370
rect 51925 65318 51977 65370
rect 51977 65318 51979 65370
rect 51923 65316 51979 65318
rect 48594 64547 48650 64549
rect 48594 64495 48596 64547
rect 48596 64495 48648 64547
rect 48648 64495 48650 64547
rect 48594 64493 48650 64495
rect 48594 64329 48650 64331
rect 48594 64277 48596 64329
rect 48596 64277 48648 64329
rect 48648 64277 48650 64329
rect 48594 64275 48650 64277
rect 48594 63777 48650 63779
rect 48594 63725 48596 63777
rect 48596 63725 48648 63777
rect 48648 63725 48650 63777
rect 48594 63723 48650 63725
rect 48594 63559 48650 63561
rect 48594 63507 48596 63559
rect 48596 63507 48648 63559
rect 48648 63507 48650 63559
rect 48594 63505 48650 63507
rect 48836 63153 48892 63155
rect 48836 63101 48838 63153
rect 48838 63101 48890 63153
rect 48890 63101 48892 63153
rect 48836 63099 48892 63101
rect 49046 63153 49102 63155
rect 49046 63101 49048 63153
rect 49048 63101 49100 63153
rect 49100 63101 49102 63153
rect 49046 63099 49102 63101
rect 49257 63153 49313 63155
rect 49257 63101 49259 63153
rect 49259 63101 49311 63153
rect 49311 63101 49313 63153
rect 49257 63099 49313 63101
rect 49469 63153 49525 63155
rect 49469 63101 49471 63153
rect 49471 63101 49523 63153
rect 49523 63101 49525 63153
rect 49469 63099 49525 63101
rect 49680 63153 49736 63155
rect 49680 63101 49682 63153
rect 49682 63101 49734 63153
rect 49734 63101 49736 63153
rect 49680 63099 49736 63101
rect 49890 63153 49946 63155
rect 49890 63101 49892 63153
rect 49892 63101 49944 63153
rect 49944 63101 49946 63153
rect 49890 63099 49946 63101
rect 48594 62747 48650 62749
rect 48594 62695 48596 62747
rect 48596 62695 48648 62747
rect 48648 62695 48650 62747
rect 48594 62693 48650 62695
rect 48594 62529 48650 62531
rect 48594 62477 48596 62529
rect 48596 62477 48648 62529
rect 48648 62477 48650 62529
rect 48594 62475 48650 62477
rect 48594 61977 48650 61979
rect 48594 61925 48596 61977
rect 48596 61925 48648 61977
rect 48648 61925 48650 61977
rect 48594 61923 48650 61925
rect 48594 61759 48650 61761
rect 48594 61707 48596 61759
rect 48596 61707 48648 61759
rect 48648 61707 48650 61759
rect 48594 61705 48650 61707
rect 48836 61353 48892 61355
rect 48836 61301 48838 61353
rect 48838 61301 48890 61353
rect 48890 61301 48892 61353
rect 48836 61299 48892 61301
rect 49046 61353 49102 61355
rect 49046 61301 49048 61353
rect 49048 61301 49100 61353
rect 49100 61301 49102 61353
rect 49046 61299 49102 61301
rect 49257 61353 49313 61355
rect 49257 61301 49259 61353
rect 49259 61301 49311 61353
rect 49311 61301 49313 61353
rect 49257 61299 49313 61301
rect 49469 61353 49525 61355
rect 49469 61301 49471 61353
rect 49471 61301 49523 61353
rect 49523 61301 49525 61353
rect 49469 61299 49525 61301
rect 49680 61353 49736 61355
rect 49680 61301 49682 61353
rect 49682 61301 49734 61353
rect 49734 61301 49736 61353
rect 49680 61299 49736 61301
rect 49890 61353 49946 61355
rect 49890 61301 49892 61353
rect 49892 61301 49944 61353
rect 49944 61301 49946 61353
rect 49890 61299 49946 61301
rect 48594 60947 48650 60949
rect 48594 60895 48596 60947
rect 48596 60895 48648 60947
rect 48648 60895 48650 60947
rect 48594 60893 48650 60895
rect 48594 60729 48650 60731
rect 48594 60677 48596 60729
rect 48596 60677 48648 60729
rect 48648 60677 48650 60729
rect 48594 60675 48650 60677
rect 48594 60177 48650 60179
rect 48594 60125 48596 60177
rect 48596 60125 48648 60177
rect 48648 60125 48650 60177
rect 48594 60123 48650 60125
rect 48594 59959 48650 59961
rect 48594 59907 48596 59959
rect 48596 59907 48648 59959
rect 48648 59907 48650 59959
rect 48594 59905 48650 59907
rect 48836 59553 48892 59555
rect 48836 59501 48838 59553
rect 48838 59501 48890 59553
rect 48890 59501 48892 59553
rect 48836 59499 48892 59501
rect 49046 59553 49102 59555
rect 49046 59501 49048 59553
rect 49048 59501 49100 59553
rect 49100 59501 49102 59553
rect 49046 59499 49102 59501
rect 49257 59553 49313 59555
rect 49257 59501 49259 59553
rect 49259 59501 49311 59553
rect 49311 59501 49313 59553
rect 49257 59499 49313 59501
rect 49469 59553 49525 59555
rect 49469 59501 49471 59553
rect 49471 59501 49523 59553
rect 49523 59501 49525 59553
rect 49469 59499 49525 59501
rect 49680 59553 49736 59555
rect 49680 59501 49682 59553
rect 49682 59501 49734 59553
rect 49734 59501 49736 59553
rect 49680 59499 49736 59501
rect 49890 59553 49946 59555
rect 49890 59501 49892 59553
rect 49892 59501 49944 59553
rect 49944 59501 49946 59553
rect 49890 59499 49946 59501
rect 48594 59147 48650 59149
rect 48594 59095 48596 59147
rect 48596 59095 48648 59147
rect 48648 59095 48650 59147
rect 48594 59093 48650 59095
rect 48594 58929 48650 58931
rect 48594 58877 48596 58929
rect 48596 58877 48648 58929
rect 48648 58877 48650 58929
rect 48594 58875 48650 58877
rect 48594 58377 48650 58379
rect 48594 58325 48596 58377
rect 48596 58325 48648 58377
rect 48648 58325 48650 58377
rect 48594 58323 48650 58325
rect 48594 58159 48650 58161
rect 48594 58107 48596 58159
rect 48596 58107 48648 58159
rect 48648 58107 48650 58159
rect 48594 58105 48650 58107
rect 48836 57753 48892 57755
rect 48836 57701 48838 57753
rect 48838 57701 48890 57753
rect 48890 57701 48892 57753
rect 48836 57699 48892 57701
rect 49046 57753 49102 57755
rect 49046 57701 49048 57753
rect 49048 57701 49100 57753
rect 49100 57701 49102 57753
rect 49046 57699 49102 57701
rect 49257 57753 49313 57755
rect 49257 57701 49259 57753
rect 49259 57701 49311 57753
rect 49311 57701 49313 57753
rect 49257 57699 49313 57701
rect 49469 57753 49525 57755
rect 49469 57701 49471 57753
rect 49471 57701 49523 57753
rect 49523 57701 49525 57753
rect 49469 57699 49525 57701
rect 49680 57753 49736 57755
rect 49680 57701 49682 57753
rect 49682 57701 49734 57753
rect 49734 57701 49736 57753
rect 49680 57699 49736 57701
rect 49890 57753 49946 57755
rect 49890 57701 49892 57753
rect 49892 57701 49944 57753
rect 49944 57701 49946 57753
rect 49890 57699 49946 57701
rect 48594 57347 48650 57349
rect 48594 57295 48596 57347
rect 48596 57295 48648 57347
rect 48648 57295 48650 57347
rect 48594 57293 48650 57295
rect 48594 57129 48650 57131
rect 48594 57077 48596 57129
rect 48596 57077 48648 57129
rect 48648 57077 48650 57129
rect 48594 57075 48650 57077
rect 48594 56577 48650 56579
rect 48594 56525 48596 56577
rect 48596 56525 48648 56577
rect 48648 56525 48650 56577
rect 48594 56523 48650 56525
rect 48594 56359 48650 56361
rect 48594 56307 48596 56359
rect 48596 56307 48648 56359
rect 48648 56307 48650 56359
rect 48594 56305 48650 56307
rect 48836 55953 48892 55955
rect 48836 55901 48838 55953
rect 48838 55901 48890 55953
rect 48890 55901 48892 55953
rect 48836 55899 48892 55901
rect 49046 55953 49102 55955
rect 49046 55901 49048 55953
rect 49048 55901 49100 55953
rect 49100 55901 49102 55953
rect 49046 55899 49102 55901
rect 49257 55953 49313 55955
rect 49257 55901 49259 55953
rect 49259 55901 49311 55953
rect 49311 55901 49313 55953
rect 49257 55899 49313 55901
rect 49469 55953 49525 55955
rect 49469 55901 49471 55953
rect 49471 55901 49523 55953
rect 49523 55901 49525 55953
rect 49469 55899 49525 55901
rect 49680 55953 49736 55955
rect 49680 55901 49682 55953
rect 49682 55901 49734 55953
rect 49734 55901 49736 55953
rect 49680 55899 49736 55901
rect 49890 55953 49946 55955
rect 49890 55901 49892 55953
rect 49892 55901 49944 55953
rect 49944 55901 49946 55953
rect 49890 55899 49946 55901
rect 48594 55547 48650 55549
rect 48594 55495 48596 55547
rect 48596 55495 48648 55547
rect 48648 55495 48650 55547
rect 48594 55493 48650 55495
rect 48594 55329 48650 55331
rect 48594 55277 48596 55329
rect 48596 55277 48648 55329
rect 48648 55277 48650 55329
rect 48594 55275 48650 55277
rect 48594 54777 48650 54779
rect 48594 54725 48596 54777
rect 48596 54725 48648 54777
rect 48648 54725 48650 54777
rect 48594 54723 48650 54725
rect 48594 54559 48650 54561
rect 48594 54507 48596 54559
rect 48596 54507 48648 54559
rect 48648 54507 48650 54559
rect 48594 54505 48650 54507
rect 48836 54153 48892 54155
rect 48836 54101 48838 54153
rect 48838 54101 48890 54153
rect 48890 54101 48892 54153
rect 48836 54099 48892 54101
rect 49046 54153 49102 54155
rect 49046 54101 49048 54153
rect 49048 54101 49100 54153
rect 49100 54101 49102 54153
rect 49046 54099 49102 54101
rect 49257 54153 49313 54155
rect 49257 54101 49259 54153
rect 49259 54101 49311 54153
rect 49311 54101 49313 54153
rect 49257 54099 49313 54101
rect 49469 54153 49525 54155
rect 49469 54101 49471 54153
rect 49471 54101 49523 54153
rect 49523 54101 49525 54153
rect 49469 54099 49525 54101
rect 49680 54153 49736 54155
rect 49680 54101 49682 54153
rect 49682 54101 49734 54153
rect 49734 54101 49736 54153
rect 49680 54099 49736 54101
rect 49890 54153 49946 54155
rect 49890 54101 49892 54153
rect 49892 54101 49944 54153
rect 49944 54101 49946 54153
rect 49890 54099 49946 54101
rect 48594 53747 48650 53749
rect 48594 53695 48596 53747
rect 48596 53695 48648 53747
rect 48648 53695 48650 53747
rect 48594 53693 48650 53695
rect 48594 53529 48650 53531
rect 48594 53477 48596 53529
rect 48596 53477 48648 53529
rect 48648 53477 48650 53529
rect 48594 53475 48650 53477
rect 48594 52977 48650 52979
rect 48594 52925 48596 52977
rect 48596 52925 48648 52977
rect 48648 52925 48650 52977
rect 48594 52923 48650 52925
rect 48594 52759 48650 52761
rect 48594 52707 48596 52759
rect 48596 52707 48648 52759
rect 48648 52707 48650 52759
rect 48594 52705 48650 52707
rect 48836 52353 48892 52355
rect 48836 52301 48838 52353
rect 48838 52301 48890 52353
rect 48890 52301 48892 52353
rect 48836 52299 48892 52301
rect 49046 52353 49102 52355
rect 49046 52301 49048 52353
rect 49048 52301 49100 52353
rect 49100 52301 49102 52353
rect 49046 52299 49102 52301
rect 49257 52353 49313 52355
rect 49257 52301 49259 52353
rect 49259 52301 49311 52353
rect 49311 52301 49313 52353
rect 49257 52299 49313 52301
rect 49469 52353 49525 52355
rect 49469 52301 49471 52353
rect 49471 52301 49523 52353
rect 49523 52301 49525 52353
rect 49469 52299 49525 52301
rect 49680 52353 49736 52355
rect 49680 52301 49682 52353
rect 49682 52301 49734 52353
rect 49734 52301 49736 52353
rect 49680 52299 49736 52301
rect 49890 52353 49946 52355
rect 49890 52301 49892 52353
rect 49892 52301 49944 52353
rect 49944 52301 49946 52353
rect 49890 52299 49946 52301
rect 48594 51947 48650 51949
rect 48594 51895 48596 51947
rect 48596 51895 48648 51947
rect 48648 51895 48650 51947
rect 48594 51893 48650 51895
rect 48594 51729 48650 51731
rect 48594 51677 48596 51729
rect 48596 51677 48648 51729
rect 48648 51677 48650 51729
rect 48594 51675 48650 51677
rect 48594 51177 48650 51179
rect 48594 51125 48596 51177
rect 48596 51125 48648 51177
rect 48648 51125 48650 51177
rect 48594 51123 48650 51125
rect 48594 50959 48650 50961
rect 48594 50907 48596 50959
rect 48596 50907 48648 50959
rect 48648 50907 48650 50959
rect 48594 50905 48650 50907
rect 48836 50553 48892 50555
rect 48836 50501 48838 50553
rect 48838 50501 48890 50553
rect 48890 50501 48892 50553
rect 48836 50499 48892 50501
rect 49046 50553 49102 50555
rect 49046 50501 49048 50553
rect 49048 50501 49100 50553
rect 49100 50501 49102 50553
rect 49046 50499 49102 50501
rect 49257 50553 49313 50555
rect 49257 50501 49259 50553
rect 49259 50501 49311 50553
rect 49311 50501 49313 50553
rect 49257 50499 49313 50501
rect 49469 50553 49525 50555
rect 49469 50501 49471 50553
rect 49471 50501 49523 50553
rect 49523 50501 49525 50553
rect 49469 50499 49525 50501
rect 49680 50553 49736 50555
rect 49680 50501 49682 50553
rect 49682 50501 49734 50553
rect 49734 50501 49736 50553
rect 49680 50499 49736 50501
rect 49890 50553 49946 50555
rect 49890 50501 49892 50553
rect 49892 50501 49944 50553
rect 49944 50501 49946 50553
rect 49890 50499 49946 50501
rect 48594 50147 48650 50149
rect 48594 50095 48596 50147
rect 48596 50095 48648 50147
rect 48648 50095 48650 50147
rect 48594 50093 48650 50095
rect 48594 49929 48650 49931
rect 48594 49877 48596 49929
rect 48596 49877 48648 49929
rect 48648 49877 48650 49929
rect 48594 49875 48650 49877
rect 48594 49377 48650 49379
rect 48594 49325 48596 49377
rect 48596 49325 48648 49377
rect 48648 49325 48650 49377
rect 48594 49323 48650 49325
rect 48594 49159 48650 49161
rect 48594 49107 48596 49159
rect 48596 49107 48648 49159
rect 48648 49107 48650 49159
rect 48594 49105 48650 49107
rect 48836 48753 48892 48755
rect 48836 48701 48838 48753
rect 48838 48701 48890 48753
rect 48890 48701 48892 48753
rect 48836 48699 48892 48701
rect 49046 48753 49102 48755
rect 49046 48701 49048 48753
rect 49048 48701 49100 48753
rect 49100 48701 49102 48753
rect 49046 48699 49102 48701
rect 49257 48753 49313 48755
rect 49257 48701 49259 48753
rect 49259 48701 49311 48753
rect 49311 48701 49313 48753
rect 49257 48699 49313 48701
rect 49469 48753 49525 48755
rect 49469 48701 49471 48753
rect 49471 48701 49523 48753
rect 49523 48701 49525 48753
rect 49469 48699 49525 48701
rect 49680 48753 49736 48755
rect 49680 48701 49682 48753
rect 49682 48701 49734 48753
rect 49734 48701 49736 48753
rect 49680 48699 49736 48701
rect 49890 48753 49946 48755
rect 49890 48701 49892 48753
rect 49892 48701 49944 48753
rect 49944 48701 49946 48753
rect 49890 48699 49946 48701
rect 48594 48347 48650 48349
rect 48594 48295 48596 48347
rect 48596 48295 48648 48347
rect 48648 48295 48650 48347
rect 48594 48293 48650 48295
rect 48594 48129 48650 48131
rect 48594 48077 48596 48129
rect 48596 48077 48648 48129
rect 48648 48077 48650 48129
rect 48594 48075 48650 48077
rect 48594 47577 48650 47579
rect 48594 47525 48596 47577
rect 48596 47525 48648 47577
rect 48648 47525 48650 47577
rect 48594 47523 48650 47525
rect 48594 47359 48650 47361
rect 48594 47307 48596 47359
rect 48596 47307 48648 47359
rect 48648 47307 48650 47359
rect 48594 47305 48650 47307
rect 48836 46953 48892 46955
rect 48836 46901 48838 46953
rect 48838 46901 48890 46953
rect 48890 46901 48892 46953
rect 48836 46899 48892 46901
rect 49046 46953 49102 46955
rect 49046 46901 49048 46953
rect 49048 46901 49100 46953
rect 49100 46901 49102 46953
rect 49046 46899 49102 46901
rect 49257 46953 49313 46955
rect 49257 46901 49259 46953
rect 49259 46901 49311 46953
rect 49311 46901 49313 46953
rect 49257 46899 49313 46901
rect 49469 46953 49525 46955
rect 49469 46901 49471 46953
rect 49471 46901 49523 46953
rect 49523 46901 49525 46953
rect 49469 46899 49525 46901
rect 49680 46953 49736 46955
rect 49680 46901 49682 46953
rect 49682 46901 49734 46953
rect 49734 46901 49736 46953
rect 49680 46899 49736 46901
rect 49890 46953 49946 46955
rect 49890 46901 49892 46953
rect 49892 46901 49944 46953
rect 49944 46901 49946 46953
rect 49890 46899 49946 46901
rect 48594 46547 48650 46549
rect 48594 46495 48596 46547
rect 48596 46495 48648 46547
rect 48648 46495 48650 46547
rect 48594 46493 48650 46495
rect 48594 46329 48650 46331
rect 48594 46277 48596 46329
rect 48596 46277 48648 46329
rect 48648 46277 48650 46329
rect 48594 46275 48650 46277
rect 48594 45777 48650 45779
rect 48594 45725 48596 45777
rect 48596 45725 48648 45777
rect 48648 45725 48650 45777
rect 48594 45723 48650 45725
rect 48594 45559 48650 45561
rect 48594 45507 48596 45559
rect 48596 45507 48648 45559
rect 48648 45507 48650 45559
rect 48594 45505 48650 45507
rect 48836 45153 48892 45155
rect 48836 45101 48838 45153
rect 48838 45101 48890 45153
rect 48890 45101 48892 45153
rect 48836 45099 48892 45101
rect 49046 45153 49102 45155
rect 49046 45101 49048 45153
rect 49048 45101 49100 45153
rect 49100 45101 49102 45153
rect 49046 45099 49102 45101
rect 49257 45153 49313 45155
rect 49257 45101 49259 45153
rect 49259 45101 49311 45153
rect 49311 45101 49313 45153
rect 49257 45099 49313 45101
rect 49469 45153 49525 45155
rect 49469 45101 49471 45153
rect 49471 45101 49523 45153
rect 49523 45101 49525 45153
rect 49469 45099 49525 45101
rect 49680 45153 49736 45155
rect 49680 45101 49682 45153
rect 49682 45101 49734 45153
rect 49734 45101 49736 45153
rect 49680 45099 49736 45101
rect 49890 45153 49946 45155
rect 49890 45101 49892 45153
rect 49892 45101 49944 45153
rect 49944 45101 49946 45153
rect 49890 45099 49946 45101
rect 48594 44747 48650 44749
rect 48594 44695 48596 44747
rect 48596 44695 48648 44747
rect 48648 44695 48650 44747
rect 48594 44693 48650 44695
rect 48594 44529 48650 44531
rect 48594 44477 48596 44529
rect 48596 44477 48648 44529
rect 48648 44477 48650 44529
rect 48594 44475 48650 44477
rect 48594 43977 48650 43979
rect 48594 43925 48596 43977
rect 48596 43925 48648 43977
rect 48648 43925 48650 43977
rect 48594 43923 48650 43925
rect 48594 43759 48650 43761
rect 48594 43707 48596 43759
rect 48596 43707 48648 43759
rect 48648 43707 48650 43759
rect 48594 43705 48650 43707
rect 48836 43353 48892 43355
rect 48836 43301 48838 43353
rect 48838 43301 48890 43353
rect 48890 43301 48892 43353
rect 48836 43299 48892 43301
rect 49046 43353 49102 43355
rect 49046 43301 49048 43353
rect 49048 43301 49100 43353
rect 49100 43301 49102 43353
rect 49046 43299 49102 43301
rect 49257 43353 49313 43355
rect 49257 43301 49259 43353
rect 49259 43301 49311 43353
rect 49311 43301 49313 43353
rect 49257 43299 49313 43301
rect 49469 43353 49525 43355
rect 49469 43301 49471 43353
rect 49471 43301 49523 43353
rect 49523 43301 49525 43353
rect 49469 43299 49525 43301
rect 49680 43353 49736 43355
rect 49680 43301 49682 43353
rect 49682 43301 49734 43353
rect 49734 43301 49736 43353
rect 49680 43299 49736 43301
rect 49890 43353 49946 43355
rect 49890 43301 49892 43353
rect 49892 43301 49944 43353
rect 49944 43301 49946 43353
rect 49890 43299 49946 43301
rect 48594 42947 48650 42949
rect 48594 42895 48596 42947
rect 48596 42895 48648 42947
rect 48648 42895 48650 42947
rect 48594 42893 48650 42895
rect 48594 42729 48650 42731
rect 48594 42677 48596 42729
rect 48596 42677 48648 42729
rect 48648 42677 48650 42729
rect 48594 42675 48650 42677
rect 48594 42177 48650 42179
rect 48594 42125 48596 42177
rect 48596 42125 48648 42177
rect 48648 42125 48650 42177
rect 48594 42123 48650 42125
rect 48594 41959 48650 41961
rect 48594 41907 48596 41959
rect 48596 41907 48648 41959
rect 48648 41907 48650 41959
rect 48594 41905 48650 41907
rect 48836 41553 48892 41555
rect 48836 41501 48838 41553
rect 48838 41501 48890 41553
rect 48890 41501 48892 41553
rect 48836 41499 48892 41501
rect 49046 41553 49102 41555
rect 49046 41501 49048 41553
rect 49048 41501 49100 41553
rect 49100 41501 49102 41553
rect 49046 41499 49102 41501
rect 49257 41553 49313 41555
rect 49257 41501 49259 41553
rect 49259 41501 49311 41553
rect 49311 41501 49313 41553
rect 49257 41499 49313 41501
rect 49469 41553 49525 41555
rect 49469 41501 49471 41553
rect 49471 41501 49523 41553
rect 49523 41501 49525 41553
rect 49469 41499 49525 41501
rect 49680 41553 49736 41555
rect 49680 41501 49682 41553
rect 49682 41501 49734 41553
rect 49734 41501 49736 41553
rect 49680 41499 49736 41501
rect 49890 41553 49946 41555
rect 49890 41501 49892 41553
rect 49892 41501 49944 41553
rect 49944 41501 49946 41553
rect 49890 41499 49946 41501
rect 48594 41147 48650 41149
rect 48594 41095 48596 41147
rect 48596 41095 48648 41147
rect 48648 41095 48650 41147
rect 48594 41093 48650 41095
rect 48594 40929 48650 40931
rect 48594 40877 48596 40929
rect 48596 40877 48648 40929
rect 48648 40877 48650 40929
rect 48594 40875 48650 40877
rect 48594 40377 48650 40379
rect 48594 40325 48596 40377
rect 48596 40325 48648 40377
rect 48648 40325 48650 40377
rect 48594 40323 48650 40325
rect 48594 40159 48650 40161
rect 48594 40107 48596 40159
rect 48596 40107 48648 40159
rect 48648 40107 48650 40159
rect 48594 40105 48650 40107
rect 48836 39753 48892 39755
rect 48836 39701 48838 39753
rect 48838 39701 48890 39753
rect 48890 39701 48892 39753
rect 48836 39699 48892 39701
rect 49046 39753 49102 39755
rect 49046 39701 49048 39753
rect 49048 39701 49100 39753
rect 49100 39701 49102 39753
rect 49046 39699 49102 39701
rect 49257 39753 49313 39755
rect 49257 39701 49259 39753
rect 49259 39701 49311 39753
rect 49311 39701 49313 39753
rect 49257 39699 49313 39701
rect 49469 39753 49525 39755
rect 49469 39701 49471 39753
rect 49471 39701 49523 39753
rect 49523 39701 49525 39753
rect 49469 39699 49525 39701
rect 49680 39753 49736 39755
rect 49680 39701 49682 39753
rect 49682 39701 49734 39753
rect 49734 39701 49736 39753
rect 49680 39699 49736 39701
rect 49890 39753 49946 39755
rect 49890 39701 49892 39753
rect 49892 39701 49944 39753
rect 49944 39701 49946 39753
rect 49890 39699 49946 39701
rect 48594 39347 48650 39349
rect 48594 39295 48596 39347
rect 48596 39295 48648 39347
rect 48648 39295 48650 39347
rect 48594 39293 48650 39295
rect 48594 39129 48650 39131
rect 48594 39077 48596 39129
rect 48596 39077 48648 39129
rect 48648 39077 48650 39129
rect 48594 39075 48650 39077
rect 48594 38577 48650 38579
rect 48594 38525 48596 38577
rect 48596 38525 48648 38577
rect 48648 38525 48650 38577
rect 48594 38523 48650 38525
rect 48594 38359 48650 38361
rect 48594 38307 48596 38359
rect 48596 38307 48648 38359
rect 48648 38307 48650 38359
rect 48594 38305 48650 38307
rect 48836 37953 48892 37955
rect 48836 37901 48838 37953
rect 48838 37901 48890 37953
rect 48890 37901 48892 37953
rect 48836 37899 48892 37901
rect 49046 37953 49102 37955
rect 49046 37901 49048 37953
rect 49048 37901 49100 37953
rect 49100 37901 49102 37953
rect 49046 37899 49102 37901
rect 49257 37953 49313 37955
rect 49257 37901 49259 37953
rect 49259 37901 49311 37953
rect 49311 37901 49313 37953
rect 49257 37899 49313 37901
rect 49469 37953 49525 37955
rect 49469 37901 49471 37953
rect 49471 37901 49523 37953
rect 49523 37901 49525 37953
rect 49469 37899 49525 37901
rect 49680 37953 49736 37955
rect 49680 37901 49682 37953
rect 49682 37901 49734 37953
rect 49734 37901 49736 37953
rect 49680 37899 49736 37901
rect 49890 37953 49946 37955
rect 49890 37901 49892 37953
rect 49892 37901 49944 37953
rect 49944 37901 49946 37953
rect 49890 37899 49946 37901
rect 48594 37547 48650 37549
rect 48594 37495 48596 37547
rect 48596 37495 48648 37547
rect 48648 37495 48650 37547
rect 48594 37493 48650 37495
rect 48594 37329 48650 37331
rect 48594 37277 48596 37329
rect 48596 37277 48648 37329
rect 48648 37277 48650 37329
rect 48594 37275 48650 37277
rect 48594 36777 48650 36779
rect 48594 36725 48596 36777
rect 48596 36725 48648 36777
rect 48648 36725 48650 36777
rect 48594 36723 48650 36725
rect 48594 36559 48650 36561
rect 48594 36507 48596 36559
rect 48596 36507 48648 36559
rect 48648 36507 48650 36559
rect 48594 36505 48650 36507
rect 48836 36153 48892 36155
rect 48836 36101 48838 36153
rect 48838 36101 48890 36153
rect 48890 36101 48892 36153
rect 48836 36099 48892 36101
rect 49046 36153 49102 36155
rect 49046 36101 49048 36153
rect 49048 36101 49100 36153
rect 49100 36101 49102 36153
rect 49046 36099 49102 36101
rect 49257 36153 49313 36155
rect 49257 36101 49259 36153
rect 49259 36101 49311 36153
rect 49311 36101 49313 36153
rect 49257 36099 49313 36101
rect 49469 36153 49525 36155
rect 49469 36101 49471 36153
rect 49471 36101 49523 36153
rect 49523 36101 49525 36153
rect 49469 36099 49525 36101
rect 49680 36153 49736 36155
rect 49680 36101 49682 36153
rect 49682 36101 49734 36153
rect 49734 36101 49736 36153
rect 49680 36099 49736 36101
rect 49890 36153 49946 36155
rect 49890 36101 49892 36153
rect 49892 36101 49944 36153
rect 49944 36101 49946 36153
rect 49890 36099 49946 36101
rect 52314 64953 52370 64955
rect 52314 64901 52316 64953
rect 52316 64901 52368 64953
rect 52368 64901 52370 64953
rect 52314 64899 52370 64901
rect 52525 64953 52581 64955
rect 52525 64901 52527 64953
rect 52527 64901 52579 64953
rect 52579 64901 52581 64953
rect 52525 64899 52581 64901
rect 52736 64953 52792 64955
rect 52736 64901 52738 64953
rect 52738 64901 52790 64953
rect 52790 64901 52792 64953
rect 52736 64899 52792 64901
rect 52946 64953 53002 64955
rect 52946 64901 52948 64953
rect 52948 64901 53000 64953
rect 53000 64901 53002 64953
rect 52946 64899 53002 64901
rect 53157 64953 53213 64955
rect 53157 64901 53159 64953
rect 53159 64901 53211 64953
rect 53211 64901 53213 64953
rect 53157 64899 53213 64901
rect 53369 64953 53425 64955
rect 53369 64901 53371 64953
rect 53371 64901 53423 64953
rect 53423 64901 53425 64953
rect 53369 64899 53425 64901
rect 53580 64953 53636 64955
rect 53580 64901 53582 64953
rect 53582 64901 53634 64953
rect 53634 64901 53636 64953
rect 53580 64899 53636 64901
rect 53790 64953 53846 64955
rect 53790 64901 53792 64953
rect 53792 64901 53844 64953
rect 53844 64901 53846 64953
rect 53790 64899 53846 64901
rect 54001 64953 54057 64955
rect 54001 64901 54003 64953
rect 54003 64901 54055 64953
rect 54055 64901 54057 64953
rect 54001 64899 54057 64901
rect 54212 64953 54268 64955
rect 54212 64901 54214 64953
rect 54214 64901 54266 64953
rect 54266 64901 54268 64953
rect 54212 64899 54268 64901
rect 51071 64459 51127 64515
rect 51251 64459 51307 64515
rect 51833 64459 51889 64515
rect 52013 64459 52069 64515
rect 50161 64053 50217 64055
rect 50161 64001 50190 64053
rect 50190 64001 50217 64053
rect 50161 63999 50217 64001
rect 50372 63999 50428 64055
rect 50584 63999 50640 64055
rect 50795 63999 50851 64055
rect 51071 63539 51127 63595
rect 51251 63539 51307 63595
rect 51833 63539 51889 63595
rect 52013 63539 52069 63595
rect 52314 63153 52370 63155
rect 52314 63101 52316 63153
rect 52316 63101 52368 63153
rect 52368 63101 52370 63153
rect 52314 63099 52370 63101
rect 52525 63153 52581 63155
rect 52525 63101 52527 63153
rect 52527 63101 52579 63153
rect 52579 63101 52581 63153
rect 52525 63099 52581 63101
rect 52736 63153 52792 63155
rect 52736 63101 52738 63153
rect 52738 63101 52790 63153
rect 52790 63101 52792 63153
rect 52736 63099 52792 63101
rect 52946 63153 53002 63155
rect 52946 63101 52948 63153
rect 52948 63101 53000 63153
rect 53000 63101 53002 63153
rect 52946 63099 53002 63101
rect 53157 63153 53213 63155
rect 53157 63101 53159 63153
rect 53159 63101 53211 63153
rect 53211 63101 53213 63153
rect 53157 63099 53213 63101
rect 53369 63153 53425 63155
rect 53369 63101 53371 63153
rect 53371 63101 53423 63153
rect 53423 63101 53425 63153
rect 53369 63099 53425 63101
rect 53580 63153 53636 63155
rect 53580 63101 53582 63153
rect 53582 63101 53634 63153
rect 53634 63101 53636 63153
rect 53580 63099 53636 63101
rect 53790 63153 53846 63155
rect 53790 63101 53792 63153
rect 53792 63101 53844 63153
rect 53844 63101 53846 63153
rect 53790 63099 53846 63101
rect 54001 63153 54057 63155
rect 54001 63101 54003 63153
rect 54003 63101 54055 63153
rect 54055 63101 54057 63153
rect 54001 63099 54057 63101
rect 54212 63153 54268 63155
rect 54212 63101 54214 63153
rect 54214 63101 54266 63153
rect 54266 63101 54268 63153
rect 54212 63099 54268 63101
rect 51071 62659 51127 62715
rect 51251 62659 51307 62715
rect 51833 62659 51889 62715
rect 52013 62659 52069 62715
rect 50161 62253 50217 62255
rect 50161 62201 50190 62253
rect 50190 62201 50217 62253
rect 50161 62199 50217 62201
rect 50372 62199 50428 62255
rect 50584 62199 50640 62255
rect 50795 62199 50851 62255
rect 51071 61739 51127 61795
rect 51251 61739 51307 61795
rect 51833 61739 51889 61795
rect 52013 61739 52069 61795
rect 52314 61353 52370 61355
rect 52314 61301 52316 61353
rect 52316 61301 52368 61353
rect 52368 61301 52370 61353
rect 52314 61299 52370 61301
rect 52525 61353 52581 61355
rect 52525 61301 52527 61353
rect 52527 61301 52579 61353
rect 52579 61301 52581 61353
rect 52525 61299 52581 61301
rect 52736 61353 52792 61355
rect 52736 61301 52738 61353
rect 52738 61301 52790 61353
rect 52790 61301 52792 61353
rect 52736 61299 52792 61301
rect 52946 61353 53002 61355
rect 52946 61301 52948 61353
rect 52948 61301 53000 61353
rect 53000 61301 53002 61353
rect 52946 61299 53002 61301
rect 53157 61353 53213 61355
rect 53157 61301 53159 61353
rect 53159 61301 53211 61353
rect 53211 61301 53213 61353
rect 53157 61299 53213 61301
rect 53369 61353 53425 61355
rect 53369 61301 53371 61353
rect 53371 61301 53423 61353
rect 53423 61301 53425 61353
rect 53369 61299 53425 61301
rect 53580 61353 53636 61355
rect 53580 61301 53582 61353
rect 53582 61301 53634 61353
rect 53634 61301 53636 61353
rect 53580 61299 53636 61301
rect 53790 61353 53846 61355
rect 53790 61301 53792 61353
rect 53792 61301 53844 61353
rect 53844 61301 53846 61353
rect 53790 61299 53846 61301
rect 54001 61353 54057 61355
rect 54001 61301 54003 61353
rect 54003 61301 54055 61353
rect 54055 61301 54057 61353
rect 54001 61299 54057 61301
rect 54212 61353 54268 61355
rect 54212 61301 54214 61353
rect 54214 61301 54266 61353
rect 54266 61301 54268 61353
rect 54212 61299 54268 61301
rect 51071 60859 51127 60915
rect 51251 60859 51307 60915
rect 51833 60859 51889 60915
rect 52013 60859 52069 60915
rect 50161 60453 50217 60455
rect 50161 60401 50190 60453
rect 50190 60401 50217 60453
rect 50161 60399 50217 60401
rect 50372 60399 50428 60455
rect 50584 60399 50640 60455
rect 50795 60399 50851 60455
rect 51071 59939 51127 59995
rect 51251 59939 51307 59995
rect 51833 59939 51889 59995
rect 52013 59939 52069 59995
rect 52314 59553 52370 59555
rect 52314 59501 52316 59553
rect 52316 59501 52368 59553
rect 52368 59501 52370 59553
rect 52314 59499 52370 59501
rect 52525 59553 52581 59555
rect 52525 59501 52527 59553
rect 52527 59501 52579 59553
rect 52579 59501 52581 59553
rect 52525 59499 52581 59501
rect 52736 59553 52792 59555
rect 52736 59501 52738 59553
rect 52738 59501 52790 59553
rect 52790 59501 52792 59553
rect 52736 59499 52792 59501
rect 52946 59553 53002 59555
rect 52946 59501 52948 59553
rect 52948 59501 53000 59553
rect 53000 59501 53002 59553
rect 52946 59499 53002 59501
rect 53157 59553 53213 59555
rect 53157 59501 53159 59553
rect 53159 59501 53211 59553
rect 53211 59501 53213 59553
rect 53157 59499 53213 59501
rect 53369 59553 53425 59555
rect 53369 59501 53371 59553
rect 53371 59501 53423 59553
rect 53423 59501 53425 59553
rect 53369 59499 53425 59501
rect 53580 59553 53636 59555
rect 53580 59501 53582 59553
rect 53582 59501 53634 59553
rect 53634 59501 53636 59553
rect 53580 59499 53636 59501
rect 53790 59553 53846 59555
rect 53790 59501 53792 59553
rect 53792 59501 53844 59553
rect 53844 59501 53846 59553
rect 53790 59499 53846 59501
rect 54001 59553 54057 59555
rect 54001 59501 54003 59553
rect 54003 59501 54055 59553
rect 54055 59501 54057 59553
rect 54001 59499 54057 59501
rect 54212 59553 54268 59555
rect 54212 59501 54214 59553
rect 54214 59501 54266 59553
rect 54266 59501 54268 59553
rect 54212 59499 54268 59501
rect 51071 59059 51127 59115
rect 51251 59059 51307 59115
rect 51833 59059 51889 59115
rect 52013 59059 52069 59115
rect 50161 58653 50217 58655
rect 50161 58601 50190 58653
rect 50190 58601 50217 58653
rect 50161 58599 50217 58601
rect 50372 58599 50428 58655
rect 50584 58599 50640 58655
rect 50795 58599 50851 58655
rect 51071 58139 51127 58195
rect 51251 58139 51307 58195
rect 51833 58139 51889 58195
rect 52013 58139 52069 58195
rect 52314 57753 52370 57755
rect 52314 57701 52316 57753
rect 52316 57701 52368 57753
rect 52368 57701 52370 57753
rect 52314 57699 52370 57701
rect 52525 57753 52581 57755
rect 52525 57701 52527 57753
rect 52527 57701 52579 57753
rect 52579 57701 52581 57753
rect 52525 57699 52581 57701
rect 52736 57753 52792 57755
rect 52736 57701 52738 57753
rect 52738 57701 52790 57753
rect 52790 57701 52792 57753
rect 52736 57699 52792 57701
rect 52946 57753 53002 57755
rect 52946 57701 52948 57753
rect 52948 57701 53000 57753
rect 53000 57701 53002 57753
rect 52946 57699 53002 57701
rect 53157 57753 53213 57755
rect 53157 57701 53159 57753
rect 53159 57701 53211 57753
rect 53211 57701 53213 57753
rect 53157 57699 53213 57701
rect 53369 57753 53425 57755
rect 53369 57701 53371 57753
rect 53371 57701 53423 57753
rect 53423 57701 53425 57753
rect 53369 57699 53425 57701
rect 53580 57753 53636 57755
rect 53580 57701 53582 57753
rect 53582 57701 53634 57753
rect 53634 57701 53636 57753
rect 53580 57699 53636 57701
rect 53790 57753 53846 57755
rect 53790 57701 53792 57753
rect 53792 57701 53844 57753
rect 53844 57701 53846 57753
rect 53790 57699 53846 57701
rect 54001 57753 54057 57755
rect 54001 57701 54003 57753
rect 54003 57701 54055 57753
rect 54055 57701 54057 57753
rect 54001 57699 54057 57701
rect 54212 57753 54268 57755
rect 54212 57701 54214 57753
rect 54214 57701 54266 57753
rect 54266 57701 54268 57753
rect 54212 57699 54268 57701
rect 51071 57259 51127 57315
rect 51251 57259 51307 57315
rect 51833 57259 51889 57315
rect 52013 57259 52069 57315
rect 50161 56853 50217 56855
rect 50161 56801 50190 56853
rect 50190 56801 50217 56853
rect 50161 56799 50217 56801
rect 50372 56799 50428 56855
rect 50584 56799 50640 56855
rect 50795 56799 50851 56855
rect 51071 56339 51127 56395
rect 51251 56339 51307 56395
rect 51833 56339 51889 56395
rect 52013 56339 52069 56395
rect 52314 55953 52370 55955
rect 52314 55901 52316 55953
rect 52316 55901 52368 55953
rect 52368 55901 52370 55953
rect 52314 55899 52370 55901
rect 52525 55953 52581 55955
rect 52525 55901 52527 55953
rect 52527 55901 52579 55953
rect 52579 55901 52581 55953
rect 52525 55899 52581 55901
rect 52736 55953 52792 55955
rect 52736 55901 52738 55953
rect 52738 55901 52790 55953
rect 52790 55901 52792 55953
rect 52736 55899 52792 55901
rect 52946 55953 53002 55955
rect 52946 55901 52948 55953
rect 52948 55901 53000 55953
rect 53000 55901 53002 55953
rect 52946 55899 53002 55901
rect 53157 55953 53213 55955
rect 53157 55901 53159 55953
rect 53159 55901 53211 55953
rect 53211 55901 53213 55953
rect 53157 55899 53213 55901
rect 53369 55953 53425 55955
rect 53369 55901 53371 55953
rect 53371 55901 53423 55953
rect 53423 55901 53425 55953
rect 53369 55899 53425 55901
rect 53580 55953 53636 55955
rect 53580 55901 53582 55953
rect 53582 55901 53634 55953
rect 53634 55901 53636 55953
rect 53580 55899 53636 55901
rect 53790 55953 53846 55955
rect 53790 55901 53792 55953
rect 53792 55901 53844 55953
rect 53844 55901 53846 55953
rect 53790 55899 53846 55901
rect 54001 55953 54057 55955
rect 54001 55901 54003 55953
rect 54003 55901 54055 55953
rect 54055 55901 54057 55953
rect 54001 55899 54057 55901
rect 54212 55953 54268 55955
rect 54212 55901 54214 55953
rect 54214 55901 54266 55953
rect 54266 55901 54268 55953
rect 54212 55899 54268 55901
rect 51071 55459 51127 55515
rect 51251 55459 51307 55515
rect 51833 55459 51889 55515
rect 52013 55459 52069 55515
rect 50161 55053 50217 55055
rect 50161 55001 50190 55053
rect 50190 55001 50217 55053
rect 50161 54999 50217 55001
rect 50372 54999 50428 55055
rect 50584 54999 50640 55055
rect 50795 54999 50851 55055
rect 51071 54539 51127 54595
rect 51251 54539 51307 54595
rect 51833 54539 51889 54595
rect 52013 54539 52069 54595
rect 52314 54153 52370 54155
rect 52314 54101 52316 54153
rect 52316 54101 52368 54153
rect 52368 54101 52370 54153
rect 52314 54099 52370 54101
rect 52525 54153 52581 54155
rect 52525 54101 52527 54153
rect 52527 54101 52579 54153
rect 52579 54101 52581 54153
rect 52525 54099 52581 54101
rect 52736 54153 52792 54155
rect 52736 54101 52738 54153
rect 52738 54101 52790 54153
rect 52790 54101 52792 54153
rect 52736 54099 52792 54101
rect 52946 54153 53002 54155
rect 52946 54101 52948 54153
rect 52948 54101 53000 54153
rect 53000 54101 53002 54153
rect 52946 54099 53002 54101
rect 53157 54153 53213 54155
rect 53157 54101 53159 54153
rect 53159 54101 53211 54153
rect 53211 54101 53213 54153
rect 53157 54099 53213 54101
rect 53369 54153 53425 54155
rect 53369 54101 53371 54153
rect 53371 54101 53423 54153
rect 53423 54101 53425 54153
rect 53369 54099 53425 54101
rect 53580 54153 53636 54155
rect 53580 54101 53582 54153
rect 53582 54101 53634 54153
rect 53634 54101 53636 54153
rect 53580 54099 53636 54101
rect 53790 54153 53846 54155
rect 53790 54101 53792 54153
rect 53792 54101 53844 54153
rect 53844 54101 53846 54153
rect 53790 54099 53846 54101
rect 54001 54153 54057 54155
rect 54001 54101 54003 54153
rect 54003 54101 54055 54153
rect 54055 54101 54057 54153
rect 54001 54099 54057 54101
rect 54212 54153 54268 54155
rect 54212 54101 54214 54153
rect 54214 54101 54266 54153
rect 54266 54101 54268 54153
rect 54212 54099 54268 54101
rect 51071 53659 51127 53715
rect 51251 53659 51307 53715
rect 51833 53659 51889 53715
rect 52013 53659 52069 53715
rect 50161 53253 50217 53255
rect 50161 53201 50190 53253
rect 50190 53201 50217 53253
rect 50161 53199 50217 53201
rect 50372 53199 50428 53255
rect 50584 53199 50640 53255
rect 50795 53199 50851 53255
rect 51071 52739 51127 52795
rect 51251 52739 51307 52795
rect 51833 52739 51889 52795
rect 52013 52739 52069 52795
rect 52314 52353 52370 52355
rect 52314 52301 52316 52353
rect 52316 52301 52368 52353
rect 52368 52301 52370 52353
rect 52314 52299 52370 52301
rect 52525 52353 52581 52355
rect 52525 52301 52527 52353
rect 52527 52301 52579 52353
rect 52579 52301 52581 52353
rect 52525 52299 52581 52301
rect 52736 52353 52792 52355
rect 52736 52301 52738 52353
rect 52738 52301 52790 52353
rect 52790 52301 52792 52353
rect 52736 52299 52792 52301
rect 52946 52353 53002 52355
rect 52946 52301 52948 52353
rect 52948 52301 53000 52353
rect 53000 52301 53002 52353
rect 52946 52299 53002 52301
rect 53157 52353 53213 52355
rect 53157 52301 53159 52353
rect 53159 52301 53211 52353
rect 53211 52301 53213 52353
rect 53157 52299 53213 52301
rect 53369 52353 53425 52355
rect 53369 52301 53371 52353
rect 53371 52301 53423 52353
rect 53423 52301 53425 52353
rect 53369 52299 53425 52301
rect 53580 52353 53636 52355
rect 53580 52301 53582 52353
rect 53582 52301 53634 52353
rect 53634 52301 53636 52353
rect 53580 52299 53636 52301
rect 53790 52353 53846 52355
rect 53790 52301 53792 52353
rect 53792 52301 53844 52353
rect 53844 52301 53846 52353
rect 53790 52299 53846 52301
rect 54001 52353 54057 52355
rect 54001 52301 54003 52353
rect 54003 52301 54055 52353
rect 54055 52301 54057 52353
rect 54001 52299 54057 52301
rect 54212 52353 54268 52355
rect 54212 52301 54214 52353
rect 54214 52301 54266 52353
rect 54266 52301 54268 52353
rect 54212 52299 54268 52301
rect 51071 51859 51127 51915
rect 51251 51859 51307 51915
rect 51833 51859 51889 51915
rect 52013 51859 52069 51915
rect 50161 51453 50217 51455
rect 50161 51401 50190 51453
rect 50190 51401 50217 51453
rect 50161 51399 50217 51401
rect 50372 51399 50428 51455
rect 50584 51399 50640 51455
rect 50795 51399 50851 51455
rect 51071 50939 51127 50995
rect 51251 50939 51307 50995
rect 51833 50939 51889 50995
rect 52013 50939 52069 50995
rect 52314 50553 52370 50555
rect 52314 50501 52316 50553
rect 52316 50501 52368 50553
rect 52368 50501 52370 50553
rect 52314 50499 52370 50501
rect 52525 50553 52581 50555
rect 52525 50501 52527 50553
rect 52527 50501 52579 50553
rect 52579 50501 52581 50553
rect 52525 50499 52581 50501
rect 52736 50553 52792 50555
rect 52736 50501 52738 50553
rect 52738 50501 52790 50553
rect 52790 50501 52792 50553
rect 52736 50499 52792 50501
rect 52946 50553 53002 50555
rect 52946 50501 52948 50553
rect 52948 50501 53000 50553
rect 53000 50501 53002 50553
rect 52946 50499 53002 50501
rect 53157 50553 53213 50555
rect 53157 50501 53159 50553
rect 53159 50501 53211 50553
rect 53211 50501 53213 50553
rect 53157 50499 53213 50501
rect 53369 50553 53425 50555
rect 53369 50501 53371 50553
rect 53371 50501 53423 50553
rect 53423 50501 53425 50553
rect 53369 50499 53425 50501
rect 53580 50553 53636 50555
rect 53580 50501 53582 50553
rect 53582 50501 53634 50553
rect 53634 50501 53636 50553
rect 53580 50499 53636 50501
rect 53790 50553 53846 50555
rect 53790 50501 53792 50553
rect 53792 50501 53844 50553
rect 53844 50501 53846 50553
rect 53790 50499 53846 50501
rect 54001 50553 54057 50555
rect 54001 50501 54003 50553
rect 54003 50501 54055 50553
rect 54055 50501 54057 50553
rect 54001 50499 54057 50501
rect 54212 50553 54268 50555
rect 54212 50501 54214 50553
rect 54214 50501 54266 50553
rect 54266 50501 54268 50553
rect 54212 50499 54268 50501
rect 51071 50059 51127 50115
rect 51251 50059 51307 50115
rect 51833 50059 51889 50115
rect 52013 50059 52069 50115
rect 50161 49653 50217 49655
rect 50161 49601 50190 49653
rect 50190 49601 50217 49653
rect 50161 49599 50217 49601
rect 50372 49599 50428 49655
rect 50584 49599 50640 49655
rect 50795 49599 50851 49655
rect 51071 49139 51127 49195
rect 51251 49139 51307 49195
rect 51833 49139 51889 49195
rect 52013 49139 52069 49195
rect 52314 48753 52370 48755
rect 52314 48701 52316 48753
rect 52316 48701 52368 48753
rect 52368 48701 52370 48753
rect 52314 48699 52370 48701
rect 52525 48753 52581 48755
rect 52525 48701 52527 48753
rect 52527 48701 52579 48753
rect 52579 48701 52581 48753
rect 52525 48699 52581 48701
rect 52736 48753 52792 48755
rect 52736 48701 52738 48753
rect 52738 48701 52790 48753
rect 52790 48701 52792 48753
rect 52736 48699 52792 48701
rect 52946 48753 53002 48755
rect 52946 48701 52948 48753
rect 52948 48701 53000 48753
rect 53000 48701 53002 48753
rect 52946 48699 53002 48701
rect 53157 48753 53213 48755
rect 53157 48701 53159 48753
rect 53159 48701 53211 48753
rect 53211 48701 53213 48753
rect 53157 48699 53213 48701
rect 53369 48753 53425 48755
rect 53369 48701 53371 48753
rect 53371 48701 53423 48753
rect 53423 48701 53425 48753
rect 53369 48699 53425 48701
rect 53580 48753 53636 48755
rect 53580 48701 53582 48753
rect 53582 48701 53634 48753
rect 53634 48701 53636 48753
rect 53580 48699 53636 48701
rect 53790 48753 53846 48755
rect 53790 48701 53792 48753
rect 53792 48701 53844 48753
rect 53844 48701 53846 48753
rect 53790 48699 53846 48701
rect 54001 48753 54057 48755
rect 54001 48701 54003 48753
rect 54003 48701 54055 48753
rect 54055 48701 54057 48753
rect 54001 48699 54057 48701
rect 54212 48753 54268 48755
rect 54212 48701 54214 48753
rect 54214 48701 54266 48753
rect 54266 48701 54268 48753
rect 54212 48699 54268 48701
rect 51071 48259 51127 48315
rect 51251 48259 51307 48315
rect 51833 48259 51889 48315
rect 52013 48259 52069 48315
rect 50161 47853 50217 47855
rect 50161 47801 50190 47853
rect 50190 47801 50217 47853
rect 50161 47799 50217 47801
rect 50372 47799 50428 47855
rect 50584 47799 50640 47855
rect 50795 47799 50851 47855
rect 51071 47339 51127 47395
rect 51251 47339 51307 47395
rect 51833 47339 51889 47395
rect 52013 47339 52069 47395
rect 52314 46953 52370 46955
rect 52314 46901 52316 46953
rect 52316 46901 52368 46953
rect 52368 46901 52370 46953
rect 52314 46899 52370 46901
rect 52525 46953 52581 46955
rect 52525 46901 52527 46953
rect 52527 46901 52579 46953
rect 52579 46901 52581 46953
rect 52525 46899 52581 46901
rect 52736 46953 52792 46955
rect 52736 46901 52738 46953
rect 52738 46901 52790 46953
rect 52790 46901 52792 46953
rect 52736 46899 52792 46901
rect 52946 46953 53002 46955
rect 52946 46901 52948 46953
rect 52948 46901 53000 46953
rect 53000 46901 53002 46953
rect 52946 46899 53002 46901
rect 53157 46953 53213 46955
rect 53157 46901 53159 46953
rect 53159 46901 53211 46953
rect 53211 46901 53213 46953
rect 53157 46899 53213 46901
rect 53369 46953 53425 46955
rect 53369 46901 53371 46953
rect 53371 46901 53423 46953
rect 53423 46901 53425 46953
rect 53369 46899 53425 46901
rect 53580 46953 53636 46955
rect 53580 46901 53582 46953
rect 53582 46901 53634 46953
rect 53634 46901 53636 46953
rect 53580 46899 53636 46901
rect 53790 46953 53846 46955
rect 53790 46901 53792 46953
rect 53792 46901 53844 46953
rect 53844 46901 53846 46953
rect 53790 46899 53846 46901
rect 54001 46953 54057 46955
rect 54001 46901 54003 46953
rect 54003 46901 54055 46953
rect 54055 46901 54057 46953
rect 54001 46899 54057 46901
rect 54212 46953 54268 46955
rect 54212 46901 54214 46953
rect 54214 46901 54266 46953
rect 54266 46901 54268 46953
rect 54212 46899 54268 46901
rect 51071 46459 51127 46515
rect 51251 46459 51307 46515
rect 51833 46459 51889 46515
rect 52013 46459 52069 46515
rect 50161 46053 50217 46055
rect 50161 46001 50190 46053
rect 50190 46001 50217 46053
rect 50161 45999 50217 46001
rect 50372 45999 50428 46055
rect 50584 45999 50640 46055
rect 50795 45999 50851 46055
rect 51071 45539 51127 45595
rect 51251 45539 51307 45595
rect 51833 45539 51889 45595
rect 52013 45539 52069 45595
rect 52314 45153 52370 45155
rect 52314 45101 52316 45153
rect 52316 45101 52368 45153
rect 52368 45101 52370 45153
rect 52314 45099 52370 45101
rect 52525 45153 52581 45155
rect 52525 45101 52527 45153
rect 52527 45101 52579 45153
rect 52579 45101 52581 45153
rect 52525 45099 52581 45101
rect 52736 45153 52792 45155
rect 52736 45101 52738 45153
rect 52738 45101 52790 45153
rect 52790 45101 52792 45153
rect 52736 45099 52792 45101
rect 52946 45153 53002 45155
rect 52946 45101 52948 45153
rect 52948 45101 53000 45153
rect 53000 45101 53002 45153
rect 52946 45099 53002 45101
rect 53157 45153 53213 45155
rect 53157 45101 53159 45153
rect 53159 45101 53211 45153
rect 53211 45101 53213 45153
rect 53157 45099 53213 45101
rect 53369 45153 53425 45155
rect 53369 45101 53371 45153
rect 53371 45101 53423 45153
rect 53423 45101 53425 45153
rect 53369 45099 53425 45101
rect 53580 45153 53636 45155
rect 53580 45101 53582 45153
rect 53582 45101 53634 45153
rect 53634 45101 53636 45153
rect 53580 45099 53636 45101
rect 53790 45153 53846 45155
rect 53790 45101 53792 45153
rect 53792 45101 53844 45153
rect 53844 45101 53846 45153
rect 53790 45099 53846 45101
rect 54001 45153 54057 45155
rect 54001 45101 54003 45153
rect 54003 45101 54055 45153
rect 54055 45101 54057 45153
rect 54001 45099 54057 45101
rect 54212 45153 54268 45155
rect 54212 45101 54214 45153
rect 54214 45101 54266 45153
rect 54266 45101 54268 45153
rect 54212 45099 54268 45101
rect 51071 44659 51127 44715
rect 51251 44659 51307 44715
rect 51833 44659 51889 44715
rect 52013 44659 52069 44715
rect 50161 44253 50217 44255
rect 50161 44201 50190 44253
rect 50190 44201 50217 44253
rect 50161 44199 50217 44201
rect 50372 44199 50428 44255
rect 50584 44199 50640 44255
rect 50795 44199 50851 44255
rect 51071 43739 51127 43795
rect 51251 43739 51307 43795
rect 51833 43739 51889 43795
rect 52013 43739 52069 43795
rect 52314 43353 52370 43355
rect 52314 43301 52316 43353
rect 52316 43301 52368 43353
rect 52368 43301 52370 43353
rect 52314 43299 52370 43301
rect 52525 43353 52581 43355
rect 52525 43301 52527 43353
rect 52527 43301 52579 43353
rect 52579 43301 52581 43353
rect 52525 43299 52581 43301
rect 52736 43353 52792 43355
rect 52736 43301 52738 43353
rect 52738 43301 52790 43353
rect 52790 43301 52792 43353
rect 52736 43299 52792 43301
rect 52946 43353 53002 43355
rect 52946 43301 52948 43353
rect 52948 43301 53000 43353
rect 53000 43301 53002 43353
rect 52946 43299 53002 43301
rect 53157 43353 53213 43355
rect 53157 43301 53159 43353
rect 53159 43301 53211 43353
rect 53211 43301 53213 43353
rect 53157 43299 53213 43301
rect 53369 43353 53425 43355
rect 53369 43301 53371 43353
rect 53371 43301 53423 43353
rect 53423 43301 53425 43353
rect 53369 43299 53425 43301
rect 53580 43353 53636 43355
rect 53580 43301 53582 43353
rect 53582 43301 53634 43353
rect 53634 43301 53636 43353
rect 53580 43299 53636 43301
rect 53790 43353 53846 43355
rect 53790 43301 53792 43353
rect 53792 43301 53844 43353
rect 53844 43301 53846 43353
rect 53790 43299 53846 43301
rect 54001 43353 54057 43355
rect 54001 43301 54003 43353
rect 54003 43301 54055 43353
rect 54055 43301 54057 43353
rect 54001 43299 54057 43301
rect 54212 43353 54268 43355
rect 54212 43301 54214 43353
rect 54214 43301 54266 43353
rect 54266 43301 54268 43353
rect 54212 43299 54268 43301
rect 51071 42859 51127 42915
rect 51251 42859 51307 42915
rect 51833 42859 51889 42915
rect 52013 42859 52069 42915
rect 50161 42453 50217 42455
rect 50161 42401 50190 42453
rect 50190 42401 50217 42453
rect 50161 42399 50217 42401
rect 50372 42399 50428 42455
rect 50584 42399 50640 42455
rect 50795 42399 50851 42455
rect 51071 41939 51127 41995
rect 51251 41939 51307 41995
rect 51833 41939 51889 41995
rect 52013 41939 52069 41995
rect 52314 41553 52370 41555
rect 52314 41501 52316 41553
rect 52316 41501 52368 41553
rect 52368 41501 52370 41553
rect 52314 41499 52370 41501
rect 52525 41553 52581 41555
rect 52525 41501 52527 41553
rect 52527 41501 52579 41553
rect 52579 41501 52581 41553
rect 52525 41499 52581 41501
rect 52736 41553 52792 41555
rect 52736 41501 52738 41553
rect 52738 41501 52790 41553
rect 52790 41501 52792 41553
rect 52736 41499 52792 41501
rect 52946 41553 53002 41555
rect 52946 41501 52948 41553
rect 52948 41501 53000 41553
rect 53000 41501 53002 41553
rect 52946 41499 53002 41501
rect 53157 41553 53213 41555
rect 53157 41501 53159 41553
rect 53159 41501 53211 41553
rect 53211 41501 53213 41553
rect 53157 41499 53213 41501
rect 53369 41553 53425 41555
rect 53369 41501 53371 41553
rect 53371 41501 53423 41553
rect 53423 41501 53425 41553
rect 53369 41499 53425 41501
rect 53580 41553 53636 41555
rect 53580 41501 53582 41553
rect 53582 41501 53634 41553
rect 53634 41501 53636 41553
rect 53580 41499 53636 41501
rect 53790 41553 53846 41555
rect 53790 41501 53792 41553
rect 53792 41501 53844 41553
rect 53844 41501 53846 41553
rect 53790 41499 53846 41501
rect 54001 41553 54057 41555
rect 54001 41501 54003 41553
rect 54003 41501 54055 41553
rect 54055 41501 54057 41553
rect 54001 41499 54057 41501
rect 54212 41553 54268 41555
rect 54212 41501 54214 41553
rect 54214 41501 54266 41553
rect 54266 41501 54268 41553
rect 54212 41499 54268 41501
rect 51071 41059 51127 41115
rect 51251 41059 51307 41115
rect 51833 41059 51889 41115
rect 52013 41059 52069 41115
rect 50161 40653 50217 40655
rect 50161 40601 50190 40653
rect 50190 40601 50217 40653
rect 50161 40599 50217 40601
rect 50372 40599 50428 40655
rect 50584 40599 50640 40655
rect 50795 40599 50851 40655
rect 51071 40139 51127 40195
rect 51251 40139 51307 40195
rect 51833 40139 51889 40195
rect 52013 40139 52069 40195
rect 52314 39753 52370 39755
rect 52314 39701 52316 39753
rect 52316 39701 52368 39753
rect 52368 39701 52370 39753
rect 52314 39699 52370 39701
rect 52525 39753 52581 39755
rect 52525 39701 52527 39753
rect 52527 39701 52579 39753
rect 52579 39701 52581 39753
rect 52525 39699 52581 39701
rect 52736 39753 52792 39755
rect 52736 39701 52738 39753
rect 52738 39701 52790 39753
rect 52790 39701 52792 39753
rect 52736 39699 52792 39701
rect 52946 39753 53002 39755
rect 52946 39701 52948 39753
rect 52948 39701 53000 39753
rect 53000 39701 53002 39753
rect 52946 39699 53002 39701
rect 53157 39753 53213 39755
rect 53157 39701 53159 39753
rect 53159 39701 53211 39753
rect 53211 39701 53213 39753
rect 53157 39699 53213 39701
rect 53369 39753 53425 39755
rect 53369 39701 53371 39753
rect 53371 39701 53423 39753
rect 53423 39701 53425 39753
rect 53369 39699 53425 39701
rect 53580 39753 53636 39755
rect 53580 39701 53582 39753
rect 53582 39701 53634 39753
rect 53634 39701 53636 39753
rect 53580 39699 53636 39701
rect 53790 39753 53846 39755
rect 53790 39701 53792 39753
rect 53792 39701 53844 39753
rect 53844 39701 53846 39753
rect 53790 39699 53846 39701
rect 54001 39753 54057 39755
rect 54001 39701 54003 39753
rect 54003 39701 54055 39753
rect 54055 39701 54057 39753
rect 54001 39699 54057 39701
rect 54212 39753 54268 39755
rect 54212 39701 54214 39753
rect 54214 39701 54266 39753
rect 54266 39701 54268 39753
rect 54212 39699 54268 39701
rect 51071 39259 51127 39315
rect 51251 39259 51307 39315
rect 51833 39259 51889 39315
rect 52013 39259 52069 39315
rect 50161 38853 50217 38855
rect 50161 38801 50190 38853
rect 50190 38801 50217 38853
rect 50161 38799 50217 38801
rect 50372 38799 50428 38855
rect 50584 38799 50640 38855
rect 50795 38799 50851 38855
rect 51071 38339 51127 38395
rect 51251 38339 51307 38395
rect 51833 38339 51889 38395
rect 52013 38339 52069 38395
rect 52314 37953 52370 37955
rect 52314 37901 52316 37953
rect 52316 37901 52368 37953
rect 52368 37901 52370 37953
rect 52314 37899 52370 37901
rect 52525 37953 52581 37955
rect 52525 37901 52527 37953
rect 52527 37901 52579 37953
rect 52579 37901 52581 37953
rect 52525 37899 52581 37901
rect 52736 37953 52792 37955
rect 52736 37901 52738 37953
rect 52738 37901 52790 37953
rect 52790 37901 52792 37953
rect 52736 37899 52792 37901
rect 52946 37953 53002 37955
rect 52946 37901 52948 37953
rect 52948 37901 53000 37953
rect 53000 37901 53002 37953
rect 52946 37899 53002 37901
rect 53157 37953 53213 37955
rect 53157 37901 53159 37953
rect 53159 37901 53211 37953
rect 53211 37901 53213 37953
rect 53157 37899 53213 37901
rect 53369 37953 53425 37955
rect 53369 37901 53371 37953
rect 53371 37901 53423 37953
rect 53423 37901 53425 37953
rect 53369 37899 53425 37901
rect 53580 37953 53636 37955
rect 53580 37901 53582 37953
rect 53582 37901 53634 37953
rect 53634 37901 53636 37953
rect 53580 37899 53636 37901
rect 53790 37953 53846 37955
rect 53790 37901 53792 37953
rect 53792 37901 53844 37953
rect 53844 37901 53846 37953
rect 53790 37899 53846 37901
rect 54001 37953 54057 37955
rect 54001 37901 54003 37953
rect 54003 37901 54055 37953
rect 54055 37901 54057 37953
rect 54001 37899 54057 37901
rect 54212 37953 54268 37955
rect 54212 37901 54214 37953
rect 54214 37901 54266 37953
rect 54266 37901 54268 37953
rect 54212 37899 54268 37901
rect 51071 37459 51127 37515
rect 51251 37459 51307 37515
rect 51833 37459 51889 37515
rect 52013 37459 52069 37515
rect 50161 37053 50217 37055
rect 50161 37001 50190 37053
rect 50190 37001 50217 37053
rect 50161 36999 50217 37001
rect 50372 36999 50428 37055
rect 50584 36999 50640 37055
rect 50795 36999 50851 37055
rect 51071 36539 51127 36595
rect 51251 36539 51307 36595
rect 51833 36539 51889 36595
rect 52013 36539 52069 36595
rect 52314 36153 52370 36155
rect 52314 36101 52316 36153
rect 52316 36101 52368 36153
rect 52368 36101 52370 36153
rect 52314 36099 52370 36101
rect 52525 36153 52581 36155
rect 52525 36101 52527 36153
rect 52527 36101 52579 36153
rect 52579 36101 52581 36153
rect 52525 36099 52581 36101
rect 52736 36153 52792 36155
rect 52736 36101 52738 36153
rect 52738 36101 52790 36153
rect 52790 36101 52792 36153
rect 52736 36099 52792 36101
rect 52946 36153 53002 36155
rect 52946 36101 52948 36153
rect 52948 36101 53000 36153
rect 53000 36101 53002 36153
rect 52946 36099 53002 36101
rect 53157 36153 53213 36155
rect 53157 36101 53159 36153
rect 53159 36101 53211 36153
rect 53211 36101 53213 36153
rect 53157 36099 53213 36101
rect 53369 36153 53425 36155
rect 53369 36101 53371 36153
rect 53371 36101 53423 36153
rect 53423 36101 53425 36153
rect 53369 36099 53425 36101
rect 53580 36153 53636 36155
rect 53580 36101 53582 36153
rect 53582 36101 53634 36153
rect 53634 36101 53636 36153
rect 53580 36099 53636 36101
rect 53790 36153 53846 36155
rect 53790 36101 53792 36153
rect 53792 36101 53844 36153
rect 53844 36101 53846 36153
rect 53790 36099 53846 36101
rect 54001 36153 54057 36155
rect 54001 36101 54003 36153
rect 54003 36101 54055 36153
rect 54055 36101 54057 36153
rect 54001 36099 54057 36101
rect 54212 36153 54268 36155
rect 54212 36101 54214 36153
rect 54214 36101 54266 36153
rect 54266 36101 54268 36153
rect 54212 36099 54268 36101
rect 56013 65853 56069 65855
rect 56013 65801 56015 65853
rect 56015 65801 56067 65853
rect 56067 65801 56069 65853
rect 56013 65799 56069 65801
rect 56224 65853 56280 65855
rect 56224 65801 56226 65853
rect 56226 65801 56278 65853
rect 56278 65801 56280 65853
rect 56224 65799 56280 65801
rect 56435 65853 56491 65855
rect 56435 65801 56437 65853
rect 56437 65801 56489 65853
rect 56489 65801 56491 65853
rect 56435 65799 56491 65801
rect 56646 65853 56702 65855
rect 56646 65801 56648 65853
rect 56648 65801 56700 65853
rect 56700 65801 56702 65853
rect 56646 65799 56702 65801
rect 56857 65853 56913 65855
rect 56857 65801 56859 65853
rect 56859 65801 56911 65853
rect 56911 65801 56913 65853
rect 56857 65799 56913 65801
rect 57068 65853 57124 65855
rect 57068 65801 57070 65853
rect 57070 65801 57122 65853
rect 57122 65801 57124 65853
rect 57068 65799 57124 65801
rect 57279 65853 57335 65855
rect 57279 65801 57281 65853
rect 57281 65801 57333 65853
rect 57333 65801 57335 65853
rect 57279 65799 57335 65801
rect 54853 64953 54909 64955
rect 54853 64901 54855 64953
rect 54855 64901 54907 64953
rect 54907 64901 54909 64953
rect 54853 64899 54909 64901
rect 55064 64953 55120 64955
rect 55064 64901 55066 64953
rect 55066 64901 55118 64953
rect 55118 64901 55120 64953
rect 55064 64899 55120 64901
rect 55276 64953 55332 64955
rect 55276 64901 55278 64953
rect 55278 64901 55330 64953
rect 55330 64901 55332 64953
rect 55276 64899 55332 64901
rect 55487 64953 55543 64955
rect 55487 64901 55489 64953
rect 55489 64901 55541 64953
rect 55541 64901 55543 64953
rect 55487 64899 55543 64901
rect 56013 64053 56069 64055
rect 56013 64001 56015 64053
rect 56015 64001 56067 64053
rect 56067 64001 56069 64053
rect 56013 63999 56069 64001
rect 56224 64053 56280 64055
rect 56224 64001 56226 64053
rect 56226 64001 56278 64053
rect 56278 64001 56280 64053
rect 56224 63999 56280 64001
rect 56435 64053 56491 64055
rect 56435 64001 56437 64053
rect 56437 64001 56489 64053
rect 56489 64001 56491 64053
rect 56435 63999 56491 64001
rect 56646 64053 56702 64055
rect 56646 64001 56648 64053
rect 56648 64001 56700 64053
rect 56700 64001 56702 64053
rect 56646 63999 56702 64001
rect 56857 64053 56913 64055
rect 56857 64001 56859 64053
rect 56859 64001 56911 64053
rect 56911 64001 56913 64053
rect 56857 63999 56913 64001
rect 57068 64053 57124 64055
rect 57068 64001 57070 64053
rect 57070 64001 57122 64053
rect 57122 64001 57124 64053
rect 57068 63999 57124 64001
rect 57279 64053 57335 64055
rect 57279 64001 57281 64053
rect 57281 64001 57333 64053
rect 57333 64001 57335 64053
rect 57279 63999 57335 64001
rect 54853 63153 54909 63155
rect 54853 63101 54855 63153
rect 54855 63101 54907 63153
rect 54907 63101 54909 63153
rect 54853 63099 54909 63101
rect 55064 63153 55120 63155
rect 55064 63101 55066 63153
rect 55066 63101 55118 63153
rect 55118 63101 55120 63153
rect 55064 63099 55120 63101
rect 55276 63153 55332 63155
rect 55276 63101 55278 63153
rect 55278 63101 55330 63153
rect 55330 63101 55332 63153
rect 55276 63099 55332 63101
rect 55487 63153 55543 63155
rect 55487 63101 55489 63153
rect 55489 63101 55541 63153
rect 55541 63101 55543 63153
rect 55487 63099 55543 63101
rect 56013 62253 56069 62255
rect 56013 62201 56015 62253
rect 56015 62201 56067 62253
rect 56067 62201 56069 62253
rect 56013 62199 56069 62201
rect 56224 62253 56280 62255
rect 56224 62201 56226 62253
rect 56226 62201 56278 62253
rect 56278 62201 56280 62253
rect 56224 62199 56280 62201
rect 56435 62253 56491 62255
rect 56435 62201 56437 62253
rect 56437 62201 56489 62253
rect 56489 62201 56491 62253
rect 56435 62199 56491 62201
rect 56646 62253 56702 62255
rect 56646 62201 56648 62253
rect 56648 62201 56700 62253
rect 56700 62201 56702 62253
rect 56646 62199 56702 62201
rect 56857 62253 56913 62255
rect 56857 62201 56859 62253
rect 56859 62201 56911 62253
rect 56911 62201 56913 62253
rect 56857 62199 56913 62201
rect 57068 62253 57124 62255
rect 57068 62201 57070 62253
rect 57070 62201 57122 62253
rect 57122 62201 57124 62253
rect 57068 62199 57124 62201
rect 57279 62253 57335 62255
rect 57279 62201 57281 62253
rect 57281 62201 57333 62253
rect 57333 62201 57335 62253
rect 57279 62199 57335 62201
rect 54853 61353 54909 61355
rect 54853 61301 54855 61353
rect 54855 61301 54907 61353
rect 54907 61301 54909 61353
rect 54853 61299 54909 61301
rect 55064 61353 55120 61355
rect 55064 61301 55066 61353
rect 55066 61301 55118 61353
rect 55118 61301 55120 61353
rect 55064 61299 55120 61301
rect 55276 61353 55332 61355
rect 55276 61301 55278 61353
rect 55278 61301 55330 61353
rect 55330 61301 55332 61353
rect 55276 61299 55332 61301
rect 55487 61353 55543 61355
rect 55487 61301 55489 61353
rect 55489 61301 55541 61353
rect 55541 61301 55543 61353
rect 55487 61299 55543 61301
rect 56013 60453 56069 60455
rect 56013 60401 56015 60453
rect 56015 60401 56067 60453
rect 56067 60401 56069 60453
rect 56013 60399 56069 60401
rect 56224 60453 56280 60455
rect 56224 60401 56226 60453
rect 56226 60401 56278 60453
rect 56278 60401 56280 60453
rect 56224 60399 56280 60401
rect 56435 60453 56491 60455
rect 56435 60401 56437 60453
rect 56437 60401 56489 60453
rect 56489 60401 56491 60453
rect 56435 60399 56491 60401
rect 56646 60453 56702 60455
rect 56646 60401 56648 60453
rect 56648 60401 56700 60453
rect 56700 60401 56702 60453
rect 56646 60399 56702 60401
rect 56857 60453 56913 60455
rect 56857 60401 56859 60453
rect 56859 60401 56911 60453
rect 56911 60401 56913 60453
rect 56857 60399 56913 60401
rect 57068 60453 57124 60455
rect 57068 60401 57070 60453
rect 57070 60401 57122 60453
rect 57122 60401 57124 60453
rect 57068 60399 57124 60401
rect 57279 60453 57335 60455
rect 57279 60401 57281 60453
rect 57281 60401 57333 60453
rect 57333 60401 57335 60453
rect 57279 60399 57335 60401
rect 54853 59553 54909 59555
rect 54853 59501 54855 59553
rect 54855 59501 54907 59553
rect 54907 59501 54909 59553
rect 54853 59499 54909 59501
rect 55064 59553 55120 59555
rect 55064 59501 55066 59553
rect 55066 59501 55118 59553
rect 55118 59501 55120 59553
rect 55064 59499 55120 59501
rect 55276 59553 55332 59555
rect 55276 59501 55278 59553
rect 55278 59501 55330 59553
rect 55330 59501 55332 59553
rect 55276 59499 55332 59501
rect 55487 59553 55543 59555
rect 55487 59501 55489 59553
rect 55489 59501 55541 59553
rect 55541 59501 55543 59553
rect 55487 59499 55543 59501
rect 56013 58653 56069 58655
rect 56013 58601 56015 58653
rect 56015 58601 56067 58653
rect 56067 58601 56069 58653
rect 56013 58599 56069 58601
rect 56224 58653 56280 58655
rect 56224 58601 56226 58653
rect 56226 58601 56278 58653
rect 56278 58601 56280 58653
rect 56224 58599 56280 58601
rect 56435 58653 56491 58655
rect 56435 58601 56437 58653
rect 56437 58601 56489 58653
rect 56489 58601 56491 58653
rect 56435 58599 56491 58601
rect 56646 58653 56702 58655
rect 56646 58601 56648 58653
rect 56648 58601 56700 58653
rect 56700 58601 56702 58653
rect 56646 58599 56702 58601
rect 56857 58653 56913 58655
rect 56857 58601 56859 58653
rect 56859 58601 56911 58653
rect 56911 58601 56913 58653
rect 56857 58599 56913 58601
rect 57068 58653 57124 58655
rect 57068 58601 57070 58653
rect 57070 58601 57122 58653
rect 57122 58601 57124 58653
rect 57068 58599 57124 58601
rect 57279 58653 57335 58655
rect 57279 58601 57281 58653
rect 57281 58601 57333 58653
rect 57333 58601 57335 58653
rect 57279 58599 57335 58601
rect 54853 57753 54909 57755
rect 54853 57701 54855 57753
rect 54855 57701 54907 57753
rect 54907 57701 54909 57753
rect 54853 57699 54909 57701
rect 55064 57753 55120 57755
rect 55064 57701 55066 57753
rect 55066 57701 55118 57753
rect 55118 57701 55120 57753
rect 55064 57699 55120 57701
rect 55276 57753 55332 57755
rect 55276 57701 55278 57753
rect 55278 57701 55330 57753
rect 55330 57701 55332 57753
rect 55276 57699 55332 57701
rect 55487 57753 55543 57755
rect 55487 57701 55489 57753
rect 55489 57701 55541 57753
rect 55541 57701 55543 57753
rect 55487 57699 55543 57701
rect 56013 56853 56069 56855
rect 56013 56801 56015 56853
rect 56015 56801 56067 56853
rect 56067 56801 56069 56853
rect 56013 56799 56069 56801
rect 56224 56853 56280 56855
rect 56224 56801 56226 56853
rect 56226 56801 56278 56853
rect 56278 56801 56280 56853
rect 56224 56799 56280 56801
rect 56435 56853 56491 56855
rect 56435 56801 56437 56853
rect 56437 56801 56489 56853
rect 56489 56801 56491 56853
rect 56435 56799 56491 56801
rect 56646 56853 56702 56855
rect 56646 56801 56648 56853
rect 56648 56801 56700 56853
rect 56700 56801 56702 56853
rect 56646 56799 56702 56801
rect 56857 56853 56913 56855
rect 56857 56801 56859 56853
rect 56859 56801 56911 56853
rect 56911 56801 56913 56853
rect 56857 56799 56913 56801
rect 57068 56853 57124 56855
rect 57068 56801 57070 56853
rect 57070 56801 57122 56853
rect 57122 56801 57124 56853
rect 57068 56799 57124 56801
rect 57279 56853 57335 56855
rect 57279 56801 57281 56853
rect 57281 56801 57333 56853
rect 57333 56801 57335 56853
rect 57279 56799 57335 56801
rect 54853 55953 54909 55955
rect 54853 55901 54855 55953
rect 54855 55901 54907 55953
rect 54907 55901 54909 55953
rect 54853 55899 54909 55901
rect 55064 55953 55120 55955
rect 55064 55901 55066 55953
rect 55066 55901 55118 55953
rect 55118 55901 55120 55953
rect 55064 55899 55120 55901
rect 55276 55953 55332 55955
rect 55276 55901 55278 55953
rect 55278 55901 55330 55953
rect 55330 55901 55332 55953
rect 55276 55899 55332 55901
rect 55487 55953 55543 55955
rect 55487 55901 55489 55953
rect 55489 55901 55541 55953
rect 55541 55901 55543 55953
rect 55487 55899 55543 55901
rect 56013 55053 56069 55055
rect 56013 55001 56015 55053
rect 56015 55001 56067 55053
rect 56067 55001 56069 55053
rect 56013 54999 56069 55001
rect 56224 55053 56280 55055
rect 56224 55001 56226 55053
rect 56226 55001 56278 55053
rect 56278 55001 56280 55053
rect 56224 54999 56280 55001
rect 56435 55053 56491 55055
rect 56435 55001 56437 55053
rect 56437 55001 56489 55053
rect 56489 55001 56491 55053
rect 56435 54999 56491 55001
rect 56646 55053 56702 55055
rect 56646 55001 56648 55053
rect 56648 55001 56700 55053
rect 56700 55001 56702 55053
rect 56646 54999 56702 55001
rect 56857 55053 56913 55055
rect 56857 55001 56859 55053
rect 56859 55001 56911 55053
rect 56911 55001 56913 55053
rect 56857 54999 56913 55001
rect 57068 55053 57124 55055
rect 57068 55001 57070 55053
rect 57070 55001 57122 55053
rect 57122 55001 57124 55053
rect 57068 54999 57124 55001
rect 57279 55053 57335 55055
rect 57279 55001 57281 55053
rect 57281 55001 57333 55053
rect 57333 55001 57335 55053
rect 57279 54999 57335 55001
rect 54853 54153 54909 54155
rect 54853 54101 54855 54153
rect 54855 54101 54907 54153
rect 54907 54101 54909 54153
rect 54853 54099 54909 54101
rect 55064 54153 55120 54155
rect 55064 54101 55066 54153
rect 55066 54101 55118 54153
rect 55118 54101 55120 54153
rect 55064 54099 55120 54101
rect 55276 54153 55332 54155
rect 55276 54101 55278 54153
rect 55278 54101 55330 54153
rect 55330 54101 55332 54153
rect 55276 54099 55332 54101
rect 55487 54153 55543 54155
rect 55487 54101 55489 54153
rect 55489 54101 55541 54153
rect 55541 54101 55543 54153
rect 55487 54099 55543 54101
rect 56013 53253 56069 53255
rect 56013 53201 56015 53253
rect 56015 53201 56067 53253
rect 56067 53201 56069 53253
rect 56013 53199 56069 53201
rect 56224 53253 56280 53255
rect 56224 53201 56226 53253
rect 56226 53201 56278 53253
rect 56278 53201 56280 53253
rect 56224 53199 56280 53201
rect 56435 53253 56491 53255
rect 56435 53201 56437 53253
rect 56437 53201 56489 53253
rect 56489 53201 56491 53253
rect 56435 53199 56491 53201
rect 56646 53253 56702 53255
rect 56646 53201 56648 53253
rect 56648 53201 56700 53253
rect 56700 53201 56702 53253
rect 56646 53199 56702 53201
rect 56857 53253 56913 53255
rect 56857 53201 56859 53253
rect 56859 53201 56911 53253
rect 56911 53201 56913 53253
rect 56857 53199 56913 53201
rect 57068 53253 57124 53255
rect 57068 53201 57070 53253
rect 57070 53201 57122 53253
rect 57122 53201 57124 53253
rect 57068 53199 57124 53201
rect 57279 53253 57335 53255
rect 57279 53201 57281 53253
rect 57281 53201 57333 53253
rect 57333 53201 57335 53253
rect 57279 53199 57335 53201
rect 54853 52353 54909 52355
rect 54853 52301 54855 52353
rect 54855 52301 54907 52353
rect 54907 52301 54909 52353
rect 54853 52299 54909 52301
rect 55064 52353 55120 52355
rect 55064 52301 55066 52353
rect 55066 52301 55118 52353
rect 55118 52301 55120 52353
rect 55064 52299 55120 52301
rect 55276 52353 55332 52355
rect 55276 52301 55278 52353
rect 55278 52301 55330 52353
rect 55330 52301 55332 52353
rect 55276 52299 55332 52301
rect 55487 52353 55543 52355
rect 55487 52301 55489 52353
rect 55489 52301 55541 52353
rect 55541 52301 55543 52353
rect 55487 52299 55543 52301
rect 56013 51453 56069 51455
rect 56013 51401 56015 51453
rect 56015 51401 56067 51453
rect 56067 51401 56069 51453
rect 56013 51399 56069 51401
rect 56224 51453 56280 51455
rect 56224 51401 56226 51453
rect 56226 51401 56278 51453
rect 56278 51401 56280 51453
rect 56224 51399 56280 51401
rect 56435 51453 56491 51455
rect 56435 51401 56437 51453
rect 56437 51401 56489 51453
rect 56489 51401 56491 51453
rect 56435 51399 56491 51401
rect 56646 51453 56702 51455
rect 56646 51401 56648 51453
rect 56648 51401 56700 51453
rect 56700 51401 56702 51453
rect 56646 51399 56702 51401
rect 56857 51453 56913 51455
rect 56857 51401 56859 51453
rect 56859 51401 56911 51453
rect 56911 51401 56913 51453
rect 56857 51399 56913 51401
rect 57068 51453 57124 51455
rect 57068 51401 57070 51453
rect 57070 51401 57122 51453
rect 57122 51401 57124 51453
rect 57068 51399 57124 51401
rect 57279 51453 57335 51455
rect 57279 51401 57281 51453
rect 57281 51401 57333 51453
rect 57333 51401 57335 51453
rect 57279 51399 57335 51401
rect 54853 50553 54909 50555
rect 54853 50501 54855 50553
rect 54855 50501 54907 50553
rect 54907 50501 54909 50553
rect 54853 50499 54909 50501
rect 55064 50553 55120 50555
rect 55064 50501 55066 50553
rect 55066 50501 55118 50553
rect 55118 50501 55120 50553
rect 55064 50499 55120 50501
rect 55276 50553 55332 50555
rect 55276 50501 55278 50553
rect 55278 50501 55330 50553
rect 55330 50501 55332 50553
rect 55276 50499 55332 50501
rect 55487 50553 55543 50555
rect 55487 50501 55489 50553
rect 55489 50501 55541 50553
rect 55541 50501 55543 50553
rect 55487 50499 55543 50501
rect 56013 49653 56069 49655
rect 56013 49601 56015 49653
rect 56015 49601 56067 49653
rect 56067 49601 56069 49653
rect 56013 49599 56069 49601
rect 56224 49653 56280 49655
rect 56224 49601 56226 49653
rect 56226 49601 56278 49653
rect 56278 49601 56280 49653
rect 56224 49599 56280 49601
rect 56435 49653 56491 49655
rect 56435 49601 56437 49653
rect 56437 49601 56489 49653
rect 56489 49601 56491 49653
rect 56435 49599 56491 49601
rect 56646 49653 56702 49655
rect 56646 49601 56648 49653
rect 56648 49601 56700 49653
rect 56700 49601 56702 49653
rect 56646 49599 56702 49601
rect 56857 49653 56913 49655
rect 56857 49601 56859 49653
rect 56859 49601 56911 49653
rect 56911 49601 56913 49653
rect 56857 49599 56913 49601
rect 57068 49653 57124 49655
rect 57068 49601 57070 49653
rect 57070 49601 57122 49653
rect 57122 49601 57124 49653
rect 57068 49599 57124 49601
rect 57279 49653 57335 49655
rect 57279 49601 57281 49653
rect 57281 49601 57333 49653
rect 57333 49601 57335 49653
rect 57279 49599 57335 49601
rect 54853 48753 54909 48755
rect 54853 48701 54855 48753
rect 54855 48701 54907 48753
rect 54907 48701 54909 48753
rect 54853 48699 54909 48701
rect 55064 48753 55120 48755
rect 55064 48701 55066 48753
rect 55066 48701 55118 48753
rect 55118 48701 55120 48753
rect 55064 48699 55120 48701
rect 55276 48753 55332 48755
rect 55276 48701 55278 48753
rect 55278 48701 55330 48753
rect 55330 48701 55332 48753
rect 55276 48699 55332 48701
rect 55487 48753 55543 48755
rect 55487 48701 55489 48753
rect 55489 48701 55541 48753
rect 55541 48701 55543 48753
rect 55487 48699 55543 48701
rect 56013 47853 56069 47855
rect 56013 47801 56015 47853
rect 56015 47801 56067 47853
rect 56067 47801 56069 47853
rect 56013 47799 56069 47801
rect 56224 47853 56280 47855
rect 56224 47801 56226 47853
rect 56226 47801 56278 47853
rect 56278 47801 56280 47853
rect 56224 47799 56280 47801
rect 56435 47853 56491 47855
rect 56435 47801 56437 47853
rect 56437 47801 56489 47853
rect 56489 47801 56491 47853
rect 56435 47799 56491 47801
rect 56646 47853 56702 47855
rect 56646 47801 56648 47853
rect 56648 47801 56700 47853
rect 56700 47801 56702 47853
rect 56646 47799 56702 47801
rect 56857 47853 56913 47855
rect 56857 47801 56859 47853
rect 56859 47801 56911 47853
rect 56911 47801 56913 47853
rect 56857 47799 56913 47801
rect 57068 47853 57124 47855
rect 57068 47801 57070 47853
rect 57070 47801 57122 47853
rect 57122 47801 57124 47853
rect 57068 47799 57124 47801
rect 57279 47853 57335 47855
rect 57279 47801 57281 47853
rect 57281 47801 57333 47853
rect 57333 47801 57335 47853
rect 57279 47799 57335 47801
rect 54853 46953 54909 46955
rect 54853 46901 54855 46953
rect 54855 46901 54907 46953
rect 54907 46901 54909 46953
rect 54853 46899 54909 46901
rect 55064 46953 55120 46955
rect 55064 46901 55066 46953
rect 55066 46901 55118 46953
rect 55118 46901 55120 46953
rect 55064 46899 55120 46901
rect 55276 46953 55332 46955
rect 55276 46901 55278 46953
rect 55278 46901 55330 46953
rect 55330 46901 55332 46953
rect 55276 46899 55332 46901
rect 55487 46953 55543 46955
rect 55487 46901 55489 46953
rect 55489 46901 55541 46953
rect 55541 46901 55543 46953
rect 55487 46899 55543 46901
rect 56013 46053 56069 46055
rect 56013 46001 56015 46053
rect 56015 46001 56067 46053
rect 56067 46001 56069 46053
rect 56013 45999 56069 46001
rect 56224 46053 56280 46055
rect 56224 46001 56226 46053
rect 56226 46001 56278 46053
rect 56278 46001 56280 46053
rect 56224 45999 56280 46001
rect 56435 46053 56491 46055
rect 56435 46001 56437 46053
rect 56437 46001 56489 46053
rect 56489 46001 56491 46053
rect 56435 45999 56491 46001
rect 56646 46053 56702 46055
rect 56646 46001 56648 46053
rect 56648 46001 56700 46053
rect 56700 46001 56702 46053
rect 56646 45999 56702 46001
rect 56857 46053 56913 46055
rect 56857 46001 56859 46053
rect 56859 46001 56911 46053
rect 56911 46001 56913 46053
rect 56857 45999 56913 46001
rect 57068 46053 57124 46055
rect 57068 46001 57070 46053
rect 57070 46001 57122 46053
rect 57122 46001 57124 46053
rect 57068 45999 57124 46001
rect 57279 46053 57335 46055
rect 57279 46001 57281 46053
rect 57281 46001 57333 46053
rect 57333 46001 57335 46053
rect 57279 45999 57335 46001
rect 54853 45153 54909 45155
rect 54853 45101 54855 45153
rect 54855 45101 54907 45153
rect 54907 45101 54909 45153
rect 54853 45099 54909 45101
rect 55064 45153 55120 45155
rect 55064 45101 55066 45153
rect 55066 45101 55118 45153
rect 55118 45101 55120 45153
rect 55064 45099 55120 45101
rect 55276 45153 55332 45155
rect 55276 45101 55278 45153
rect 55278 45101 55330 45153
rect 55330 45101 55332 45153
rect 55276 45099 55332 45101
rect 55487 45153 55543 45155
rect 55487 45101 55489 45153
rect 55489 45101 55541 45153
rect 55541 45101 55543 45153
rect 55487 45099 55543 45101
rect 56013 44253 56069 44255
rect 56013 44201 56015 44253
rect 56015 44201 56067 44253
rect 56067 44201 56069 44253
rect 56013 44199 56069 44201
rect 56224 44253 56280 44255
rect 56224 44201 56226 44253
rect 56226 44201 56278 44253
rect 56278 44201 56280 44253
rect 56224 44199 56280 44201
rect 56435 44253 56491 44255
rect 56435 44201 56437 44253
rect 56437 44201 56489 44253
rect 56489 44201 56491 44253
rect 56435 44199 56491 44201
rect 56646 44253 56702 44255
rect 56646 44201 56648 44253
rect 56648 44201 56700 44253
rect 56700 44201 56702 44253
rect 56646 44199 56702 44201
rect 56857 44253 56913 44255
rect 56857 44201 56859 44253
rect 56859 44201 56911 44253
rect 56911 44201 56913 44253
rect 56857 44199 56913 44201
rect 57068 44253 57124 44255
rect 57068 44201 57070 44253
rect 57070 44201 57122 44253
rect 57122 44201 57124 44253
rect 57068 44199 57124 44201
rect 57279 44253 57335 44255
rect 57279 44201 57281 44253
rect 57281 44201 57333 44253
rect 57333 44201 57335 44253
rect 57279 44199 57335 44201
rect 54853 43353 54909 43355
rect 54853 43301 54855 43353
rect 54855 43301 54907 43353
rect 54907 43301 54909 43353
rect 54853 43299 54909 43301
rect 55064 43353 55120 43355
rect 55064 43301 55066 43353
rect 55066 43301 55118 43353
rect 55118 43301 55120 43353
rect 55064 43299 55120 43301
rect 55276 43353 55332 43355
rect 55276 43301 55278 43353
rect 55278 43301 55330 43353
rect 55330 43301 55332 43353
rect 55276 43299 55332 43301
rect 55487 43353 55543 43355
rect 55487 43301 55489 43353
rect 55489 43301 55541 43353
rect 55541 43301 55543 43353
rect 55487 43299 55543 43301
rect 56013 42453 56069 42455
rect 56013 42401 56015 42453
rect 56015 42401 56067 42453
rect 56067 42401 56069 42453
rect 56013 42399 56069 42401
rect 56224 42453 56280 42455
rect 56224 42401 56226 42453
rect 56226 42401 56278 42453
rect 56278 42401 56280 42453
rect 56224 42399 56280 42401
rect 56435 42453 56491 42455
rect 56435 42401 56437 42453
rect 56437 42401 56489 42453
rect 56489 42401 56491 42453
rect 56435 42399 56491 42401
rect 56646 42453 56702 42455
rect 56646 42401 56648 42453
rect 56648 42401 56700 42453
rect 56700 42401 56702 42453
rect 56646 42399 56702 42401
rect 56857 42453 56913 42455
rect 56857 42401 56859 42453
rect 56859 42401 56911 42453
rect 56911 42401 56913 42453
rect 56857 42399 56913 42401
rect 57068 42453 57124 42455
rect 57068 42401 57070 42453
rect 57070 42401 57122 42453
rect 57122 42401 57124 42453
rect 57068 42399 57124 42401
rect 57279 42453 57335 42455
rect 57279 42401 57281 42453
rect 57281 42401 57333 42453
rect 57333 42401 57335 42453
rect 57279 42399 57335 42401
rect 54853 41553 54909 41555
rect 54853 41501 54855 41553
rect 54855 41501 54907 41553
rect 54907 41501 54909 41553
rect 54853 41499 54909 41501
rect 55064 41553 55120 41555
rect 55064 41501 55066 41553
rect 55066 41501 55118 41553
rect 55118 41501 55120 41553
rect 55064 41499 55120 41501
rect 55276 41553 55332 41555
rect 55276 41501 55278 41553
rect 55278 41501 55330 41553
rect 55330 41501 55332 41553
rect 55276 41499 55332 41501
rect 55487 41553 55543 41555
rect 55487 41501 55489 41553
rect 55489 41501 55541 41553
rect 55541 41501 55543 41553
rect 55487 41499 55543 41501
rect 56013 40653 56069 40655
rect 56013 40601 56015 40653
rect 56015 40601 56067 40653
rect 56067 40601 56069 40653
rect 56013 40599 56069 40601
rect 56224 40653 56280 40655
rect 56224 40601 56226 40653
rect 56226 40601 56278 40653
rect 56278 40601 56280 40653
rect 56224 40599 56280 40601
rect 56435 40653 56491 40655
rect 56435 40601 56437 40653
rect 56437 40601 56489 40653
rect 56489 40601 56491 40653
rect 56435 40599 56491 40601
rect 56646 40653 56702 40655
rect 56646 40601 56648 40653
rect 56648 40601 56700 40653
rect 56700 40601 56702 40653
rect 56646 40599 56702 40601
rect 56857 40653 56913 40655
rect 56857 40601 56859 40653
rect 56859 40601 56911 40653
rect 56911 40601 56913 40653
rect 56857 40599 56913 40601
rect 57068 40653 57124 40655
rect 57068 40601 57070 40653
rect 57070 40601 57122 40653
rect 57122 40601 57124 40653
rect 57068 40599 57124 40601
rect 57279 40653 57335 40655
rect 57279 40601 57281 40653
rect 57281 40601 57333 40653
rect 57333 40601 57335 40653
rect 57279 40599 57335 40601
rect 54853 39753 54909 39755
rect 54853 39701 54855 39753
rect 54855 39701 54907 39753
rect 54907 39701 54909 39753
rect 54853 39699 54909 39701
rect 55064 39753 55120 39755
rect 55064 39701 55066 39753
rect 55066 39701 55118 39753
rect 55118 39701 55120 39753
rect 55064 39699 55120 39701
rect 55276 39753 55332 39755
rect 55276 39701 55278 39753
rect 55278 39701 55330 39753
rect 55330 39701 55332 39753
rect 55276 39699 55332 39701
rect 55487 39753 55543 39755
rect 55487 39701 55489 39753
rect 55489 39701 55541 39753
rect 55541 39701 55543 39753
rect 55487 39699 55543 39701
rect 56013 38853 56069 38855
rect 56013 38801 56015 38853
rect 56015 38801 56067 38853
rect 56067 38801 56069 38853
rect 56013 38799 56069 38801
rect 56224 38853 56280 38855
rect 56224 38801 56226 38853
rect 56226 38801 56278 38853
rect 56278 38801 56280 38853
rect 56224 38799 56280 38801
rect 56435 38853 56491 38855
rect 56435 38801 56437 38853
rect 56437 38801 56489 38853
rect 56489 38801 56491 38853
rect 56435 38799 56491 38801
rect 56646 38853 56702 38855
rect 56646 38801 56648 38853
rect 56648 38801 56700 38853
rect 56700 38801 56702 38853
rect 56646 38799 56702 38801
rect 56857 38853 56913 38855
rect 56857 38801 56859 38853
rect 56859 38801 56911 38853
rect 56911 38801 56913 38853
rect 56857 38799 56913 38801
rect 57068 38853 57124 38855
rect 57068 38801 57070 38853
rect 57070 38801 57122 38853
rect 57122 38801 57124 38853
rect 57068 38799 57124 38801
rect 57279 38853 57335 38855
rect 57279 38801 57281 38853
rect 57281 38801 57333 38853
rect 57333 38801 57335 38853
rect 57279 38799 57335 38801
rect 54853 37953 54909 37955
rect 54853 37901 54855 37953
rect 54855 37901 54907 37953
rect 54907 37901 54909 37953
rect 54853 37899 54909 37901
rect 55064 37953 55120 37955
rect 55064 37901 55066 37953
rect 55066 37901 55118 37953
rect 55118 37901 55120 37953
rect 55064 37899 55120 37901
rect 55276 37953 55332 37955
rect 55276 37901 55278 37953
rect 55278 37901 55330 37953
rect 55330 37901 55332 37953
rect 55276 37899 55332 37901
rect 55487 37953 55543 37955
rect 55487 37901 55489 37953
rect 55489 37901 55541 37953
rect 55541 37901 55543 37953
rect 55487 37899 55543 37901
rect 56013 37053 56069 37055
rect 56013 37001 56015 37053
rect 56015 37001 56067 37053
rect 56067 37001 56069 37053
rect 56013 36999 56069 37001
rect 56224 37053 56280 37055
rect 56224 37001 56226 37053
rect 56226 37001 56278 37053
rect 56278 37001 56280 37053
rect 56224 36999 56280 37001
rect 56435 37053 56491 37055
rect 56435 37001 56437 37053
rect 56437 37001 56489 37053
rect 56489 37001 56491 37053
rect 56435 36999 56491 37001
rect 56646 37053 56702 37055
rect 56646 37001 56648 37053
rect 56648 37001 56700 37053
rect 56700 37001 56702 37053
rect 56646 36999 56702 37001
rect 56857 37053 56913 37055
rect 56857 37001 56859 37053
rect 56859 37001 56911 37053
rect 56911 37001 56913 37053
rect 56857 36999 56913 37001
rect 57068 37053 57124 37055
rect 57068 37001 57070 37053
rect 57070 37001 57122 37053
rect 57122 37001 57124 37053
rect 57068 36999 57124 37001
rect 57279 37053 57335 37055
rect 57279 37001 57281 37053
rect 57281 37001 57333 37053
rect 57333 37001 57335 37053
rect 57279 36999 57335 37001
rect 54853 36153 54909 36155
rect 54853 36101 54855 36153
rect 54855 36101 54907 36153
rect 54907 36101 54909 36153
rect 54853 36099 54909 36101
rect 55064 36153 55120 36155
rect 55064 36101 55066 36153
rect 55066 36101 55118 36153
rect 55118 36101 55120 36153
rect 55064 36099 55120 36101
rect 55276 36153 55332 36155
rect 55276 36101 55278 36153
rect 55278 36101 55330 36153
rect 55330 36101 55332 36153
rect 55276 36099 55332 36101
rect 55487 36153 55543 36155
rect 55487 36101 55489 36153
rect 55489 36101 55541 36153
rect 55541 36101 55543 36153
rect 55487 36099 55543 36101
rect 57996 33955 58052 34011
rect 58208 33955 58264 34011
rect 57996 33737 58052 33793
rect 58208 33737 58264 33793
rect 57996 33520 58052 33576
rect 58208 33520 58264 33576
rect 27474 33085 27530 33141
rect 27686 33085 27742 33141
rect 27474 32867 27530 32923
rect 27686 32867 27742 32923
rect 27474 32649 27530 32705
rect 27686 32649 27742 32705
rect 27474 32431 27530 32487
rect 27686 32431 27742 32487
rect 27474 31204 27476 31252
rect 27476 31204 27528 31252
rect 27528 31204 27530 31252
rect 27474 31196 27530 31204
rect 27686 31204 27688 31252
rect 27688 31204 27740 31252
rect 27740 31204 27742 31252
rect 27686 31196 27742 31204
rect 27474 30986 27476 31034
rect 27476 30986 27528 31034
rect 27528 30986 27530 31034
rect 27474 30978 27530 30986
rect 27686 30986 27688 31034
rect 27688 30986 27740 31034
rect 27740 30986 27742 31034
rect 27686 30978 27742 30986
rect 27474 30769 27476 30816
rect 27476 30769 27528 30816
rect 27528 30769 27530 30816
rect 27474 30760 27530 30769
rect 27686 30769 27688 30816
rect 27688 30769 27740 30816
rect 27740 30769 27742 30816
rect 27686 30760 27742 30769
rect 27474 30551 27476 30598
rect 27476 30551 27528 30598
rect 27528 30551 27530 30598
rect 27474 30542 27530 30551
rect 27686 30551 27688 30598
rect 27688 30551 27740 30598
rect 27740 30551 27742 30598
rect 27686 30542 27742 30551
rect 25404 27267 25460 27323
rect 25528 27267 25584 27323
rect 25652 27267 25708 27323
rect 25776 27267 25832 27323
rect 25900 27267 25956 27323
rect 25404 27143 25460 27199
rect 25528 27143 25584 27199
rect 25652 27143 25708 27199
rect 25776 27143 25832 27199
rect 25900 27143 25956 27199
rect 25404 27019 25460 27075
rect 25528 27019 25584 27075
rect 25652 27019 25708 27075
rect 25776 27019 25832 27075
rect 25900 27019 25956 27075
rect 25404 26895 25460 26951
rect 25528 26895 25584 26951
rect 25652 26895 25708 26951
rect 25776 26895 25832 26951
rect 25900 26895 25956 26951
rect 25404 26771 25460 26827
rect 25528 26771 25584 26827
rect 25652 26771 25708 26827
rect 25776 26771 25832 26827
rect 25900 26771 25956 26827
rect 25404 26647 25460 26703
rect 25528 26647 25584 26703
rect 25652 26647 25708 26703
rect 25776 26647 25832 26703
rect 25900 26647 25956 26703
rect 25404 26523 25460 26579
rect 25528 26523 25584 26579
rect 25652 26523 25708 26579
rect 25776 26523 25832 26579
rect 25900 26523 25956 26579
rect 26450 26126 26610 26286
rect 26092 25807 26252 25967
rect 25756 25487 25916 25647
rect 25421 25168 25581 25328
rect 25081 24477 25241 24637
rect 24744 24156 24904 24316
rect 24416 23835 24576 23995
rect 24057 23513 24217 23673
rect 26465 19532 26625 19692
rect 26858 24074 27122 24075
rect 26858 24022 26861 24074
rect 26861 24022 26913 24074
rect 26913 24022 27073 24074
rect 27073 24022 27122 24074
rect 26858 23857 27122 24022
rect 26858 23805 26861 23857
rect 26861 23805 26913 23857
rect 26913 23805 27073 23857
rect 27073 23805 27122 23857
rect 26858 23639 27122 23805
rect 26858 23587 26861 23639
rect 26861 23587 26913 23639
rect 26913 23587 27073 23639
rect 27073 23587 27122 23639
rect 26858 23421 27122 23587
rect 26858 23369 26861 23421
rect 26861 23369 26913 23421
rect 26913 23369 27073 23421
rect 27073 23369 27122 23421
rect 26858 23204 27122 23369
rect 26858 23187 26861 23204
rect 26861 23187 26913 23204
rect 26913 23187 27073 23204
rect 27073 23187 27122 23204
rect 26924 20540 27073 20570
rect 27073 20540 27084 20570
rect 26924 20410 27084 20540
rect 26924 20157 27084 20226
rect 26924 20105 27073 20157
rect 27073 20105 27084 20157
rect 26924 20066 27084 20105
rect 26107 19187 26267 19347
rect 25771 18867 25931 19027
rect 25434 18524 25594 18684
rect 25094 18190 25254 18350
rect 24757 17817 24917 17977
rect 24429 17496 24589 17656
rect 24069 17157 24229 17317
rect 26859 14063 26915 14119
rect 27071 14063 27127 14119
rect 26859 13846 26915 13902
rect 27071 13846 27127 13902
rect 26859 13628 26915 13684
rect 27071 13628 27127 13684
rect 26859 13411 26915 13467
rect 27071 13411 27127 13467
rect 26859 13193 26915 13249
rect 27071 13193 27127 13249
rect 26859 12975 26915 13031
rect 27071 12975 27127 13031
rect 26859 12757 26915 12813
rect 27071 12757 27127 12813
rect 26859 12540 26915 12596
rect 27071 12540 27127 12596
rect 26859 12322 26915 12378
rect 27071 12322 27127 12378
rect 26859 12105 26915 12161
rect 27071 12105 27127 12161
rect 26859 9351 26915 9407
rect 27071 9351 27127 9407
rect 26859 9134 26915 9190
rect 27071 9134 27127 9190
rect 26859 8916 26915 8972
rect 27071 8916 27127 8972
rect 26859 8698 26915 8754
rect 27071 8698 27127 8754
rect 26859 8480 26915 8536
rect 27071 8480 27127 8536
rect 26859 8263 26915 8319
rect 27071 8263 27127 8319
rect 26859 5523 26861 5539
rect 26861 5523 26913 5539
rect 26913 5523 26915 5539
rect 26859 5483 26915 5523
rect 27071 5523 27073 5539
rect 27073 5523 27125 5539
rect 27125 5523 27127 5539
rect 27071 5483 27127 5523
rect 26859 5306 26861 5321
rect 26861 5306 26913 5321
rect 26913 5306 26915 5321
rect 26859 5265 26915 5306
rect 27071 5306 27073 5321
rect 27073 5306 27125 5321
rect 27125 5306 27127 5321
rect 27071 5265 27127 5306
rect 27474 26743 27530 26799
rect 27686 26743 27742 26799
rect 27474 26525 27530 26581
rect 27686 26525 27742 26581
rect 27474 24972 27530 25028
rect 27686 24972 27742 25028
rect 27474 24754 27530 24810
rect 27686 24754 27742 24810
rect 27475 22934 27476 22936
rect 27476 22934 27528 22936
rect 27528 22934 27688 22936
rect 27688 22934 27739 22936
rect 27475 22768 27739 22934
rect 27475 22716 27476 22768
rect 27476 22716 27528 22768
rect 27528 22716 27688 22768
rect 27688 22716 27739 22768
rect 27475 22551 27739 22716
rect 27475 22499 27476 22551
rect 27476 22499 27528 22551
rect 27528 22499 27688 22551
rect 27688 22499 27739 22551
rect 27475 22333 27739 22499
rect 27475 22281 27476 22333
rect 27476 22281 27528 22333
rect 27528 22281 27688 22333
rect 27688 22281 27739 22333
rect 27475 22115 27739 22281
rect 27475 22063 27476 22115
rect 27476 22063 27528 22115
rect 27528 22063 27688 22115
rect 27688 22063 27739 22115
rect 27475 22048 27739 22063
rect 27474 16457 27530 16470
rect 27474 16414 27476 16457
rect 27476 16414 27528 16457
rect 27528 16414 27530 16457
rect 27686 16457 27742 16470
rect 27686 16414 27688 16457
rect 27688 16414 27740 16457
rect 27740 16414 27742 16457
rect 27474 16239 27530 16253
rect 27474 16197 27476 16239
rect 27476 16197 27528 16239
rect 27528 16197 27530 16239
rect 27686 16239 27742 16253
rect 27686 16197 27688 16239
rect 27688 16197 27740 16239
rect 27740 16197 27742 16239
rect 27474 16022 27530 16035
rect 27474 15979 27476 16022
rect 27476 15979 27528 16022
rect 27528 15979 27530 16022
rect 27686 16022 27742 16035
rect 27686 15979 27688 16022
rect 27688 15979 27740 16022
rect 27740 15979 27742 16022
rect 27474 15804 27530 15818
rect 27474 15762 27476 15804
rect 27476 15762 27528 15804
rect 27528 15762 27530 15804
rect 27686 15804 27742 15818
rect 27686 15762 27688 15804
rect 27688 15762 27740 15804
rect 27740 15762 27742 15804
rect 27474 15586 27530 15600
rect 27474 15544 27476 15586
rect 27476 15544 27528 15586
rect 27528 15544 27530 15586
rect 27686 15586 27742 15600
rect 27686 15544 27688 15586
rect 27688 15544 27740 15586
rect 27740 15544 27742 15586
rect 27474 15369 27530 15382
rect 27474 15326 27476 15369
rect 27476 15326 27528 15369
rect 27528 15326 27530 15369
rect 27686 15369 27742 15382
rect 27686 15326 27688 15369
rect 27688 15326 27740 15369
rect 27740 15326 27742 15369
rect 27474 15151 27530 15164
rect 27474 15108 27476 15151
rect 27476 15108 27528 15151
rect 27528 15108 27530 15151
rect 27686 15151 27742 15164
rect 27686 15108 27688 15151
rect 27688 15108 27740 15151
rect 27740 15108 27742 15151
rect 27474 14933 27530 14947
rect 27474 14891 27476 14933
rect 27476 14891 27528 14933
rect 27528 14891 27530 14933
rect 27686 14933 27742 14947
rect 27686 14891 27688 14933
rect 27688 14891 27740 14933
rect 27740 14891 27742 14933
rect 27474 14716 27530 14729
rect 27474 14673 27476 14716
rect 27476 14673 27528 14716
rect 27528 14673 27530 14716
rect 27686 14716 27742 14729
rect 27686 14673 27688 14716
rect 27688 14673 27740 14716
rect 27740 14673 27742 14716
rect 27474 14498 27530 14512
rect 27474 14456 27476 14498
rect 27476 14456 27528 14498
rect 27528 14456 27530 14498
rect 27686 14498 27742 14512
rect 27686 14456 27688 14498
rect 27688 14456 27740 14498
rect 27740 14456 27742 14498
rect 27474 14229 27476 14231
rect 27476 14229 27528 14231
rect 27528 14229 27530 14231
rect 27474 14175 27530 14229
rect 27686 14229 27688 14231
rect 27688 14229 27740 14231
rect 27740 14229 27742 14231
rect 27686 14175 27742 14229
rect 27474 14011 27476 14014
rect 27476 14011 27528 14014
rect 27528 14011 27530 14014
rect 27474 13958 27530 14011
rect 27686 14011 27688 14014
rect 27688 14011 27740 14014
rect 27740 14011 27742 14014
rect 27686 13958 27742 14011
rect 27474 13793 27476 13796
rect 27476 13793 27528 13796
rect 27528 13793 27530 13796
rect 27474 13740 27530 13793
rect 27686 13793 27688 13796
rect 27688 13793 27740 13796
rect 27740 13793 27742 13796
rect 27686 13740 27742 13793
rect 27474 13576 27476 13578
rect 27476 13576 27528 13578
rect 27528 13576 27530 13578
rect 27474 13522 27530 13576
rect 27686 13576 27688 13578
rect 27688 13576 27740 13578
rect 27740 13576 27742 13578
rect 27686 13522 27742 13576
rect 27474 13358 27476 13361
rect 27476 13358 27528 13361
rect 27528 13358 27530 13361
rect 27474 13305 27530 13358
rect 27686 13358 27688 13361
rect 27688 13358 27740 13361
rect 27740 13358 27742 13361
rect 27686 13305 27742 13358
rect 27474 11399 27476 11406
rect 27476 11399 27528 11406
rect 27528 11399 27530 11406
rect 27474 11350 27530 11399
rect 27686 11399 27688 11406
rect 27688 11399 27740 11406
rect 27740 11399 27742 11406
rect 27686 11350 27742 11399
rect 27474 11182 27476 11189
rect 27476 11182 27528 11189
rect 27528 11182 27530 11189
rect 27474 11133 27530 11182
rect 27686 11182 27688 11189
rect 27688 11182 27740 11189
rect 27740 11182 27742 11189
rect 27686 11133 27742 11182
rect 27474 10964 27476 10971
rect 27476 10964 27528 10971
rect 27528 10964 27530 10971
rect 27474 10915 27530 10964
rect 27686 10964 27688 10971
rect 27688 10964 27740 10971
rect 27740 10964 27742 10971
rect 27686 10915 27742 10964
rect 27474 10746 27476 10753
rect 27476 10746 27528 10753
rect 27528 10746 27530 10753
rect 27474 10697 27530 10746
rect 27686 10746 27688 10753
rect 27688 10746 27740 10753
rect 27740 10746 27742 10753
rect 27686 10697 27742 10746
rect 27474 10529 27476 10535
rect 27476 10529 27528 10535
rect 27528 10529 27530 10535
rect 27474 10479 27530 10529
rect 27686 10529 27688 10535
rect 27688 10529 27740 10535
rect 27740 10529 27742 10535
rect 27686 10479 27742 10529
rect 27474 10311 27476 10318
rect 27476 10311 27528 10318
rect 27528 10311 27530 10318
rect 27474 10262 27530 10311
rect 27686 10311 27688 10318
rect 27688 10311 27740 10318
rect 27740 10311 27742 10318
rect 27686 10262 27742 10311
rect 57381 33085 57437 33141
rect 57593 33085 57649 33141
rect 57381 32867 57437 32923
rect 57593 32867 57649 32923
rect 57381 32649 57437 32705
rect 57593 32649 57649 32705
rect 57381 32431 57437 32487
rect 57593 32431 57649 32487
rect 57381 31204 57383 31252
rect 57383 31204 57435 31252
rect 57435 31204 57437 31252
rect 57381 31196 57437 31204
rect 57593 31204 57595 31252
rect 57595 31204 57647 31252
rect 57647 31204 57649 31252
rect 57593 31196 57649 31204
rect 57381 30986 57383 31034
rect 57383 30986 57435 31034
rect 57435 30986 57437 31034
rect 57381 30978 57437 30986
rect 57593 30986 57595 31034
rect 57595 30986 57647 31034
rect 57647 30986 57649 31034
rect 57593 30978 57649 30986
rect 57381 30769 57383 30816
rect 57383 30769 57435 30816
rect 57435 30769 57437 30816
rect 57381 30760 57437 30769
rect 57593 30769 57595 30816
rect 57595 30769 57647 30816
rect 57647 30769 57649 30816
rect 57593 30760 57649 30769
rect 57381 30551 57383 30598
rect 57383 30551 57435 30598
rect 57435 30551 57437 30598
rect 57381 30542 57437 30551
rect 57593 30551 57595 30598
rect 57595 30551 57647 30598
rect 57647 30551 57649 30598
rect 57593 30542 57649 30551
rect 57381 26743 57437 26799
rect 57593 26743 57649 26799
rect 57381 26525 57437 26581
rect 57593 26525 57649 26581
rect 57363 22768 57627 22923
rect 57363 22716 57383 22768
rect 57383 22716 57435 22768
rect 57435 22716 57595 22768
rect 57595 22716 57627 22768
rect 57363 22551 57627 22716
rect 57363 22499 57383 22551
rect 57383 22499 57435 22551
rect 57435 22499 57595 22551
rect 57595 22499 57627 22551
rect 57363 22333 57627 22499
rect 57363 22281 57383 22333
rect 57383 22281 57435 22333
rect 57435 22281 57595 22333
rect 57595 22281 57627 22333
rect 57363 22115 57627 22281
rect 57363 22063 57383 22115
rect 57383 22063 57435 22115
rect 57435 22063 57595 22115
rect 57595 22063 57627 22115
rect 57363 22035 57627 22063
rect 57381 16675 57437 16678
rect 57381 16623 57383 16675
rect 57383 16623 57435 16675
rect 57435 16623 57437 16675
rect 57381 16622 57437 16623
rect 57593 16675 57649 16678
rect 57593 16623 57595 16675
rect 57595 16623 57647 16675
rect 57647 16623 57649 16675
rect 57593 16622 57649 16623
rect 57381 16457 57437 16461
rect 57381 16405 57383 16457
rect 57383 16405 57435 16457
rect 57435 16405 57437 16457
rect 57593 16457 57649 16461
rect 57593 16405 57595 16457
rect 57595 16405 57647 16457
rect 57647 16405 57649 16457
rect 57381 16239 57437 16243
rect 57381 16187 57383 16239
rect 57383 16187 57435 16239
rect 57435 16187 57437 16239
rect 57593 16239 57649 16243
rect 57593 16187 57595 16239
rect 57595 16187 57647 16239
rect 57647 16187 57649 16239
rect 57381 16022 57437 16026
rect 57381 15970 57383 16022
rect 57383 15970 57435 16022
rect 57435 15970 57437 16022
rect 57593 16022 57649 16026
rect 57593 15970 57595 16022
rect 57595 15970 57647 16022
rect 57647 15970 57649 16022
rect 57381 15804 57437 15808
rect 57381 15752 57383 15804
rect 57383 15752 57435 15804
rect 57435 15752 57437 15804
rect 57593 15804 57649 15808
rect 57593 15752 57595 15804
rect 57595 15752 57647 15804
rect 57647 15752 57649 15804
rect 57381 15586 57437 15590
rect 57381 15534 57383 15586
rect 57383 15534 57435 15586
rect 57435 15534 57437 15586
rect 57593 15586 57649 15590
rect 57593 15534 57595 15586
rect 57595 15534 57647 15586
rect 57647 15534 57649 15586
rect 57381 15369 57437 15372
rect 57381 15317 57383 15369
rect 57383 15317 57435 15369
rect 57435 15317 57437 15369
rect 57381 15316 57437 15317
rect 57593 15369 57649 15372
rect 57593 15317 57595 15369
rect 57595 15317 57647 15369
rect 57647 15317 57649 15369
rect 57593 15316 57649 15317
rect 57381 15151 57437 15155
rect 57381 15099 57383 15151
rect 57383 15099 57435 15151
rect 57435 15099 57437 15151
rect 57593 15151 57649 15155
rect 57593 15099 57595 15151
rect 57595 15099 57647 15151
rect 57647 15099 57649 15151
rect 57381 14933 57437 14937
rect 57381 14881 57383 14933
rect 57383 14881 57435 14933
rect 57435 14881 57437 14933
rect 57593 14933 57649 14937
rect 57593 14881 57595 14933
rect 57595 14881 57647 14933
rect 57647 14881 57649 14933
rect 57381 14716 57437 14720
rect 57381 14664 57383 14716
rect 57383 14664 57435 14716
rect 57435 14664 57437 14716
rect 57593 14716 57649 14720
rect 57593 14664 57595 14716
rect 57595 14664 57647 14716
rect 57647 14664 57649 14716
rect 57381 11399 57383 11406
rect 57383 11399 57435 11406
rect 57435 11399 57437 11406
rect 57381 11350 57437 11399
rect 57593 11399 57595 11406
rect 57595 11399 57647 11406
rect 57647 11399 57649 11406
rect 57593 11350 57649 11399
rect 57381 11182 57383 11189
rect 57383 11182 57435 11189
rect 57435 11182 57437 11189
rect 57381 11133 57437 11182
rect 57593 11182 57595 11189
rect 57595 11182 57647 11189
rect 57647 11182 57649 11189
rect 57593 11133 57649 11182
rect 57381 10964 57383 10971
rect 57383 10964 57435 10971
rect 57435 10964 57437 10971
rect 57381 10915 57437 10964
rect 57593 10964 57595 10971
rect 57595 10964 57647 10971
rect 57647 10964 57649 10971
rect 57593 10915 57649 10964
rect 57381 10746 57383 10753
rect 57383 10746 57435 10753
rect 57435 10746 57437 10753
rect 57381 10697 57437 10746
rect 57593 10746 57595 10753
rect 57595 10746 57647 10753
rect 57647 10746 57649 10753
rect 57593 10697 57649 10746
rect 57381 10529 57383 10535
rect 57383 10529 57435 10535
rect 57435 10529 57437 10535
rect 57381 10479 57437 10529
rect 57593 10529 57595 10535
rect 57595 10529 57647 10535
rect 57647 10529 57649 10535
rect 57593 10479 57649 10529
rect 57381 10311 57383 10318
rect 57383 10311 57435 10318
rect 57435 10311 57437 10318
rect 57381 10262 57437 10311
rect 57593 10311 57595 10318
rect 57595 10311 57647 10318
rect 57647 10311 57649 10318
rect 57593 10262 57649 10311
rect 51766 9811 51822 9971
rect 49906 8897 50066 8953
rect 27474 7534 27530 7535
rect 27474 7482 27476 7534
rect 27476 7482 27528 7534
rect 27528 7482 27530 7534
rect 27474 7479 27530 7482
rect 27686 7534 27742 7535
rect 27686 7482 27688 7534
rect 27688 7482 27740 7534
rect 27740 7482 27742 7534
rect 27686 7479 27742 7482
rect 27474 7316 27530 7317
rect 27474 7264 27476 7316
rect 27476 7264 27528 7316
rect 27528 7264 27530 7316
rect 27474 7261 27530 7264
rect 27686 7316 27742 7317
rect 27686 7264 27688 7316
rect 27688 7264 27740 7316
rect 27740 7264 27742 7316
rect 27686 7261 27742 7264
rect 27474 7047 27476 7099
rect 27476 7047 27528 7099
rect 27528 7047 27530 7099
rect 27474 7043 27530 7047
rect 27686 7047 27688 7099
rect 27688 7047 27740 7099
rect 27740 7047 27742 7099
rect 27686 7043 27742 7047
rect 28273 6780 28329 6836
rect 28484 6780 28540 6836
rect 28696 6780 28752 6836
rect 28907 6780 28963 6836
rect 28273 6562 28329 6618
rect 28484 6562 28540 6618
rect 28696 6562 28752 6618
rect 28907 6562 28963 6618
rect 28273 6344 28329 6400
rect 28484 6344 28540 6400
rect 28696 6344 28752 6400
rect 28907 6344 28963 6400
rect 27474 6064 27530 6120
rect 27686 6064 27742 6120
rect 27474 5846 27530 5902
rect 27686 5846 27742 5902
rect 26859 4472 26915 4528
rect 27071 4472 27127 4528
rect 26859 4254 26915 4310
rect 27071 4254 27127 4310
rect 27474 3781 27530 3837
rect 27686 3781 27742 3837
rect 27474 3563 27530 3619
rect 27686 3563 27742 3619
rect 28801 3781 28857 3837
rect 28801 3563 28857 3619
rect 43800 2988 43960 3044
rect 57381 8840 57437 8854
rect 57381 8798 57383 8840
rect 57383 8798 57435 8840
rect 57435 8798 57437 8840
rect 57593 8840 57649 8854
rect 57593 8798 57595 8840
rect 57595 8798 57647 8840
rect 57647 8798 57649 8840
rect 57381 8622 57437 8636
rect 57381 8580 57383 8622
rect 57383 8580 57435 8622
rect 57435 8580 57437 8622
rect 57593 8622 57649 8636
rect 57593 8580 57595 8622
rect 57595 8580 57647 8622
rect 57647 8580 57649 8622
rect 57381 8404 57437 8419
rect 57381 8363 57383 8404
rect 57383 8363 57435 8404
rect 57435 8363 57437 8404
rect 57593 8404 57649 8419
rect 57593 8363 57595 8404
rect 57595 8363 57647 8404
rect 57647 8363 57649 8404
rect 57381 8187 57437 8201
rect 57381 8145 57383 8187
rect 57383 8145 57435 8187
rect 57435 8145 57437 8187
rect 57593 8187 57649 8201
rect 57593 8145 57595 8187
rect 57595 8145 57647 8187
rect 57647 8145 57649 8187
rect 57381 7969 57437 7983
rect 57381 7927 57383 7969
rect 57383 7927 57435 7969
rect 57435 7927 57437 7969
rect 57593 7969 57649 7983
rect 57593 7927 57595 7969
rect 57595 7927 57647 7969
rect 57647 7927 57649 7969
rect 57381 7752 57437 7766
rect 57381 7710 57383 7752
rect 57383 7710 57435 7752
rect 57435 7710 57437 7752
rect 57593 7752 57649 7766
rect 57593 7710 57595 7752
rect 57595 7710 57647 7752
rect 57647 7710 57649 7752
rect 57381 7534 57437 7548
rect 57381 7492 57383 7534
rect 57383 7492 57435 7534
rect 57435 7492 57437 7534
rect 57593 7534 57649 7548
rect 57593 7492 57595 7534
rect 57595 7492 57647 7534
rect 57647 7492 57649 7534
rect 57381 7316 57437 7330
rect 57381 7274 57383 7316
rect 57383 7274 57435 7316
rect 57435 7274 57437 7316
rect 57593 7316 57649 7330
rect 57593 7274 57595 7316
rect 57595 7274 57647 7316
rect 57647 7274 57649 7316
rect 57381 7099 57437 7113
rect 57381 7057 57383 7099
rect 57383 7057 57435 7099
rect 57435 7057 57437 7099
rect 57593 7099 57649 7113
rect 57593 7057 57595 7099
rect 57595 7057 57647 7099
rect 57647 7057 57649 7099
rect 56160 6780 56216 6836
rect 56371 6780 56427 6836
rect 56583 6780 56639 6836
rect 56794 6780 56850 6836
rect 56160 6562 56216 6618
rect 56371 6562 56427 6618
rect 56583 6562 56639 6618
rect 56794 6562 56850 6618
rect 56160 6344 56216 6400
rect 56371 6344 56427 6400
rect 56583 6344 56639 6400
rect 56794 6344 56850 6400
rect 57381 6064 57437 6120
rect 57593 6064 57649 6120
rect 57381 5846 57437 5902
rect 57593 5846 57649 5902
rect 57381 3781 57437 3837
rect 57593 3781 57649 3837
rect 57381 3563 57437 3619
rect 57593 3563 57649 3619
rect 57996 33302 58052 33358
rect 58208 33302 58264 33358
rect 57996 33084 58052 33140
rect 58208 33084 58264 33140
rect 57996 32866 58052 32922
rect 58208 32866 58264 32922
rect 57996 32649 58052 32705
rect 58208 32649 58264 32705
rect 57996 32431 58052 32487
rect 58208 32431 58264 32487
rect 57996 32075 57998 32088
rect 57998 32075 58050 32088
rect 58050 32075 58052 32088
rect 57996 32032 58052 32075
rect 58208 32075 58210 32088
rect 58210 32075 58262 32088
rect 58262 32075 58264 32088
rect 58208 32032 58264 32075
rect 57996 31857 57998 31870
rect 57998 31857 58050 31870
rect 58050 31857 58052 31870
rect 57996 31814 58052 31857
rect 58208 31857 58210 31870
rect 58210 31857 58262 31870
rect 58262 31857 58264 31870
rect 58208 31814 58264 31857
rect 57996 31639 57998 31652
rect 57998 31639 58050 31652
rect 58050 31639 58052 31652
rect 57996 31596 58052 31639
rect 58208 31639 58210 31652
rect 58210 31639 58262 31652
rect 58262 31639 58264 31652
rect 58208 31596 58264 31639
rect 57996 29950 58052 29968
rect 57996 29912 57998 29950
rect 57998 29912 58050 29950
rect 58050 29912 58052 29950
rect 58208 29950 58264 29968
rect 58208 29912 58210 29950
rect 58210 29912 58262 29950
rect 58262 29912 58264 29950
rect 57996 29733 58052 29750
rect 57996 29694 57998 29733
rect 57998 29694 58050 29733
rect 58050 29694 58052 29733
rect 58208 29733 58264 29750
rect 58208 29694 58210 29733
rect 58210 29694 58262 29733
rect 58262 29694 58264 29733
rect 57996 29515 58052 29533
rect 57996 29477 57998 29515
rect 57998 29477 58050 29515
rect 58050 29477 58052 29515
rect 58208 29515 58264 29533
rect 58208 29477 58210 29515
rect 58210 29477 58262 29515
rect 58262 29477 58264 29515
rect 57996 29297 58052 29315
rect 57996 29259 57998 29297
rect 57998 29259 58050 29297
rect 58050 29259 58052 29297
rect 58208 29297 58264 29315
rect 58208 29259 58210 29297
rect 58210 29259 58262 29297
rect 58262 29259 58264 29297
rect 57996 29080 58052 29098
rect 57996 29042 57998 29080
rect 57998 29042 58050 29080
rect 58050 29042 58052 29080
rect 58208 29080 58264 29098
rect 58208 29042 58210 29080
rect 58210 29042 58262 29080
rect 58262 29042 58264 29080
rect 57996 28862 58052 28880
rect 57996 28824 57998 28862
rect 57998 28824 58050 28862
rect 58050 28824 58052 28862
rect 58208 28862 58264 28880
rect 58208 28824 58210 28862
rect 58210 28824 58262 28862
rect 58262 28824 58264 28862
rect 57996 28644 58052 28662
rect 57996 28606 57998 28644
rect 57998 28606 58050 28644
rect 58050 28606 58052 28644
rect 58208 28644 58264 28662
rect 58208 28606 58210 28644
rect 58210 28606 58262 28644
rect 58262 28606 58264 28644
rect 57996 28427 58052 28444
rect 57996 28388 57998 28427
rect 57998 28388 58050 28427
rect 58050 28388 58052 28427
rect 58208 28427 58264 28444
rect 58208 28388 58210 28427
rect 58210 28388 58262 28427
rect 58262 28388 58264 28427
rect 57996 28209 58052 28227
rect 57996 28171 57998 28209
rect 57998 28171 58050 28209
rect 58050 28171 58052 28209
rect 58208 28209 58264 28227
rect 58208 28171 58210 28209
rect 58210 28171 58262 28209
rect 58262 28171 58264 28209
rect 57996 27992 58052 28009
rect 57996 27953 57998 27992
rect 57998 27953 58050 27992
rect 58050 27953 58052 27992
rect 58208 27992 58264 28009
rect 58208 27953 58210 27992
rect 58210 27953 58262 27992
rect 58262 27953 58264 27992
rect 57996 27774 58052 27792
rect 57996 27736 57998 27774
rect 57998 27736 58050 27774
rect 58050 27736 58052 27774
rect 58208 27774 58264 27792
rect 58208 27736 58210 27774
rect 58210 27736 58262 27774
rect 58262 27736 58264 27774
rect 57996 27556 58052 27574
rect 57996 27518 57998 27556
rect 57998 27518 58050 27556
rect 58050 27518 58052 27556
rect 58208 27556 58264 27574
rect 58208 27518 58210 27556
rect 58210 27518 58262 27556
rect 58262 27518 58264 27556
rect 58856 65914 58912 65916
rect 58856 65862 58858 65914
rect 58858 65862 58910 65914
rect 58910 65862 58912 65914
rect 58856 65860 58912 65862
rect 58980 65914 59036 65916
rect 58980 65862 58982 65914
rect 58982 65862 59034 65914
rect 59034 65862 59036 65914
rect 58980 65860 59036 65862
rect 59104 65914 59160 65916
rect 59104 65862 59106 65914
rect 59106 65862 59158 65914
rect 59158 65862 59160 65914
rect 59104 65860 59160 65862
rect 59228 65914 59284 65916
rect 59228 65862 59230 65914
rect 59230 65862 59282 65914
rect 59282 65862 59284 65914
rect 59228 65860 59284 65862
rect 59352 65914 59408 65916
rect 59352 65862 59354 65914
rect 59354 65862 59406 65914
rect 59406 65862 59408 65914
rect 59352 65860 59408 65862
rect 58856 65790 58912 65792
rect 58856 65738 58858 65790
rect 58858 65738 58910 65790
rect 58910 65738 58912 65790
rect 58856 65736 58912 65738
rect 58980 65790 59036 65792
rect 58980 65738 58982 65790
rect 58982 65738 59034 65790
rect 59034 65738 59036 65790
rect 58980 65736 59036 65738
rect 59104 65790 59160 65792
rect 59104 65738 59106 65790
rect 59106 65738 59158 65790
rect 59158 65738 59160 65790
rect 59104 65736 59160 65738
rect 59228 65790 59284 65792
rect 59228 65738 59230 65790
rect 59230 65738 59282 65790
rect 59282 65738 59284 65790
rect 59228 65736 59284 65738
rect 59352 65790 59408 65792
rect 59352 65738 59354 65790
rect 59354 65738 59406 65790
rect 59406 65738 59408 65790
rect 59352 65736 59408 65738
rect 58822 34979 58878 34981
rect 58822 34927 58824 34979
rect 58824 34927 58876 34979
rect 58876 34927 58878 34979
rect 58822 34925 58878 34927
rect 58946 34979 59002 34981
rect 58946 34927 58948 34979
rect 58948 34927 59000 34979
rect 59000 34927 59002 34979
rect 58946 34925 59002 34927
rect 59070 34979 59126 34981
rect 59070 34927 59072 34979
rect 59072 34927 59124 34979
rect 59124 34927 59126 34979
rect 59070 34925 59126 34927
rect 59194 34979 59250 34981
rect 59194 34927 59196 34979
rect 59196 34927 59248 34979
rect 59248 34927 59250 34979
rect 59194 34925 59250 34927
rect 59318 34979 59374 34981
rect 59318 34927 59320 34979
rect 59320 34927 59372 34979
rect 59372 34927 59374 34979
rect 59318 34925 59374 34927
rect 59442 34979 59498 34981
rect 59442 34927 59444 34979
rect 59444 34927 59496 34979
rect 59496 34927 59498 34979
rect 59442 34925 59498 34927
rect 58822 34855 58878 34857
rect 58822 34803 58824 34855
rect 58824 34803 58876 34855
rect 58876 34803 58878 34855
rect 58822 34801 58878 34803
rect 58946 34855 59002 34857
rect 58946 34803 58948 34855
rect 58948 34803 59000 34855
rect 59000 34803 59002 34855
rect 58946 34801 59002 34803
rect 59070 34855 59126 34857
rect 59070 34803 59072 34855
rect 59072 34803 59124 34855
rect 59124 34803 59126 34855
rect 59070 34801 59126 34803
rect 59194 34855 59250 34857
rect 59194 34803 59196 34855
rect 59196 34803 59248 34855
rect 59248 34803 59250 34855
rect 59194 34801 59250 34803
rect 59318 34855 59374 34857
rect 59318 34803 59320 34855
rect 59320 34803 59372 34855
rect 59372 34803 59374 34855
rect 59318 34801 59374 34803
rect 59442 34855 59498 34857
rect 59442 34803 59444 34855
rect 59444 34803 59496 34855
rect 59496 34803 59498 34855
rect 59442 34801 59498 34803
rect 58822 34731 58878 34733
rect 58822 34679 58824 34731
rect 58824 34679 58876 34731
rect 58876 34679 58878 34731
rect 58822 34677 58878 34679
rect 58946 34731 59002 34733
rect 58946 34679 58948 34731
rect 58948 34679 59000 34731
rect 59000 34679 59002 34731
rect 58946 34677 59002 34679
rect 59070 34731 59126 34733
rect 59070 34679 59072 34731
rect 59072 34679 59124 34731
rect 59124 34679 59126 34731
rect 59070 34677 59126 34679
rect 59194 34731 59250 34733
rect 59194 34679 59196 34731
rect 59196 34679 59248 34731
rect 59248 34679 59250 34731
rect 59194 34677 59250 34679
rect 59318 34731 59374 34733
rect 59318 34679 59320 34731
rect 59320 34679 59372 34731
rect 59372 34679 59374 34731
rect 59318 34677 59374 34679
rect 59442 34731 59498 34733
rect 59442 34679 59444 34731
rect 59444 34679 59496 34731
rect 59496 34679 59498 34731
rect 59442 34677 59498 34679
rect 58873 31242 58929 31298
rect 58997 31242 59053 31298
rect 59121 31242 59177 31298
rect 59245 31242 59301 31298
rect 59369 31242 59425 31298
rect 58873 31118 58929 31174
rect 58997 31118 59053 31174
rect 59121 31118 59177 31174
rect 59245 31118 59301 31174
rect 59369 31118 59425 31174
rect 58873 30994 58929 31050
rect 58997 30994 59053 31050
rect 59121 30994 59177 31050
rect 59245 30994 59301 31050
rect 59369 30994 59425 31050
rect 58873 30797 58929 30853
rect 58997 30797 59053 30853
rect 59121 30797 59177 30853
rect 59245 30797 59301 30853
rect 59369 30797 59425 30853
rect 58873 30673 58929 30729
rect 58997 30673 59053 30729
rect 59121 30673 59177 30729
rect 59245 30673 59301 30729
rect 59369 30673 59425 30729
rect 58873 30549 58929 30605
rect 58997 30549 59053 30605
rect 59121 30549 59177 30605
rect 59245 30549 59301 30605
rect 59369 30549 59425 30605
rect 58859 28265 58915 28321
rect 58983 28265 59039 28321
rect 59107 28265 59163 28321
rect 59231 28265 59287 28321
rect 59355 28265 59411 28321
rect 58859 28141 58915 28197
rect 58983 28141 59039 28197
rect 59107 28141 59163 28197
rect 59231 28141 59287 28197
rect 59355 28141 59411 28197
rect 58859 28017 58915 28073
rect 58983 28017 59039 28073
rect 59107 28017 59163 28073
rect 59231 28017 59287 28073
rect 59355 28017 59411 28073
rect 58859 27893 58915 27949
rect 58983 27893 59039 27949
rect 59107 27893 59163 27949
rect 59231 27893 59287 27949
rect 59355 27893 59411 27949
rect 58859 27769 58915 27825
rect 58983 27769 59039 27825
rect 59107 27769 59163 27825
rect 59231 27769 59287 27825
rect 59355 27769 59411 27825
rect 58859 27645 58915 27701
rect 58983 27645 59039 27701
rect 59107 27645 59163 27701
rect 59231 27645 59287 27701
rect 59355 27645 59411 27701
rect 58859 27521 58915 27577
rect 58983 27521 59039 27577
rect 59107 27521 59163 27577
rect 59231 27521 59287 27577
rect 59355 27521 59411 27577
rect 58859 27397 58915 27453
rect 58983 27397 59039 27453
rect 59107 27397 59163 27453
rect 59231 27397 59287 27453
rect 59355 27397 59411 27453
rect 58859 27273 58915 27329
rect 58983 27273 59039 27329
rect 59107 27273 59163 27329
rect 59231 27273 59287 27329
rect 59355 27273 59411 27329
rect 58859 27149 58915 27205
rect 58983 27149 59039 27205
rect 59107 27149 59163 27205
rect 59231 27149 59287 27205
rect 59355 27149 59411 27205
rect 58859 27025 58915 27081
rect 58983 27025 59039 27081
rect 59107 27025 59163 27081
rect 59231 27025 59287 27081
rect 59355 27025 59411 27081
rect 58859 26901 58915 26957
rect 58983 26901 59039 26957
rect 59107 26901 59163 26957
rect 59231 26901 59287 26957
rect 59355 26901 59411 26957
rect 58859 26777 58915 26833
rect 58983 26777 59039 26833
rect 59107 26777 59163 26833
rect 59231 26777 59287 26833
rect 59355 26777 59411 26833
rect 58859 26653 58915 26709
rect 58983 26653 59039 26709
rect 59107 26653 59163 26709
rect 59231 26653 59287 26709
rect 59355 26653 59411 26709
rect 58859 26529 58915 26585
rect 58983 26529 59039 26585
rect 59107 26529 59163 26585
rect 59231 26529 59287 26585
rect 59355 26529 59411 26585
rect 57994 24074 58258 24075
rect 57994 24022 57998 24074
rect 57998 24022 58050 24074
rect 58050 24022 58210 24074
rect 58210 24022 58258 24074
rect 57994 23857 58258 24022
rect 57994 23805 57998 23857
rect 57998 23805 58050 23857
rect 58050 23805 58210 23857
rect 58210 23805 58258 23857
rect 57994 23639 58258 23805
rect 57994 23587 57998 23639
rect 57998 23587 58050 23639
rect 58050 23587 58210 23639
rect 58210 23587 58258 23639
rect 57994 23421 58258 23587
rect 57994 23369 57998 23421
rect 57998 23369 58050 23421
rect 58050 23369 58210 23421
rect 58210 23369 58258 23421
rect 57994 23204 58258 23369
rect 57994 23187 57998 23204
rect 57998 23187 58050 23204
rect 58050 23187 58210 23204
rect 58210 23187 58258 23204
rect 58048 20540 58050 20570
rect 58050 20540 58208 20570
rect 58048 20410 58208 20540
rect 58048 20157 58208 20226
rect 58048 20105 58050 20157
rect 58050 20105 58208 20157
rect 58048 20066 58208 20105
rect 57996 13734 58052 13790
rect 58208 13734 58264 13790
rect 57996 13517 58052 13573
rect 58208 13517 58264 13573
rect 57996 13299 58052 13355
rect 58208 13299 58264 13355
rect 57996 13082 58052 13138
rect 58208 13082 58264 13138
rect 57996 12864 58052 12920
rect 58208 12864 58264 12920
rect 57996 12646 58052 12702
rect 58208 12646 58264 12702
rect 57996 12428 58052 12484
rect 58208 12428 58264 12484
rect 57996 12211 58052 12267
rect 58208 12211 58264 12267
rect 57996 11993 58052 12049
rect 58208 11993 58264 12049
rect 57996 11776 58052 11832
rect 58208 11776 58264 11832
rect 57996 9351 58052 9407
rect 58208 9351 58264 9407
rect 57996 9134 58052 9190
rect 58208 9134 58264 9190
rect 57996 8916 58052 8972
rect 58208 8916 58264 8972
rect 57996 8698 58052 8754
rect 58208 8698 58264 8754
rect 57996 8480 58052 8536
rect 58208 8480 58264 8536
rect 57996 8263 58052 8319
rect 58208 8263 58264 8319
rect 57996 5523 57998 5539
rect 57998 5523 58050 5539
rect 58050 5523 58052 5539
rect 57996 5483 58052 5523
rect 58208 5523 58210 5539
rect 58210 5523 58262 5539
rect 58262 5523 58264 5539
rect 58208 5483 58264 5523
rect 57996 5306 57998 5321
rect 57998 5306 58050 5321
rect 58050 5306 58052 5321
rect 57996 5265 58052 5306
rect 58208 5306 58210 5321
rect 58210 5306 58262 5321
rect 58262 5306 58264 5321
rect 58208 5265 58264 5306
rect 61287 5323 61289 5462
rect 61289 5323 61445 5462
rect 61445 5323 61447 5462
rect 61287 5302 61447 5323
rect 57996 4472 58052 4528
rect 58208 4472 58264 4528
rect 57996 4254 58052 4310
rect 58208 4254 58264 4310
<< metal3 >>
rect 1401 67376 2401 68176
rect 2626 67568 3626 68176
rect 4137 67376 5137 68176
rect 5362 67568 6362 68176
rect 6801 67376 7801 68176
rect 8026 67568 9026 68176
rect 9537 67376 10537 68176
rect 10762 67568 11762 68176
rect 12201 67376 13201 68176
rect 13426 67568 14426 68176
rect 14937 67376 15937 68176
rect 16162 67568 17162 68176
rect 17601 67376 18601 68176
rect 18826 67568 19826 68176
rect 20653 67376 21653 68176
rect 22258 67568 23258 68176
rect 23483 67376 24483 68176
rect 25158 67568 26158 68176
rect 26572 67376 27572 68176
rect 27877 67568 28877 68176
rect 29273 67568 30273 68176
rect 30710 67376 31710 68176
rect 32381 67568 33381 68176
rect 34024 67568 35024 68176
rect 35415 67376 36415 68176
rect 36948 67568 37948 68176
rect 38585 67376 39585 68176
rect 39882 67568 40882 68176
rect 41230 67376 42230 68176
rect 42430 67568 43430 68176
rect 43713 67568 44713 68176
rect 45069 67376 46069 68176
rect 46313 67376 47313 68176
rect 47538 67568 48538 68176
rect 48901 67376 49901 68176
rect 50465 67568 51465 68176
rect 52569 67376 53569 68176
rect 54262 67376 55262 68176
rect 55990 67568 56990 68176
rect 57547 67376 58547 68176
rect 58791 67568 59791 68176
rect 60977 67376 61977 68176
rect 62202 67568 63202 68176
rect 63713 67376 64713 68176
rect 64938 67568 65938 68176
rect 66377 67568 67378 68176
rect 67602 67568 68603 68176
rect 66378 67376 67378 67568
rect 69113 67376 70113 68176
rect 70338 67568 71338 68176
rect 71777 67376 72777 68176
rect 73002 67568 74002 68176
rect 74513 67376 75513 68176
rect 75738 67568 76738 68176
rect 77177 67376 78177 68176
rect 78402 67568 79402 68176
rect 80229 67376 81229 68176
rect 81834 67568 82834 68176
rect 83059 67376 84059 68176
rect 84666 67376 85666 68176
rect 0 66376 86372 67376
rect 0 65976 1014 66176
rect 85358 65976 86372 66176
rect 0 65928 27272 65976
rect 0 65926 57494 65928
rect 60471 65926 86372 65976
rect 0 65916 86372 65926
rect 0 65860 25378 65916
rect 25434 65860 25502 65916
rect 25558 65860 25626 65916
rect 25682 65860 25750 65916
rect 25806 65860 25874 65916
rect 25930 65860 58856 65916
rect 58912 65860 58980 65916
rect 59036 65860 59104 65916
rect 59160 65860 59228 65916
rect 59284 65860 59352 65916
rect 59408 65860 86372 65916
rect 0 65855 86372 65860
rect 0 65799 27788 65855
rect 27844 65799 27999 65855
rect 28055 65799 28210 65855
rect 28266 65799 28421 65855
rect 28477 65799 28632 65855
rect 28688 65799 28843 65855
rect 28899 65799 29054 65855
rect 29110 65799 34288 65855
rect 34344 65799 34499 65855
rect 34555 65799 34710 65855
rect 34766 65799 34921 65855
rect 34977 65799 40250 65855
rect 40306 65799 40430 65855
rect 40486 65799 50135 65855
rect 50191 65799 50346 65855
rect 50402 65799 50557 65855
rect 50613 65799 50768 65855
rect 50824 65799 56013 65855
rect 56069 65799 56224 65855
rect 56280 65799 56435 65855
rect 56491 65799 56646 65855
rect 56702 65799 56857 65855
rect 56913 65799 57068 65855
rect 57124 65799 57279 65855
rect 57335 65799 86372 65855
rect 0 65792 86372 65799
rect 0 65736 25378 65792
rect 25434 65736 25502 65792
rect 25558 65736 25626 65792
rect 25682 65736 25750 65792
rect 25806 65736 25874 65792
rect 25930 65736 58856 65792
rect 58912 65736 58980 65792
rect 59036 65736 59104 65792
rect 59160 65736 59228 65792
rect 59284 65736 59352 65792
rect 59408 65736 86372 65792
rect 0 65727 86372 65736
rect 0 65726 27779 65727
rect 30402 65726 54622 65727
rect 57410 65726 86372 65727
rect 0 65676 27272 65726
rect 60471 65676 86372 65726
rect 0 65476 1014 65676
rect 85358 65476 86372 65676
rect 28677 65434 33984 65468
rect 28676 65374 33984 65434
rect 28676 65318 33048 65374
rect 33104 65318 33259 65374
rect 33315 65318 33470 65374
rect 33526 65318 33681 65374
rect 33737 65318 33892 65374
rect 33948 65318 33984 65374
rect 28676 65300 33984 65318
rect 0 64576 1706 65276
rect 28677 65266 33984 65300
rect 36863 65372 42155 65411
rect 36863 65316 36899 65372
rect 36955 65316 37110 65372
rect 37166 65316 37321 65372
rect 37377 65316 37532 65372
rect 37588 65316 41008 65372
rect 41064 65316 41219 65372
rect 41275 65316 41430 65372
rect 41486 65316 41641 65372
rect 41697 65316 41852 65372
rect 41908 65316 42062 65372
rect 42118 65316 42155 65372
rect 42671 65365 43222 65404
rect 42671 65330 42708 65365
rect 36863 65277 42155 65316
rect 42670 65309 42708 65330
rect 42764 65309 42919 65365
rect 42975 65309 43130 65365
rect 43186 65309 43222 65365
rect 42670 65271 43222 65309
rect 51042 65372 61644 65468
rect 51042 65316 51079 65372
rect 51135 65316 51290 65372
rect 51346 65316 51501 65372
rect 51557 65316 51712 65372
rect 51768 65316 51923 65372
rect 51979 65316 61644 65372
rect 42670 65028 42769 65271
rect 51042 65266 61644 65316
rect 24298 64955 60825 65028
rect 24298 64899 29580 64955
rect 29636 64899 29791 64955
rect 29847 64899 30003 64955
rect 30059 64899 30214 64955
rect 30270 64899 30852 64955
rect 30908 64899 31063 64955
rect 31119 64899 31274 64955
rect 31330 64899 31484 64955
rect 31540 64899 31695 64955
rect 31751 64899 31907 64955
rect 31963 64899 32118 64955
rect 32174 64899 32328 64955
rect 32384 64899 32539 64955
rect 32595 64899 32750 64955
rect 32806 64899 35218 64955
rect 35274 64899 35428 64955
rect 35484 64899 35639 64955
rect 35695 64899 35851 64955
rect 35907 64899 36062 64955
rect 36118 64899 36272 64955
rect 36328 64899 39050 64955
rect 39106 64899 39230 64955
rect 39286 64899 40777 64955
rect 40833 64899 40988 64955
rect 41044 64899 41199 64955
rect 41255 64954 44832 64955
rect 41255 64899 41881 64954
rect 24298 64898 41881 64899
rect 42041 64899 44832 64954
rect 44888 64899 45043 64955
rect 45099 64899 45254 64955
rect 45310 64899 48836 64955
rect 48892 64899 49046 64955
rect 49102 64899 49257 64955
rect 49313 64899 49469 64955
rect 49525 64899 49680 64955
rect 49736 64899 49890 64955
rect 49946 64899 52314 64955
rect 52370 64899 52525 64955
rect 52581 64899 52736 64955
rect 52792 64899 52946 64955
rect 53002 64899 53157 64955
rect 53213 64899 53369 64955
rect 53425 64899 53580 64955
rect 53636 64899 53790 64955
rect 53846 64899 54001 64955
rect 54057 64899 54212 64955
rect 54268 64899 54853 64955
rect 54909 64899 55064 64955
rect 55120 64899 55276 64955
rect 55332 64899 55487 64955
rect 55543 64899 60825 64955
rect 42041 64898 60825 64899
rect 24298 64827 60825 64898
rect 30403 64826 54622 64827
rect 36648 64601 40041 64602
rect 24298 64522 34090 64588
rect 24298 64466 33055 64522
rect 33111 64466 33235 64522
rect 33291 64515 34090 64522
rect 33291 64466 33817 64515
rect 24298 64459 33817 64466
rect 33873 64459 33997 64515
rect 34053 64459 34090 64515
rect 36640 64563 40085 64601
rect 36640 64507 36676 64563
rect 36732 64507 39992 64563
rect 40048 64507 40085 64563
rect 36640 64468 40085 64507
rect 48557 64549 48687 64588
rect 48557 64493 48594 64549
rect 48650 64493 48687 64549
rect 24298 64387 34090 64459
rect 30403 64386 34090 64387
rect 0 64176 1014 64376
rect 48557 64370 48687 64493
rect 51034 64515 60825 64588
rect 84666 64576 86372 65276
rect 51034 64459 51071 64515
rect 51127 64459 51251 64515
rect 51307 64459 51833 64515
rect 51889 64459 52013 64515
rect 52069 64459 60825 64515
rect 51034 64387 60825 64459
rect 51034 64386 54622 64387
rect 37852 64332 48687 64370
rect 37852 64276 37889 64332
rect 37945 64276 38069 64332
rect 38125 64276 39773 64332
rect 39829 64331 48687 64332
rect 39829 64276 48594 64331
rect 37852 64275 48594 64276
rect 48650 64275 48687 64331
rect 37852 64237 48687 64275
rect 85358 64176 86372 64376
rect 0 64128 27272 64176
rect 60471 64128 86372 64176
rect 0 64055 86372 64128
rect 0 63999 27788 64055
rect 27844 63999 27999 64055
rect 28055 63999 28210 64055
rect 28266 63999 28421 64055
rect 28477 63999 28632 64055
rect 28688 63999 28843 64055
rect 28899 63999 29054 64055
rect 29110 63999 34282 64055
rect 34338 63999 34493 64055
rect 34549 63999 34705 64055
rect 34761 63999 34916 64055
rect 34972 63999 38328 64055
rect 38384 63999 38539 64055
rect 38595 63999 38750 64055
rect 38806 63999 40251 64055
rect 40307 63999 40431 64055
rect 40487 63999 43788 64055
rect 43844 63999 43999 64055
rect 44055 63999 44211 64055
rect 44267 63999 44422 64055
rect 44478 63999 50161 64055
rect 50217 63999 50372 64055
rect 50428 63999 50584 64055
rect 50640 63999 50795 64055
rect 50851 63999 56013 64055
rect 56069 63999 56224 64055
rect 56280 63999 56435 64055
rect 56491 63999 56646 64055
rect 56702 63999 56857 64055
rect 56913 63999 57068 64055
rect 57124 63999 57279 64055
rect 57335 63999 86372 64055
rect 0 63927 86372 63999
rect 0 63876 27272 63927
rect 30403 63926 54622 63927
rect 60471 63876 86372 63927
rect 0 63676 1014 63876
rect 37852 63779 48687 63817
rect 37852 63778 48594 63779
rect 37852 63722 37889 63778
rect 37945 63722 38069 63778
rect 38125 63722 39773 63778
rect 39829 63723 48594 63778
rect 48650 63723 48687 63779
rect 39829 63722 48687 63723
rect 37852 63684 48687 63722
rect 24298 63595 34090 63668
rect 24298 63588 33817 63595
rect 24298 63532 33055 63588
rect 33111 63532 33235 63588
rect 33291 63539 33817 63588
rect 33873 63539 33997 63595
rect 34053 63539 34090 63595
rect 33291 63532 34090 63539
rect 0 62776 1706 63476
rect 24298 63466 34090 63532
rect 36640 63547 40085 63586
rect 36640 63491 36676 63547
rect 36732 63491 39992 63547
rect 40048 63491 40085 63547
rect 36640 63453 40085 63491
rect 48557 63561 48687 63684
rect 85358 63676 86372 63876
rect 48557 63505 48594 63561
rect 48650 63505 48687 63561
rect 48557 63466 48687 63505
rect 51034 63595 60825 63668
rect 51034 63539 51071 63595
rect 51127 63539 51251 63595
rect 51307 63539 51833 63595
rect 51889 63539 52013 63595
rect 52069 63539 60825 63595
rect 51034 63466 60825 63539
rect 36648 63452 40041 63453
rect 24298 63155 60825 63228
rect 24298 63099 29580 63155
rect 29636 63099 29791 63155
rect 29847 63099 30003 63155
rect 30059 63099 30214 63155
rect 30270 63099 30852 63155
rect 30908 63099 31063 63155
rect 31119 63099 31274 63155
rect 31330 63099 31484 63155
rect 31540 63099 31695 63155
rect 31751 63099 31907 63155
rect 31963 63099 32118 63155
rect 32174 63099 32328 63155
rect 32384 63099 32539 63155
rect 32595 63099 32750 63155
rect 32806 63099 35218 63155
rect 35274 63099 35428 63155
rect 35484 63099 35639 63155
rect 35695 63099 35851 63155
rect 35907 63099 36062 63155
rect 36118 63099 36272 63155
rect 36328 63099 39050 63155
rect 39106 63099 39230 63155
rect 39286 63099 44832 63155
rect 44888 63099 45043 63155
rect 45099 63099 45254 63155
rect 45310 63099 48836 63155
rect 48892 63099 49046 63155
rect 49102 63099 49257 63155
rect 49313 63099 49469 63155
rect 49525 63099 49680 63155
rect 49736 63099 49890 63155
rect 49946 63099 52314 63155
rect 52370 63099 52525 63155
rect 52581 63099 52736 63155
rect 52792 63099 52946 63155
rect 53002 63099 53157 63155
rect 53213 63099 53369 63155
rect 53425 63099 53580 63155
rect 53636 63099 53790 63155
rect 53846 63099 54001 63155
rect 54057 63099 54212 63155
rect 54268 63099 54853 63155
rect 54909 63099 55064 63155
rect 55120 63099 55276 63155
rect 55332 63099 55487 63155
rect 55543 63099 60825 63155
rect 24298 63027 60825 63099
rect 30403 63026 54622 63027
rect 36648 62801 40041 62802
rect 24298 62722 34090 62788
rect 24298 62666 33055 62722
rect 33111 62666 33235 62722
rect 33291 62715 34090 62722
rect 33291 62666 33817 62715
rect 24298 62659 33817 62666
rect 33873 62659 33997 62715
rect 34053 62659 34090 62715
rect 36640 62763 40085 62801
rect 36640 62707 36676 62763
rect 36732 62707 39992 62763
rect 40048 62707 40085 62763
rect 36640 62668 40085 62707
rect 48557 62749 48687 62788
rect 48557 62693 48594 62749
rect 48650 62693 48687 62749
rect 24298 62587 34090 62659
rect 30403 62586 34090 62587
rect 0 62376 1014 62576
rect 48557 62570 48687 62693
rect 51034 62715 60825 62788
rect 84666 62776 86372 63476
rect 51034 62659 51071 62715
rect 51127 62659 51251 62715
rect 51307 62659 51833 62715
rect 51889 62659 52013 62715
rect 52069 62659 60825 62715
rect 51034 62587 60825 62659
rect 51034 62586 54622 62587
rect 37852 62532 48687 62570
rect 37852 62476 37889 62532
rect 37945 62476 38069 62532
rect 38125 62476 39773 62532
rect 39829 62531 48687 62532
rect 39829 62476 48594 62531
rect 37852 62475 48594 62476
rect 48650 62475 48687 62531
rect 37852 62437 48687 62475
rect 85358 62376 86372 62576
rect 0 62328 27272 62376
rect 60471 62328 86372 62376
rect 0 62255 86372 62328
rect 0 62199 27788 62255
rect 27844 62199 27999 62255
rect 28055 62199 28210 62255
rect 28266 62199 28421 62255
rect 28477 62199 28632 62255
rect 28688 62199 28843 62255
rect 28899 62199 29054 62255
rect 29110 62199 34282 62255
rect 34338 62199 34493 62255
rect 34549 62199 34705 62255
rect 34761 62199 34916 62255
rect 34972 62199 38328 62255
rect 38384 62199 38539 62255
rect 38595 62199 38750 62255
rect 38806 62199 40251 62255
rect 40307 62199 40431 62255
rect 40487 62199 43788 62255
rect 43844 62199 43999 62255
rect 44055 62199 44211 62255
rect 44267 62199 44422 62255
rect 44478 62199 50161 62255
rect 50217 62199 50372 62255
rect 50428 62199 50584 62255
rect 50640 62199 50795 62255
rect 50851 62199 56013 62255
rect 56069 62199 56224 62255
rect 56280 62199 56435 62255
rect 56491 62199 56646 62255
rect 56702 62199 56857 62255
rect 56913 62199 57068 62255
rect 57124 62199 57279 62255
rect 57335 62199 86372 62255
rect 0 62127 86372 62199
rect 0 62076 27272 62127
rect 30403 62126 54622 62127
rect 60471 62076 86372 62127
rect 0 61876 1014 62076
rect 37852 61979 48687 62017
rect 37852 61978 48594 61979
rect 37852 61922 37889 61978
rect 37945 61922 38069 61978
rect 38125 61922 39773 61978
rect 39829 61923 48594 61978
rect 48650 61923 48687 61979
rect 39829 61922 48687 61923
rect 37852 61884 48687 61922
rect 24298 61795 34090 61868
rect 24298 61788 33817 61795
rect 24298 61732 33055 61788
rect 33111 61732 33235 61788
rect 33291 61739 33817 61788
rect 33873 61739 33997 61795
rect 34053 61739 34090 61795
rect 33291 61732 34090 61739
rect 0 60976 1706 61676
rect 24298 61666 34090 61732
rect 36640 61747 40085 61786
rect 36640 61691 36676 61747
rect 36732 61691 39992 61747
rect 40048 61691 40085 61747
rect 36640 61653 40085 61691
rect 48557 61761 48687 61884
rect 85358 61876 86372 62076
rect 48557 61705 48594 61761
rect 48650 61705 48687 61761
rect 48557 61666 48687 61705
rect 51034 61795 60825 61868
rect 51034 61739 51071 61795
rect 51127 61739 51251 61795
rect 51307 61739 51833 61795
rect 51889 61739 52013 61795
rect 52069 61739 60825 61795
rect 51034 61666 60825 61739
rect 36648 61652 40041 61653
rect 24298 61355 60825 61428
rect 24298 61299 29580 61355
rect 29636 61299 29791 61355
rect 29847 61299 30003 61355
rect 30059 61299 30214 61355
rect 30270 61299 30852 61355
rect 30908 61299 31063 61355
rect 31119 61299 31274 61355
rect 31330 61299 31484 61355
rect 31540 61299 31695 61355
rect 31751 61299 31907 61355
rect 31963 61299 32118 61355
rect 32174 61299 32328 61355
rect 32384 61299 32539 61355
rect 32595 61299 32750 61355
rect 32806 61299 35218 61355
rect 35274 61299 35428 61355
rect 35484 61299 35639 61355
rect 35695 61299 35851 61355
rect 35907 61299 36062 61355
rect 36118 61299 36272 61355
rect 36328 61299 39050 61355
rect 39106 61299 39230 61355
rect 39286 61299 44832 61355
rect 44888 61299 45043 61355
rect 45099 61299 45254 61355
rect 45310 61299 48836 61355
rect 48892 61299 49046 61355
rect 49102 61299 49257 61355
rect 49313 61299 49469 61355
rect 49525 61299 49680 61355
rect 49736 61299 49890 61355
rect 49946 61299 52314 61355
rect 52370 61299 52525 61355
rect 52581 61299 52736 61355
rect 52792 61299 52946 61355
rect 53002 61299 53157 61355
rect 53213 61299 53369 61355
rect 53425 61299 53580 61355
rect 53636 61299 53790 61355
rect 53846 61299 54001 61355
rect 54057 61299 54212 61355
rect 54268 61299 54853 61355
rect 54909 61299 55064 61355
rect 55120 61299 55276 61355
rect 55332 61299 55487 61355
rect 55543 61299 60825 61355
rect 24298 61227 60825 61299
rect 30403 61226 54622 61227
rect 36648 61001 40041 61002
rect 24298 60922 34090 60988
rect 24298 60866 33055 60922
rect 33111 60866 33235 60922
rect 33291 60915 34090 60922
rect 33291 60866 33817 60915
rect 24298 60859 33817 60866
rect 33873 60859 33997 60915
rect 34053 60859 34090 60915
rect 36640 60963 40085 61001
rect 36640 60907 36676 60963
rect 36732 60907 39992 60963
rect 40048 60907 40085 60963
rect 36640 60868 40085 60907
rect 48557 60949 48687 60988
rect 48557 60893 48594 60949
rect 48650 60893 48687 60949
rect 24298 60787 34090 60859
rect 30403 60786 34090 60787
rect 0 60576 1014 60776
rect 48557 60770 48687 60893
rect 51034 60915 60825 60988
rect 84666 60976 86372 61676
rect 51034 60859 51071 60915
rect 51127 60859 51251 60915
rect 51307 60859 51833 60915
rect 51889 60859 52013 60915
rect 52069 60859 60825 60915
rect 51034 60787 60825 60859
rect 51034 60786 54622 60787
rect 37852 60732 48687 60770
rect 37852 60676 37889 60732
rect 37945 60676 38069 60732
rect 38125 60676 39773 60732
rect 39829 60731 48687 60732
rect 39829 60676 48594 60731
rect 37852 60675 48594 60676
rect 48650 60675 48687 60731
rect 37852 60637 48687 60675
rect 85358 60576 86372 60776
rect 0 60528 27272 60576
rect 60471 60528 86372 60576
rect 0 60455 86372 60528
rect 0 60399 27788 60455
rect 27844 60399 27999 60455
rect 28055 60399 28210 60455
rect 28266 60399 28421 60455
rect 28477 60399 28632 60455
rect 28688 60399 28843 60455
rect 28899 60399 29054 60455
rect 29110 60399 34282 60455
rect 34338 60399 34493 60455
rect 34549 60399 34705 60455
rect 34761 60399 34916 60455
rect 34972 60399 38328 60455
rect 38384 60399 38539 60455
rect 38595 60399 38750 60455
rect 38806 60399 40251 60455
rect 40307 60399 40431 60455
rect 40487 60399 43788 60455
rect 43844 60399 43999 60455
rect 44055 60399 44211 60455
rect 44267 60399 44422 60455
rect 44478 60399 50161 60455
rect 50217 60399 50372 60455
rect 50428 60399 50584 60455
rect 50640 60399 50795 60455
rect 50851 60399 56013 60455
rect 56069 60399 56224 60455
rect 56280 60399 56435 60455
rect 56491 60399 56646 60455
rect 56702 60399 56857 60455
rect 56913 60399 57068 60455
rect 57124 60399 57279 60455
rect 57335 60399 86372 60455
rect 0 60327 86372 60399
rect 0 60276 27272 60327
rect 30403 60326 54622 60327
rect 60471 60276 86372 60327
rect 0 60076 1014 60276
rect 37852 60179 48687 60217
rect 37852 60178 48594 60179
rect 37852 60122 37889 60178
rect 37945 60122 38069 60178
rect 38125 60122 39773 60178
rect 39829 60123 48594 60178
rect 48650 60123 48687 60179
rect 39829 60122 48687 60123
rect 37852 60084 48687 60122
rect 24298 59995 34090 60068
rect 24298 59988 33817 59995
rect 24298 59932 33055 59988
rect 33111 59932 33235 59988
rect 33291 59939 33817 59988
rect 33873 59939 33997 59995
rect 34053 59939 34090 59995
rect 33291 59932 34090 59939
rect 0 59176 1706 59876
rect 24298 59866 34090 59932
rect 36640 59947 40085 59986
rect 36640 59891 36676 59947
rect 36732 59891 39992 59947
rect 40048 59891 40085 59947
rect 36640 59853 40085 59891
rect 48557 59961 48687 60084
rect 85358 60076 86372 60276
rect 48557 59905 48594 59961
rect 48650 59905 48687 59961
rect 48557 59866 48687 59905
rect 51034 59995 60825 60068
rect 51034 59939 51071 59995
rect 51127 59939 51251 59995
rect 51307 59939 51833 59995
rect 51889 59939 52013 59995
rect 52069 59939 60825 59995
rect 51034 59866 60825 59939
rect 36648 59852 40041 59853
rect 24298 59555 60825 59628
rect 24298 59499 29580 59555
rect 29636 59499 29791 59555
rect 29847 59499 30003 59555
rect 30059 59499 30214 59555
rect 30270 59499 30852 59555
rect 30908 59499 31063 59555
rect 31119 59499 31274 59555
rect 31330 59499 31484 59555
rect 31540 59499 31695 59555
rect 31751 59499 31907 59555
rect 31963 59499 32118 59555
rect 32174 59499 32328 59555
rect 32384 59499 32539 59555
rect 32595 59499 32750 59555
rect 32806 59499 35218 59555
rect 35274 59499 35428 59555
rect 35484 59499 35639 59555
rect 35695 59499 35851 59555
rect 35907 59499 36062 59555
rect 36118 59499 36272 59555
rect 36328 59499 39050 59555
rect 39106 59499 39230 59555
rect 39286 59499 44832 59555
rect 44888 59499 45043 59555
rect 45099 59499 45254 59555
rect 45310 59499 48836 59555
rect 48892 59499 49046 59555
rect 49102 59499 49257 59555
rect 49313 59499 49469 59555
rect 49525 59499 49680 59555
rect 49736 59499 49890 59555
rect 49946 59499 52314 59555
rect 52370 59499 52525 59555
rect 52581 59499 52736 59555
rect 52792 59499 52946 59555
rect 53002 59499 53157 59555
rect 53213 59499 53369 59555
rect 53425 59499 53580 59555
rect 53636 59499 53790 59555
rect 53846 59499 54001 59555
rect 54057 59499 54212 59555
rect 54268 59499 54853 59555
rect 54909 59499 55064 59555
rect 55120 59499 55276 59555
rect 55332 59499 55487 59555
rect 55543 59499 60825 59555
rect 24298 59427 60825 59499
rect 30403 59426 54622 59427
rect 36648 59201 40041 59202
rect 24298 59122 34090 59188
rect 24298 59066 33055 59122
rect 33111 59066 33235 59122
rect 33291 59115 34090 59122
rect 33291 59066 33817 59115
rect 24298 59059 33817 59066
rect 33873 59059 33997 59115
rect 34053 59059 34090 59115
rect 36640 59163 40085 59201
rect 36640 59107 36676 59163
rect 36732 59107 39992 59163
rect 40048 59107 40085 59163
rect 36640 59068 40085 59107
rect 48557 59149 48687 59188
rect 48557 59093 48594 59149
rect 48650 59093 48687 59149
rect 24298 58987 34090 59059
rect 30403 58986 34090 58987
rect 0 58776 1014 58976
rect 48557 58970 48687 59093
rect 51034 59115 60825 59188
rect 84666 59176 86372 59876
rect 51034 59059 51071 59115
rect 51127 59059 51251 59115
rect 51307 59059 51833 59115
rect 51889 59059 52013 59115
rect 52069 59059 60825 59115
rect 51034 58987 60825 59059
rect 51034 58986 54622 58987
rect 37852 58932 48687 58970
rect 37852 58876 37889 58932
rect 37945 58876 38069 58932
rect 38125 58876 39773 58932
rect 39829 58931 48687 58932
rect 39829 58876 48594 58931
rect 37852 58875 48594 58876
rect 48650 58875 48687 58931
rect 37852 58837 48687 58875
rect 85358 58776 86372 58976
rect 0 58728 27272 58776
rect 60471 58728 86372 58776
rect 0 58655 86372 58728
rect 0 58599 27788 58655
rect 27844 58599 27999 58655
rect 28055 58599 28210 58655
rect 28266 58599 28421 58655
rect 28477 58599 28632 58655
rect 28688 58599 28843 58655
rect 28899 58599 29054 58655
rect 29110 58599 34282 58655
rect 34338 58599 34493 58655
rect 34549 58599 34705 58655
rect 34761 58599 34916 58655
rect 34972 58599 38328 58655
rect 38384 58599 38539 58655
rect 38595 58599 38750 58655
rect 38806 58599 40251 58655
rect 40307 58599 40431 58655
rect 40487 58599 43788 58655
rect 43844 58599 43999 58655
rect 44055 58599 44211 58655
rect 44267 58599 44422 58655
rect 44478 58599 50161 58655
rect 50217 58599 50372 58655
rect 50428 58599 50584 58655
rect 50640 58599 50795 58655
rect 50851 58599 56013 58655
rect 56069 58599 56224 58655
rect 56280 58599 56435 58655
rect 56491 58599 56646 58655
rect 56702 58599 56857 58655
rect 56913 58599 57068 58655
rect 57124 58599 57279 58655
rect 57335 58599 86372 58655
rect 0 58527 86372 58599
rect 0 58476 27272 58527
rect 30403 58526 54622 58527
rect 60471 58476 86372 58527
rect 0 58276 1014 58476
rect 37852 58379 48687 58417
rect 37852 58378 48594 58379
rect 37852 58322 37889 58378
rect 37945 58322 38069 58378
rect 38125 58322 39773 58378
rect 39829 58323 48594 58378
rect 48650 58323 48687 58379
rect 39829 58322 48687 58323
rect 37852 58284 48687 58322
rect 24298 58195 34090 58268
rect 24298 58188 33817 58195
rect 24298 58132 33055 58188
rect 33111 58132 33235 58188
rect 33291 58139 33817 58188
rect 33873 58139 33997 58195
rect 34053 58139 34090 58195
rect 33291 58132 34090 58139
rect 0 57376 1706 58076
rect 24298 58066 34090 58132
rect 36640 58147 40085 58186
rect 36640 58091 36676 58147
rect 36732 58091 39992 58147
rect 40048 58091 40085 58147
rect 36640 58053 40085 58091
rect 48557 58161 48687 58284
rect 85358 58276 86372 58476
rect 48557 58105 48594 58161
rect 48650 58105 48687 58161
rect 48557 58066 48687 58105
rect 51034 58195 60825 58268
rect 51034 58139 51071 58195
rect 51127 58139 51251 58195
rect 51307 58139 51833 58195
rect 51889 58139 52013 58195
rect 52069 58139 60825 58195
rect 51034 58066 60825 58139
rect 36648 58052 40041 58053
rect 24298 57755 60825 57828
rect 24298 57699 29580 57755
rect 29636 57699 29791 57755
rect 29847 57699 30003 57755
rect 30059 57699 30214 57755
rect 30270 57699 30852 57755
rect 30908 57699 31063 57755
rect 31119 57699 31274 57755
rect 31330 57699 31484 57755
rect 31540 57699 31695 57755
rect 31751 57699 31907 57755
rect 31963 57699 32118 57755
rect 32174 57699 32328 57755
rect 32384 57699 32539 57755
rect 32595 57699 32750 57755
rect 32806 57699 35218 57755
rect 35274 57699 35428 57755
rect 35484 57699 35639 57755
rect 35695 57699 35851 57755
rect 35907 57699 36062 57755
rect 36118 57699 36272 57755
rect 36328 57699 39050 57755
rect 39106 57699 39230 57755
rect 39286 57699 44832 57755
rect 44888 57699 45043 57755
rect 45099 57699 45254 57755
rect 45310 57699 48836 57755
rect 48892 57699 49046 57755
rect 49102 57699 49257 57755
rect 49313 57699 49469 57755
rect 49525 57699 49680 57755
rect 49736 57699 49890 57755
rect 49946 57699 52314 57755
rect 52370 57699 52525 57755
rect 52581 57699 52736 57755
rect 52792 57699 52946 57755
rect 53002 57699 53157 57755
rect 53213 57699 53369 57755
rect 53425 57699 53580 57755
rect 53636 57699 53790 57755
rect 53846 57699 54001 57755
rect 54057 57699 54212 57755
rect 54268 57699 54853 57755
rect 54909 57699 55064 57755
rect 55120 57699 55276 57755
rect 55332 57699 55487 57755
rect 55543 57699 60825 57755
rect 24298 57627 60825 57699
rect 30403 57626 54622 57627
rect 36648 57401 40041 57402
rect 24298 57322 34090 57388
rect 24298 57266 33055 57322
rect 33111 57266 33235 57322
rect 33291 57315 34090 57322
rect 33291 57266 33817 57315
rect 24298 57259 33817 57266
rect 33873 57259 33997 57315
rect 34053 57259 34090 57315
rect 36640 57363 40085 57401
rect 36640 57307 36676 57363
rect 36732 57307 39992 57363
rect 40048 57307 40085 57363
rect 36640 57268 40085 57307
rect 48557 57349 48687 57388
rect 48557 57293 48594 57349
rect 48650 57293 48687 57349
rect 24298 57187 34090 57259
rect 30403 57186 34090 57187
rect 0 56976 1014 57176
rect 48557 57170 48687 57293
rect 51034 57315 60825 57388
rect 84666 57376 86372 58076
rect 51034 57259 51071 57315
rect 51127 57259 51251 57315
rect 51307 57259 51833 57315
rect 51889 57259 52013 57315
rect 52069 57259 60825 57315
rect 51034 57187 60825 57259
rect 51034 57186 54622 57187
rect 37852 57132 48687 57170
rect 37852 57076 37889 57132
rect 37945 57076 38069 57132
rect 38125 57076 39773 57132
rect 39829 57131 48687 57132
rect 39829 57076 48594 57131
rect 37852 57075 48594 57076
rect 48650 57075 48687 57131
rect 37852 57037 48687 57075
rect 85358 56976 86372 57176
rect 0 56928 27272 56976
rect 60471 56928 86372 56976
rect 0 56855 86372 56928
rect 0 56799 27788 56855
rect 27844 56799 27999 56855
rect 28055 56799 28210 56855
rect 28266 56799 28421 56855
rect 28477 56799 28632 56855
rect 28688 56799 28843 56855
rect 28899 56799 29054 56855
rect 29110 56799 34282 56855
rect 34338 56799 34493 56855
rect 34549 56799 34705 56855
rect 34761 56799 34916 56855
rect 34972 56799 38328 56855
rect 38384 56799 38539 56855
rect 38595 56799 38750 56855
rect 38806 56799 40251 56855
rect 40307 56799 40431 56855
rect 40487 56799 43788 56855
rect 43844 56799 43999 56855
rect 44055 56799 44211 56855
rect 44267 56799 44422 56855
rect 44478 56799 50161 56855
rect 50217 56799 50372 56855
rect 50428 56799 50584 56855
rect 50640 56799 50795 56855
rect 50851 56799 56013 56855
rect 56069 56799 56224 56855
rect 56280 56799 56435 56855
rect 56491 56799 56646 56855
rect 56702 56799 56857 56855
rect 56913 56799 57068 56855
rect 57124 56799 57279 56855
rect 57335 56799 86372 56855
rect 0 56727 86372 56799
rect 0 56676 27272 56727
rect 30403 56726 54622 56727
rect 60471 56676 86372 56727
rect 0 56476 1014 56676
rect 37852 56579 48687 56617
rect 37852 56578 48594 56579
rect 37852 56522 37889 56578
rect 37945 56522 38069 56578
rect 38125 56522 39773 56578
rect 39829 56523 48594 56578
rect 48650 56523 48687 56579
rect 39829 56522 48687 56523
rect 37852 56484 48687 56522
rect 24298 56395 34090 56468
rect 24298 56388 33817 56395
rect 24298 56332 33055 56388
rect 33111 56332 33235 56388
rect 33291 56339 33817 56388
rect 33873 56339 33997 56395
rect 34053 56339 34090 56395
rect 33291 56332 34090 56339
rect 0 55576 1706 56276
rect 24298 56266 34090 56332
rect 36640 56347 40085 56386
rect 36640 56291 36676 56347
rect 36732 56291 39992 56347
rect 40048 56291 40085 56347
rect 36640 56253 40085 56291
rect 48557 56361 48687 56484
rect 85358 56476 86372 56676
rect 48557 56305 48594 56361
rect 48650 56305 48687 56361
rect 48557 56266 48687 56305
rect 51034 56395 60825 56468
rect 51034 56339 51071 56395
rect 51127 56339 51251 56395
rect 51307 56339 51833 56395
rect 51889 56339 52013 56395
rect 52069 56339 60825 56395
rect 51034 56266 60825 56339
rect 36648 56252 40041 56253
rect 24298 55955 60825 56028
rect 24298 55899 29580 55955
rect 29636 55899 29791 55955
rect 29847 55899 30003 55955
rect 30059 55899 30214 55955
rect 30270 55899 30852 55955
rect 30908 55899 31063 55955
rect 31119 55899 31274 55955
rect 31330 55899 31484 55955
rect 31540 55899 31695 55955
rect 31751 55899 31907 55955
rect 31963 55899 32118 55955
rect 32174 55899 32328 55955
rect 32384 55899 32539 55955
rect 32595 55899 32750 55955
rect 32806 55899 35218 55955
rect 35274 55899 35428 55955
rect 35484 55899 35639 55955
rect 35695 55899 35851 55955
rect 35907 55899 36062 55955
rect 36118 55899 36272 55955
rect 36328 55899 39050 55955
rect 39106 55899 39230 55955
rect 39286 55899 44832 55955
rect 44888 55899 45043 55955
rect 45099 55899 45254 55955
rect 45310 55899 48836 55955
rect 48892 55899 49046 55955
rect 49102 55899 49257 55955
rect 49313 55899 49469 55955
rect 49525 55899 49680 55955
rect 49736 55899 49890 55955
rect 49946 55899 52314 55955
rect 52370 55899 52525 55955
rect 52581 55899 52736 55955
rect 52792 55899 52946 55955
rect 53002 55899 53157 55955
rect 53213 55899 53369 55955
rect 53425 55899 53580 55955
rect 53636 55899 53790 55955
rect 53846 55899 54001 55955
rect 54057 55899 54212 55955
rect 54268 55899 54853 55955
rect 54909 55899 55064 55955
rect 55120 55899 55276 55955
rect 55332 55899 55487 55955
rect 55543 55899 60825 55955
rect 24298 55827 60825 55899
rect 30403 55826 54622 55827
rect 36648 55601 40041 55602
rect 24298 55522 34090 55588
rect 24298 55466 33055 55522
rect 33111 55466 33235 55522
rect 33291 55515 34090 55522
rect 33291 55466 33817 55515
rect 24298 55459 33817 55466
rect 33873 55459 33997 55515
rect 34053 55459 34090 55515
rect 36640 55563 40085 55601
rect 36640 55507 36676 55563
rect 36732 55507 39992 55563
rect 40048 55507 40085 55563
rect 36640 55468 40085 55507
rect 48557 55549 48687 55588
rect 48557 55493 48594 55549
rect 48650 55493 48687 55549
rect 24298 55387 34090 55459
rect 30403 55386 34090 55387
rect 0 55176 1014 55376
rect 48557 55370 48687 55493
rect 51034 55515 60825 55588
rect 84666 55576 86372 56276
rect 51034 55459 51071 55515
rect 51127 55459 51251 55515
rect 51307 55459 51833 55515
rect 51889 55459 52013 55515
rect 52069 55459 60825 55515
rect 51034 55387 60825 55459
rect 51034 55386 54622 55387
rect 37852 55332 48687 55370
rect 37852 55276 37889 55332
rect 37945 55276 38069 55332
rect 38125 55276 39773 55332
rect 39829 55331 48687 55332
rect 39829 55276 48594 55331
rect 37852 55275 48594 55276
rect 48650 55275 48687 55331
rect 37852 55237 48687 55275
rect 85358 55176 86372 55376
rect 0 55128 27272 55176
rect 60471 55128 86372 55176
rect 0 55055 86372 55128
rect 0 54999 27788 55055
rect 27844 54999 27999 55055
rect 28055 54999 28210 55055
rect 28266 54999 28421 55055
rect 28477 54999 28632 55055
rect 28688 54999 28843 55055
rect 28899 54999 29054 55055
rect 29110 54999 34282 55055
rect 34338 54999 34493 55055
rect 34549 54999 34705 55055
rect 34761 54999 34916 55055
rect 34972 54999 38328 55055
rect 38384 54999 38539 55055
rect 38595 54999 38750 55055
rect 38806 54999 40251 55055
rect 40307 54999 40431 55055
rect 40487 54999 43788 55055
rect 43844 54999 43999 55055
rect 44055 54999 44211 55055
rect 44267 54999 44422 55055
rect 44478 54999 50161 55055
rect 50217 54999 50372 55055
rect 50428 54999 50584 55055
rect 50640 54999 50795 55055
rect 50851 54999 56013 55055
rect 56069 54999 56224 55055
rect 56280 54999 56435 55055
rect 56491 54999 56646 55055
rect 56702 54999 56857 55055
rect 56913 54999 57068 55055
rect 57124 54999 57279 55055
rect 57335 54999 86372 55055
rect 0 54927 86372 54999
rect 0 54876 27272 54927
rect 30403 54926 54622 54927
rect 60471 54876 86372 54927
rect 0 54676 1014 54876
rect 37852 54779 48687 54817
rect 37852 54778 48594 54779
rect 37852 54722 37889 54778
rect 37945 54722 38069 54778
rect 38125 54722 39773 54778
rect 39829 54723 48594 54778
rect 48650 54723 48687 54779
rect 39829 54722 48687 54723
rect 37852 54684 48687 54722
rect 24298 54595 34090 54668
rect 24298 54588 33817 54595
rect 24298 54532 33055 54588
rect 33111 54532 33235 54588
rect 33291 54539 33817 54588
rect 33873 54539 33997 54595
rect 34053 54539 34090 54595
rect 33291 54532 34090 54539
rect 0 53776 1706 54476
rect 24298 54466 34090 54532
rect 36640 54547 40085 54586
rect 36640 54491 36676 54547
rect 36732 54491 39992 54547
rect 40048 54491 40085 54547
rect 36640 54453 40085 54491
rect 48557 54561 48687 54684
rect 85358 54676 86372 54876
rect 48557 54505 48594 54561
rect 48650 54505 48687 54561
rect 48557 54466 48687 54505
rect 51034 54595 60825 54668
rect 51034 54539 51071 54595
rect 51127 54539 51251 54595
rect 51307 54539 51833 54595
rect 51889 54539 52013 54595
rect 52069 54539 60825 54595
rect 51034 54466 60825 54539
rect 36648 54452 40041 54453
rect 24298 54155 60825 54228
rect 24298 54099 29580 54155
rect 29636 54099 29791 54155
rect 29847 54099 30003 54155
rect 30059 54099 30214 54155
rect 30270 54099 30852 54155
rect 30908 54099 31063 54155
rect 31119 54099 31274 54155
rect 31330 54099 31484 54155
rect 31540 54099 31695 54155
rect 31751 54099 31907 54155
rect 31963 54099 32118 54155
rect 32174 54099 32328 54155
rect 32384 54099 32539 54155
rect 32595 54099 32750 54155
rect 32806 54099 35218 54155
rect 35274 54099 35428 54155
rect 35484 54099 35639 54155
rect 35695 54099 35851 54155
rect 35907 54099 36062 54155
rect 36118 54099 36272 54155
rect 36328 54099 39050 54155
rect 39106 54099 39230 54155
rect 39286 54099 44832 54155
rect 44888 54099 45043 54155
rect 45099 54099 45254 54155
rect 45310 54099 48836 54155
rect 48892 54099 49046 54155
rect 49102 54099 49257 54155
rect 49313 54099 49469 54155
rect 49525 54099 49680 54155
rect 49736 54099 49890 54155
rect 49946 54099 52314 54155
rect 52370 54099 52525 54155
rect 52581 54099 52736 54155
rect 52792 54099 52946 54155
rect 53002 54099 53157 54155
rect 53213 54099 53369 54155
rect 53425 54099 53580 54155
rect 53636 54099 53790 54155
rect 53846 54099 54001 54155
rect 54057 54099 54212 54155
rect 54268 54099 54853 54155
rect 54909 54099 55064 54155
rect 55120 54099 55276 54155
rect 55332 54099 55487 54155
rect 55543 54099 60825 54155
rect 24298 54027 60825 54099
rect 30403 54026 54622 54027
rect 36648 53801 40041 53802
rect 24298 53722 34090 53788
rect 24298 53666 33055 53722
rect 33111 53666 33235 53722
rect 33291 53715 34090 53722
rect 33291 53666 33817 53715
rect 24298 53659 33817 53666
rect 33873 53659 33997 53715
rect 34053 53659 34090 53715
rect 36640 53763 40085 53801
rect 36640 53707 36676 53763
rect 36732 53707 39992 53763
rect 40048 53707 40085 53763
rect 36640 53668 40085 53707
rect 48557 53749 48687 53788
rect 48557 53693 48594 53749
rect 48650 53693 48687 53749
rect 24298 53587 34090 53659
rect 30403 53586 34090 53587
rect 0 53376 1014 53576
rect 48557 53570 48687 53693
rect 51034 53715 60825 53788
rect 84666 53776 86372 54476
rect 51034 53659 51071 53715
rect 51127 53659 51251 53715
rect 51307 53659 51833 53715
rect 51889 53659 52013 53715
rect 52069 53659 60825 53715
rect 51034 53587 60825 53659
rect 51034 53586 54622 53587
rect 37852 53532 48687 53570
rect 37852 53476 37889 53532
rect 37945 53476 38069 53532
rect 38125 53476 39773 53532
rect 39829 53531 48687 53532
rect 39829 53476 48594 53531
rect 37852 53475 48594 53476
rect 48650 53475 48687 53531
rect 37852 53437 48687 53475
rect 85358 53376 86372 53576
rect 0 53328 27272 53376
rect 60471 53328 86372 53376
rect 0 53255 86372 53328
rect 0 53199 27788 53255
rect 27844 53199 27999 53255
rect 28055 53199 28210 53255
rect 28266 53199 28421 53255
rect 28477 53199 28632 53255
rect 28688 53199 28843 53255
rect 28899 53199 29054 53255
rect 29110 53199 34282 53255
rect 34338 53199 34493 53255
rect 34549 53199 34705 53255
rect 34761 53199 34916 53255
rect 34972 53199 38328 53255
rect 38384 53199 38539 53255
rect 38595 53199 38750 53255
rect 38806 53199 40251 53255
rect 40307 53199 40431 53255
rect 40487 53199 43788 53255
rect 43844 53199 43999 53255
rect 44055 53199 44211 53255
rect 44267 53199 44422 53255
rect 44478 53199 50161 53255
rect 50217 53199 50372 53255
rect 50428 53199 50584 53255
rect 50640 53199 50795 53255
rect 50851 53199 56013 53255
rect 56069 53199 56224 53255
rect 56280 53199 56435 53255
rect 56491 53199 56646 53255
rect 56702 53199 56857 53255
rect 56913 53199 57068 53255
rect 57124 53199 57279 53255
rect 57335 53199 86372 53255
rect 0 53127 86372 53199
rect 0 53076 27272 53127
rect 30403 53126 54622 53127
rect 60471 53076 86372 53127
rect 0 52876 1014 53076
rect 37852 52979 48687 53017
rect 37852 52978 48594 52979
rect 37852 52922 37889 52978
rect 37945 52922 38069 52978
rect 38125 52922 39773 52978
rect 39829 52923 48594 52978
rect 48650 52923 48687 52979
rect 39829 52922 48687 52923
rect 37852 52884 48687 52922
rect 24298 52795 34090 52868
rect 24298 52788 33817 52795
rect 24298 52732 33055 52788
rect 33111 52732 33235 52788
rect 33291 52739 33817 52788
rect 33873 52739 33997 52795
rect 34053 52739 34090 52795
rect 33291 52732 34090 52739
rect 0 51976 1706 52676
rect 24298 52666 34090 52732
rect 36640 52747 40085 52786
rect 36640 52691 36676 52747
rect 36732 52691 39992 52747
rect 40048 52691 40085 52747
rect 36640 52653 40085 52691
rect 48557 52761 48687 52884
rect 85358 52876 86372 53076
rect 48557 52705 48594 52761
rect 48650 52705 48687 52761
rect 48557 52666 48687 52705
rect 51034 52795 60825 52868
rect 51034 52739 51071 52795
rect 51127 52739 51251 52795
rect 51307 52739 51833 52795
rect 51889 52739 52013 52795
rect 52069 52739 60825 52795
rect 51034 52666 60825 52739
rect 36648 52652 40041 52653
rect 24298 52355 60825 52428
rect 24298 52299 29580 52355
rect 29636 52299 29791 52355
rect 29847 52299 30003 52355
rect 30059 52299 30214 52355
rect 30270 52299 30852 52355
rect 30908 52299 31063 52355
rect 31119 52299 31274 52355
rect 31330 52299 31484 52355
rect 31540 52299 31695 52355
rect 31751 52299 31907 52355
rect 31963 52299 32118 52355
rect 32174 52299 32328 52355
rect 32384 52299 32539 52355
rect 32595 52299 32750 52355
rect 32806 52299 35218 52355
rect 35274 52299 35428 52355
rect 35484 52299 35639 52355
rect 35695 52299 35851 52355
rect 35907 52299 36062 52355
rect 36118 52299 36272 52355
rect 36328 52299 39050 52355
rect 39106 52299 39230 52355
rect 39286 52299 44832 52355
rect 44888 52299 45043 52355
rect 45099 52299 45254 52355
rect 45310 52299 48836 52355
rect 48892 52299 49046 52355
rect 49102 52299 49257 52355
rect 49313 52299 49469 52355
rect 49525 52299 49680 52355
rect 49736 52299 49890 52355
rect 49946 52299 52314 52355
rect 52370 52299 52525 52355
rect 52581 52299 52736 52355
rect 52792 52299 52946 52355
rect 53002 52299 53157 52355
rect 53213 52299 53369 52355
rect 53425 52299 53580 52355
rect 53636 52299 53790 52355
rect 53846 52299 54001 52355
rect 54057 52299 54212 52355
rect 54268 52299 54853 52355
rect 54909 52299 55064 52355
rect 55120 52299 55276 52355
rect 55332 52299 55487 52355
rect 55543 52299 60825 52355
rect 24298 52227 60825 52299
rect 30403 52226 54622 52227
rect 36648 52001 40041 52002
rect 24298 51922 34090 51988
rect 24298 51866 33055 51922
rect 33111 51866 33235 51922
rect 33291 51915 34090 51922
rect 33291 51866 33817 51915
rect 24298 51859 33817 51866
rect 33873 51859 33997 51915
rect 34053 51859 34090 51915
rect 36640 51963 40085 52001
rect 36640 51907 36676 51963
rect 36732 51907 39992 51963
rect 40048 51907 40085 51963
rect 36640 51868 40085 51907
rect 48557 51949 48687 51988
rect 48557 51893 48594 51949
rect 48650 51893 48687 51949
rect 24298 51787 34090 51859
rect 30403 51786 34090 51787
rect 0 51576 1014 51776
rect 48557 51770 48687 51893
rect 51034 51915 60825 51988
rect 84666 51976 86372 52676
rect 51034 51859 51071 51915
rect 51127 51859 51251 51915
rect 51307 51859 51833 51915
rect 51889 51859 52013 51915
rect 52069 51859 60825 51915
rect 51034 51787 60825 51859
rect 51034 51786 54622 51787
rect 37852 51732 48687 51770
rect 37852 51676 37889 51732
rect 37945 51676 38069 51732
rect 38125 51676 39773 51732
rect 39829 51731 48687 51732
rect 39829 51676 48594 51731
rect 37852 51675 48594 51676
rect 48650 51675 48687 51731
rect 37852 51637 48687 51675
rect 85358 51576 86372 51776
rect 0 51528 27272 51576
rect 60471 51528 86372 51576
rect 0 51455 86372 51528
rect 0 51399 27788 51455
rect 27844 51399 27999 51455
rect 28055 51399 28210 51455
rect 28266 51399 28421 51455
rect 28477 51399 28632 51455
rect 28688 51399 28843 51455
rect 28899 51399 29054 51455
rect 29110 51399 34282 51455
rect 34338 51399 34493 51455
rect 34549 51399 34705 51455
rect 34761 51399 34916 51455
rect 34972 51399 38328 51455
rect 38384 51399 38539 51455
rect 38595 51399 38750 51455
rect 38806 51399 40251 51455
rect 40307 51399 40431 51455
rect 40487 51399 43788 51455
rect 43844 51399 43999 51455
rect 44055 51399 44211 51455
rect 44267 51399 44422 51455
rect 44478 51399 50161 51455
rect 50217 51399 50372 51455
rect 50428 51399 50584 51455
rect 50640 51399 50795 51455
rect 50851 51399 56013 51455
rect 56069 51399 56224 51455
rect 56280 51399 56435 51455
rect 56491 51399 56646 51455
rect 56702 51399 56857 51455
rect 56913 51399 57068 51455
rect 57124 51399 57279 51455
rect 57335 51399 86372 51455
rect 0 51327 86372 51399
rect 0 51276 27272 51327
rect 30403 51326 54622 51327
rect 60471 51276 86372 51327
rect 0 51076 1014 51276
rect 37852 51179 48687 51217
rect 37852 51178 48594 51179
rect 37852 51122 37889 51178
rect 37945 51122 38069 51178
rect 38125 51122 39773 51178
rect 39829 51123 48594 51178
rect 48650 51123 48687 51179
rect 39829 51122 48687 51123
rect 37852 51084 48687 51122
rect 24298 50995 34090 51068
rect 24298 50988 33817 50995
rect 24298 50932 33055 50988
rect 33111 50932 33235 50988
rect 33291 50939 33817 50988
rect 33873 50939 33997 50995
rect 34053 50939 34090 50995
rect 33291 50932 34090 50939
rect 0 50176 1706 50876
rect 24298 50866 34090 50932
rect 36640 50947 40085 50986
rect 36640 50891 36676 50947
rect 36732 50891 39992 50947
rect 40048 50891 40085 50947
rect 36640 50853 40085 50891
rect 48557 50961 48687 51084
rect 85358 51076 86372 51276
rect 48557 50905 48594 50961
rect 48650 50905 48687 50961
rect 48557 50866 48687 50905
rect 51034 50995 60825 51068
rect 51034 50939 51071 50995
rect 51127 50939 51251 50995
rect 51307 50939 51833 50995
rect 51889 50939 52013 50995
rect 52069 50939 60825 50995
rect 51034 50866 60825 50939
rect 36648 50852 40041 50853
rect 24298 50555 60825 50628
rect 24298 50499 29580 50555
rect 29636 50499 29791 50555
rect 29847 50499 30003 50555
rect 30059 50499 30214 50555
rect 30270 50499 30852 50555
rect 30908 50499 31063 50555
rect 31119 50499 31274 50555
rect 31330 50499 31484 50555
rect 31540 50499 31695 50555
rect 31751 50499 31907 50555
rect 31963 50499 32118 50555
rect 32174 50499 32328 50555
rect 32384 50499 32539 50555
rect 32595 50499 32750 50555
rect 32806 50499 35218 50555
rect 35274 50499 35428 50555
rect 35484 50499 35639 50555
rect 35695 50499 35851 50555
rect 35907 50499 36062 50555
rect 36118 50499 36272 50555
rect 36328 50499 39050 50555
rect 39106 50499 39230 50555
rect 39286 50499 44832 50555
rect 44888 50499 45043 50555
rect 45099 50499 45254 50555
rect 45310 50499 48836 50555
rect 48892 50499 49046 50555
rect 49102 50499 49257 50555
rect 49313 50499 49469 50555
rect 49525 50499 49680 50555
rect 49736 50499 49890 50555
rect 49946 50499 52314 50555
rect 52370 50499 52525 50555
rect 52581 50499 52736 50555
rect 52792 50499 52946 50555
rect 53002 50499 53157 50555
rect 53213 50499 53369 50555
rect 53425 50499 53580 50555
rect 53636 50499 53790 50555
rect 53846 50499 54001 50555
rect 54057 50499 54212 50555
rect 54268 50499 54853 50555
rect 54909 50499 55064 50555
rect 55120 50499 55276 50555
rect 55332 50499 55487 50555
rect 55543 50499 60825 50555
rect 24298 50427 60825 50499
rect 30403 50426 54622 50427
rect 36648 50201 40041 50202
rect 24298 50122 34090 50188
rect 24298 50066 33055 50122
rect 33111 50066 33235 50122
rect 33291 50115 34090 50122
rect 33291 50066 33817 50115
rect 24298 50059 33817 50066
rect 33873 50059 33997 50115
rect 34053 50059 34090 50115
rect 36640 50163 40085 50201
rect 36640 50107 36676 50163
rect 36732 50107 39992 50163
rect 40048 50107 40085 50163
rect 36640 50068 40085 50107
rect 48557 50149 48687 50188
rect 48557 50093 48594 50149
rect 48650 50093 48687 50149
rect 24298 49987 34090 50059
rect 30403 49986 34090 49987
rect 0 49776 1014 49976
rect 48557 49970 48687 50093
rect 51034 50115 60825 50188
rect 84666 50176 86372 50876
rect 51034 50059 51071 50115
rect 51127 50059 51251 50115
rect 51307 50059 51833 50115
rect 51889 50059 52013 50115
rect 52069 50059 60825 50115
rect 51034 49987 60825 50059
rect 51034 49986 54622 49987
rect 37852 49932 48687 49970
rect 37852 49876 37889 49932
rect 37945 49876 38069 49932
rect 38125 49876 39773 49932
rect 39829 49931 48687 49932
rect 39829 49876 48594 49931
rect 37852 49875 48594 49876
rect 48650 49875 48687 49931
rect 37852 49837 48687 49875
rect 85358 49776 86372 49976
rect 0 49728 27272 49776
rect 60471 49728 86372 49776
rect 0 49655 86372 49728
rect 0 49599 27788 49655
rect 27844 49599 27999 49655
rect 28055 49599 28210 49655
rect 28266 49599 28421 49655
rect 28477 49599 28632 49655
rect 28688 49599 28843 49655
rect 28899 49599 29054 49655
rect 29110 49599 34282 49655
rect 34338 49599 34493 49655
rect 34549 49599 34705 49655
rect 34761 49599 34916 49655
rect 34972 49599 38328 49655
rect 38384 49599 38539 49655
rect 38595 49599 38750 49655
rect 38806 49599 40251 49655
rect 40307 49599 40431 49655
rect 40487 49599 43788 49655
rect 43844 49599 43999 49655
rect 44055 49599 44211 49655
rect 44267 49599 44422 49655
rect 44478 49599 50161 49655
rect 50217 49599 50372 49655
rect 50428 49599 50584 49655
rect 50640 49599 50795 49655
rect 50851 49599 56013 49655
rect 56069 49599 56224 49655
rect 56280 49599 56435 49655
rect 56491 49599 56646 49655
rect 56702 49599 56857 49655
rect 56913 49599 57068 49655
rect 57124 49599 57279 49655
rect 57335 49599 86372 49655
rect 0 49527 86372 49599
rect 0 49476 27272 49527
rect 30403 49526 54622 49527
rect 60471 49476 86372 49527
rect 0 49276 1014 49476
rect 37852 49379 48687 49417
rect 37852 49378 48594 49379
rect 37852 49322 37889 49378
rect 37945 49322 38069 49378
rect 38125 49322 39773 49378
rect 39829 49323 48594 49378
rect 48650 49323 48687 49379
rect 39829 49322 48687 49323
rect 37852 49284 48687 49322
rect 24298 49195 34090 49268
rect 24298 49188 33817 49195
rect 24298 49132 33055 49188
rect 33111 49132 33235 49188
rect 33291 49139 33817 49188
rect 33873 49139 33997 49195
rect 34053 49139 34090 49195
rect 33291 49132 34090 49139
rect 0 48376 1706 49076
rect 24298 49066 34090 49132
rect 36640 49147 40085 49186
rect 36640 49091 36676 49147
rect 36732 49091 39992 49147
rect 40048 49091 40085 49147
rect 36640 49053 40085 49091
rect 48557 49161 48687 49284
rect 85358 49276 86372 49476
rect 48557 49105 48594 49161
rect 48650 49105 48687 49161
rect 48557 49066 48687 49105
rect 51034 49195 60825 49268
rect 51034 49139 51071 49195
rect 51127 49139 51251 49195
rect 51307 49139 51833 49195
rect 51889 49139 52013 49195
rect 52069 49139 60825 49195
rect 51034 49066 60825 49139
rect 36648 49052 40041 49053
rect 24298 48755 60825 48828
rect 24298 48699 29580 48755
rect 29636 48699 29791 48755
rect 29847 48699 30003 48755
rect 30059 48699 30214 48755
rect 30270 48699 30852 48755
rect 30908 48699 31063 48755
rect 31119 48699 31274 48755
rect 31330 48699 31484 48755
rect 31540 48699 31695 48755
rect 31751 48699 31907 48755
rect 31963 48699 32118 48755
rect 32174 48699 32328 48755
rect 32384 48699 32539 48755
rect 32595 48699 32750 48755
rect 32806 48699 35218 48755
rect 35274 48699 35428 48755
rect 35484 48699 35639 48755
rect 35695 48699 35851 48755
rect 35907 48699 36062 48755
rect 36118 48699 36272 48755
rect 36328 48699 39050 48755
rect 39106 48699 39230 48755
rect 39286 48699 44832 48755
rect 44888 48699 45043 48755
rect 45099 48699 45254 48755
rect 45310 48699 48836 48755
rect 48892 48699 49046 48755
rect 49102 48699 49257 48755
rect 49313 48699 49469 48755
rect 49525 48699 49680 48755
rect 49736 48699 49890 48755
rect 49946 48699 52314 48755
rect 52370 48699 52525 48755
rect 52581 48699 52736 48755
rect 52792 48699 52946 48755
rect 53002 48699 53157 48755
rect 53213 48699 53369 48755
rect 53425 48699 53580 48755
rect 53636 48699 53790 48755
rect 53846 48699 54001 48755
rect 54057 48699 54212 48755
rect 54268 48699 54853 48755
rect 54909 48699 55064 48755
rect 55120 48699 55276 48755
rect 55332 48699 55487 48755
rect 55543 48699 60825 48755
rect 24298 48627 60825 48699
rect 30403 48626 54622 48627
rect 36648 48401 40041 48402
rect 24298 48322 34090 48388
rect 24298 48266 33055 48322
rect 33111 48266 33235 48322
rect 33291 48315 34090 48322
rect 33291 48266 33817 48315
rect 24298 48259 33817 48266
rect 33873 48259 33997 48315
rect 34053 48259 34090 48315
rect 36640 48363 40085 48401
rect 36640 48307 36676 48363
rect 36732 48307 39992 48363
rect 40048 48307 40085 48363
rect 36640 48268 40085 48307
rect 48557 48349 48687 48388
rect 48557 48293 48594 48349
rect 48650 48293 48687 48349
rect 24298 48187 34090 48259
rect 30403 48186 34090 48187
rect 0 47976 1014 48176
rect 48557 48170 48687 48293
rect 51034 48315 60825 48388
rect 84666 48376 86372 49076
rect 51034 48259 51071 48315
rect 51127 48259 51251 48315
rect 51307 48259 51833 48315
rect 51889 48259 52013 48315
rect 52069 48259 60825 48315
rect 51034 48187 60825 48259
rect 51034 48186 54622 48187
rect 37852 48132 48687 48170
rect 37852 48076 37889 48132
rect 37945 48076 38069 48132
rect 38125 48076 39773 48132
rect 39829 48131 48687 48132
rect 39829 48076 48594 48131
rect 37852 48075 48594 48076
rect 48650 48075 48687 48131
rect 37852 48037 48687 48075
rect 85358 47976 86372 48176
rect 0 47928 27272 47976
rect 60471 47928 86372 47976
rect 0 47855 86372 47928
rect 0 47799 27788 47855
rect 27844 47799 27999 47855
rect 28055 47799 28210 47855
rect 28266 47799 28421 47855
rect 28477 47799 28632 47855
rect 28688 47799 28843 47855
rect 28899 47799 29054 47855
rect 29110 47799 34282 47855
rect 34338 47799 34493 47855
rect 34549 47799 34705 47855
rect 34761 47799 34916 47855
rect 34972 47799 38328 47855
rect 38384 47799 38539 47855
rect 38595 47799 38750 47855
rect 38806 47799 40251 47855
rect 40307 47799 40431 47855
rect 40487 47799 43788 47855
rect 43844 47799 43999 47855
rect 44055 47799 44211 47855
rect 44267 47799 44422 47855
rect 44478 47799 50161 47855
rect 50217 47799 50372 47855
rect 50428 47799 50584 47855
rect 50640 47799 50795 47855
rect 50851 47799 56013 47855
rect 56069 47799 56224 47855
rect 56280 47799 56435 47855
rect 56491 47799 56646 47855
rect 56702 47799 56857 47855
rect 56913 47799 57068 47855
rect 57124 47799 57279 47855
rect 57335 47799 86372 47855
rect 0 47727 86372 47799
rect 0 47676 27272 47727
rect 30403 47726 54622 47727
rect 60471 47676 86372 47727
rect 0 47476 1014 47676
rect 37852 47579 48687 47617
rect 37852 47578 48594 47579
rect 37852 47522 37889 47578
rect 37945 47522 38069 47578
rect 38125 47522 39773 47578
rect 39829 47523 48594 47578
rect 48650 47523 48687 47579
rect 39829 47522 48687 47523
rect 37852 47484 48687 47522
rect 24298 47395 34090 47468
rect 24298 47388 33817 47395
rect 24298 47332 33055 47388
rect 33111 47332 33235 47388
rect 33291 47339 33817 47388
rect 33873 47339 33997 47395
rect 34053 47339 34090 47395
rect 33291 47332 34090 47339
rect 0 46576 1706 47276
rect 24298 47266 34090 47332
rect 36640 47347 40085 47386
rect 36640 47291 36676 47347
rect 36732 47291 39992 47347
rect 40048 47291 40085 47347
rect 36640 47253 40085 47291
rect 48557 47361 48687 47484
rect 85358 47476 86372 47676
rect 48557 47305 48594 47361
rect 48650 47305 48687 47361
rect 48557 47266 48687 47305
rect 51034 47395 60825 47468
rect 51034 47339 51071 47395
rect 51127 47339 51251 47395
rect 51307 47339 51833 47395
rect 51889 47339 52013 47395
rect 52069 47339 60825 47395
rect 51034 47266 60825 47339
rect 36648 47252 40041 47253
rect 24298 46955 60825 47028
rect 24298 46899 29580 46955
rect 29636 46899 29791 46955
rect 29847 46899 30003 46955
rect 30059 46899 30214 46955
rect 30270 46899 30852 46955
rect 30908 46899 31063 46955
rect 31119 46899 31274 46955
rect 31330 46899 31484 46955
rect 31540 46899 31695 46955
rect 31751 46899 31907 46955
rect 31963 46899 32118 46955
rect 32174 46899 32328 46955
rect 32384 46899 32539 46955
rect 32595 46899 32750 46955
rect 32806 46899 35218 46955
rect 35274 46899 35428 46955
rect 35484 46899 35639 46955
rect 35695 46899 35851 46955
rect 35907 46899 36062 46955
rect 36118 46899 36272 46955
rect 36328 46899 39050 46955
rect 39106 46899 39230 46955
rect 39286 46899 44832 46955
rect 44888 46899 45043 46955
rect 45099 46899 45254 46955
rect 45310 46899 48836 46955
rect 48892 46899 49046 46955
rect 49102 46899 49257 46955
rect 49313 46899 49469 46955
rect 49525 46899 49680 46955
rect 49736 46899 49890 46955
rect 49946 46899 52314 46955
rect 52370 46899 52525 46955
rect 52581 46899 52736 46955
rect 52792 46899 52946 46955
rect 53002 46899 53157 46955
rect 53213 46899 53369 46955
rect 53425 46899 53580 46955
rect 53636 46899 53790 46955
rect 53846 46899 54001 46955
rect 54057 46899 54212 46955
rect 54268 46899 54853 46955
rect 54909 46899 55064 46955
rect 55120 46899 55276 46955
rect 55332 46899 55487 46955
rect 55543 46899 60825 46955
rect 24298 46827 60825 46899
rect 30403 46826 54622 46827
rect 36648 46601 40041 46602
rect 24298 46522 34090 46588
rect 24298 46466 33055 46522
rect 33111 46466 33235 46522
rect 33291 46515 34090 46522
rect 33291 46466 33817 46515
rect 24298 46459 33817 46466
rect 33873 46459 33997 46515
rect 34053 46459 34090 46515
rect 36640 46563 40085 46601
rect 36640 46507 36676 46563
rect 36732 46507 39992 46563
rect 40048 46507 40085 46563
rect 36640 46468 40085 46507
rect 48557 46549 48687 46588
rect 48557 46493 48594 46549
rect 48650 46493 48687 46549
rect 24298 46387 34090 46459
rect 30403 46386 34090 46387
rect 0 46176 1014 46376
rect 48557 46370 48687 46493
rect 51034 46515 60825 46588
rect 84666 46576 86372 47276
rect 51034 46459 51071 46515
rect 51127 46459 51251 46515
rect 51307 46459 51833 46515
rect 51889 46459 52013 46515
rect 52069 46459 60825 46515
rect 51034 46387 60825 46459
rect 51034 46386 54622 46387
rect 37852 46332 48687 46370
rect 37852 46276 37889 46332
rect 37945 46276 38069 46332
rect 38125 46276 39773 46332
rect 39829 46331 48687 46332
rect 39829 46276 48594 46331
rect 37852 46275 48594 46276
rect 48650 46275 48687 46331
rect 37852 46237 48687 46275
rect 85358 46176 86372 46376
rect 0 46128 27272 46176
rect 60471 46128 86372 46176
rect 0 46055 86372 46128
rect 0 45999 27788 46055
rect 27844 45999 27999 46055
rect 28055 45999 28210 46055
rect 28266 45999 28421 46055
rect 28477 45999 28632 46055
rect 28688 45999 28843 46055
rect 28899 45999 29054 46055
rect 29110 45999 34282 46055
rect 34338 45999 34493 46055
rect 34549 45999 34705 46055
rect 34761 45999 34916 46055
rect 34972 45999 38328 46055
rect 38384 45999 38539 46055
rect 38595 45999 38750 46055
rect 38806 45999 40251 46055
rect 40307 45999 40431 46055
rect 40487 45999 43788 46055
rect 43844 45999 43999 46055
rect 44055 45999 44211 46055
rect 44267 45999 44422 46055
rect 44478 45999 50161 46055
rect 50217 45999 50372 46055
rect 50428 45999 50584 46055
rect 50640 45999 50795 46055
rect 50851 45999 56013 46055
rect 56069 45999 56224 46055
rect 56280 45999 56435 46055
rect 56491 45999 56646 46055
rect 56702 45999 56857 46055
rect 56913 45999 57068 46055
rect 57124 45999 57279 46055
rect 57335 45999 86372 46055
rect 0 45927 86372 45999
rect 0 45876 27272 45927
rect 30403 45926 54622 45927
rect 60471 45876 86372 45927
rect 0 45676 1014 45876
rect 37852 45779 48687 45817
rect 37852 45778 48594 45779
rect 37852 45722 37889 45778
rect 37945 45722 38069 45778
rect 38125 45722 39773 45778
rect 39829 45723 48594 45778
rect 48650 45723 48687 45779
rect 39829 45722 48687 45723
rect 37852 45684 48687 45722
rect 24298 45595 34090 45668
rect 24298 45588 33817 45595
rect 24298 45532 33055 45588
rect 33111 45532 33235 45588
rect 33291 45539 33817 45588
rect 33873 45539 33997 45595
rect 34053 45539 34090 45595
rect 33291 45532 34090 45539
rect 0 44776 1706 45476
rect 24298 45466 34090 45532
rect 36640 45547 40085 45586
rect 36640 45491 36676 45547
rect 36732 45491 39992 45547
rect 40048 45491 40085 45547
rect 36640 45453 40085 45491
rect 48557 45561 48687 45684
rect 85358 45676 86372 45876
rect 48557 45505 48594 45561
rect 48650 45505 48687 45561
rect 48557 45466 48687 45505
rect 51034 45595 60825 45668
rect 51034 45539 51071 45595
rect 51127 45539 51251 45595
rect 51307 45539 51833 45595
rect 51889 45539 52013 45595
rect 52069 45539 60825 45595
rect 51034 45466 60825 45539
rect 36648 45452 40041 45453
rect 24298 45155 60825 45228
rect 24298 45099 29580 45155
rect 29636 45099 29791 45155
rect 29847 45099 30003 45155
rect 30059 45099 30214 45155
rect 30270 45099 30852 45155
rect 30908 45099 31063 45155
rect 31119 45099 31274 45155
rect 31330 45099 31484 45155
rect 31540 45099 31695 45155
rect 31751 45099 31907 45155
rect 31963 45099 32118 45155
rect 32174 45099 32328 45155
rect 32384 45099 32539 45155
rect 32595 45099 32750 45155
rect 32806 45099 35218 45155
rect 35274 45099 35428 45155
rect 35484 45099 35639 45155
rect 35695 45099 35851 45155
rect 35907 45099 36062 45155
rect 36118 45099 36272 45155
rect 36328 45099 39050 45155
rect 39106 45099 39230 45155
rect 39286 45099 44832 45155
rect 44888 45099 45043 45155
rect 45099 45099 45254 45155
rect 45310 45099 48836 45155
rect 48892 45099 49046 45155
rect 49102 45099 49257 45155
rect 49313 45099 49469 45155
rect 49525 45099 49680 45155
rect 49736 45099 49890 45155
rect 49946 45099 52314 45155
rect 52370 45099 52525 45155
rect 52581 45099 52736 45155
rect 52792 45099 52946 45155
rect 53002 45099 53157 45155
rect 53213 45099 53369 45155
rect 53425 45099 53580 45155
rect 53636 45099 53790 45155
rect 53846 45099 54001 45155
rect 54057 45099 54212 45155
rect 54268 45099 54853 45155
rect 54909 45099 55064 45155
rect 55120 45099 55276 45155
rect 55332 45099 55487 45155
rect 55543 45099 60825 45155
rect 24298 45027 60825 45099
rect 30403 45026 54622 45027
rect 36648 44801 40041 44802
rect 24298 44722 34090 44788
rect 24298 44666 33055 44722
rect 33111 44666 33235 44722
rect 33291 44715 34090 44722
rect 33291 44666 33817 44715
rect 24298 44659 33817 44666
rect 33873 44659 33997 44715
rect 34053 44659 34090 44715
rect 36640 44763 40085 44801
rect 36640 44707 36676 44763
rect 36732 44707 39992 44763
rect 40048 44707 40085 44763
rect 36640 44668 40085 44707
rect 48557 44749 48687 44788
rect 48557 44693 48594 44749
rect 48650 44693 48687 44749
rect 24298 44587 34090 44659
rect 30403 44586 34090 44587
rect 0 44376 1014 44576
rect 48557 44570 48687 44693
rect 51034 44715 60825 44788
rect 84666 44776 86372 45476
rect 51034 44659 51071 44715
rect 51127 44659 51251 44715
rect 51307 44659 51833 44715
rect 51889 44659 52013 44715
rect 52069 44659 60825 44715
rect 51034 44587 60825 44659
rect 51034 44586 54622 44587
rect 37852 44532 48687 44570
rect 37852 44476 37889 44532
rect 37945 44476 38069 44532
rect 38125 44476 39773 44532
rect 39829 44531 48687 44532
rect 39829 44476 48594 44531
rect 37852 44475 48594 44476
rect 48650 44475 48687 44531
rect 37852 44437 48687 44475
rect 85358 44376 86372 44576
rect 0 44328 27272 44376
rect 60471 44328 86372 44376
rect 0 44255 86372 44328
rect 0 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 34282 44255
rect 34338 44199 34493 44255
rect 34549 44199 34705 44255
rect 34761 44199 34916 44255
rect 34972 44199 38328 44255
rect 38384 44199 38539 44255
rect 38595 44199 38750 44255
rect 38806 44199 40251 44255
rect 40307 44199 40431 44255
rect 40487 44199 43788 44255
rect 43844 44199 43999 44255
rect 44055 44199 44211 44255
rect 44267 44199 44422 44255
rect 44478 44199 50161 44255
rect 50217 44199 50372 44255
rect 50428 44199 50584 44255
rect 50640 44199 50795 44255
rect 50851 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 86372 44255
rect 0 44127 86372 44199
rect 0 44076 27272 44127
rect 30403 44126 54622 44127
rect 60471 44076 86372 44127
rect 0 43876 1014 44076
rect 37852 43979 48687 44017
rect 37852 43978 48594 43979
rect 37852 43922 37889 43978
rect 37945 43922 38069 43978
rect 38125 43922 39773 43978
rect 39829 43923 48594 43978
rect 48650 43923 48687 43979
rect 39829 43922 48687 43923
rect 37852 43884 48687 43922
rect 24298 43795 34090 43868
rect 24298 43788 33817 43795
rect 24298 43732 33055 43788
rect 33111 43732 33235 43788
rect 33291 43739 33817 43788
rect 33873 43739 33997 43795
rect 34053 43739 34090 43795
rect 33291 43732 34090 43739
rect 0 42976 1706 43676
rect 24298 43666 34090 43732
rect 36640 43747 40085 43786
rect 36640 43691 36676 43747
rect 36732 43691 39992 43747
rect 40048 43691 40085 43747
rect 36640 43653 40085 43691
rect 48557 43761 48687 43884
rect 85358 43876 86372 44076
rect 48557 43705 48594 43761
rect 48650 43705 48687 43761
rect 48557 43666 48687 43705
rect 51034 43795 60825 43868
rect 51034 43739 51071 43795
rect 51127 43739 51251 43795
rect 51307 43739 51833 43795
rect 51889 43739 52013 43795
rect 52069 43739 60825 43795
rect 51034 43666 60825 43739
rect 36648 43652 40041 43653
rect 24298 43355 60825 43428
rect 24298 43299 29580 43355
rect 29636 43299 29791 43355
rect 29847 43299 30003 43355
rect 30059 43299 30214 43355
rect 30270 43299 30852 43355
rect 30908 43299 31063 43355
rect 31119 43299 31274 43355
rect 31330 43299 31484 43355
rect 31540 43299 31695 43355
rect 31751 43299 31907 43355
rect 31963 43299 32118 43355
rect 32174 43299 32328 43355
rect 32384 43299 32539 43355
rect 32595 43299 32750 43355
rect 32806 43299 35218 43355
rect 35274 43299 35428 43355
rect 35484 43299 35639 43355
rect 35695 43299 35851 43355
rect 35907 43299 36062 43355
rect 36118 43299 36272 43355
rect 36328 43299 39050 43355
rect 39106 43299 39230 43355
rect 39286 43299 44832 43355
rect 44888 43299 45043 43355
rect 45099 43299 45254 43355
rect 45310 43299 48836 43355
rect 48892 43299 49046 43355
rect 49102 43299 49257 43355
rect 49313 43299 49469 43355
rect 49525 43299 49680 43355
rect 49736 43299 49890 43355
rect 49946 43299 52314 43355
rect 52370 43299 52525 43355
rect 52581 43299 52736 43355
rect 52792 43299 52946 43355
rect 53002 43299 53157 43355
rect 53213 43299 53369 43355
rect 53425 43299 53580 43355
rect 53636 43299 53790 43355
rect 53846 43299 54001 43355
rect 54057 43299 54212 43355
rect 54268 43299 54853 43355
rect 54909 43299 55064 43355
rect 55120 43299 55276 43355
rect 55332 43299 55487 43355
rect 55543 43299 60825 43355
rect 24298 43227 60825 43299
rect 30403 43226 54622 43227
rect 36648 43001 40041 43002
rect 24298 42922 34090 42988
rect 24298 42866 33055 42922
rect 33111 42866 33235 42922
rect 33291 42915 34090 42922
rect 33291 42866 33817 42915
rect 24298 42859 33817 42866
rect 33873 42859 33997 42915
rect 34053 42859 34090 42915
rect 36640 42963 40085 43001
rect 36640 42907 36676 42963
rect 36732 42907 39992 42963
rect 40048 42907 40085 42963
rect 36640 42868 40085 42907
rect 48557 42949 48687 42988
rect 48557 42893 48594 42949
rect 48650 42893 48687 42949
rect 24298 42787 34090 42859
rect 30403 42786 34090 42787
rect 0 42576 1014 42776
rect 48557 42770 48687 42893
rect 51034 42915 60825 42988
rect 84666 42976 86372 43676
rect 51034 42859 51071 42915
rect 51127 42859 51251 42915
rect 51307 42859 51833 42915
rect 51889 42859 52013 42915
rect 52069 42859 60825 42915
rect 51034 42787 60825 42859
rect 51034 42786 54622 42787
rect 37852 42732 48687 42770
rect 37852 42676 37889 42732
rect 37945 42676 38069 42732
rect 38125 42676 39773 42732
rect 39829 42731 48687 42732
rect 39829 42676 48594 42731
rect 37852 42675 48594 42676
rect 48650 42675 48687 42731
rect 37852 42637 48687 42675
rect 85358 42576 86372 42776
rect 0 42528 27272 42576
rect 60471 42528 86372 42576
rect 0 42455 86372 42528
rect 0 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 34282 42455
rect 34338 42399 34493 42455
rect 34549 42399 34705 42455
rect 34761 42399 34916 42455
rect 34972 42399 38328 42455
rect 38384 42399 38539 42455
rect 38595 42399 38750 42455
rect 38806 42399 40251 42455
rect 40307 42399 40431 42455
rect 40487 42399 43788 42455
rect 43844 42399 43999 42455
rect 44055 42399 44211 42455
rect 44267 42399 44422 42455
rect 44478 42399 50161 42455
rect 50217 42399 50372 42455
rect 50428 42399 50584 42455
rect 50640 42399 50795 42455
rect 50851 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 86372 42455
rect 0 42327 86372 42399
rect 0 42276 27272 42327
rect 30403 42326 54622 42327
rect 60471 42276 86372 42327
rect 0 42076 1014 42276
rect 37852 42179 48687 42217
rect 37852 42178 48594 42179
rect 37852 42122 37889 42178
rect 37945 42122 38069 42178
rect 38125 42122 39773 42178
rect 39829 42123 48594 42178
rect 48650 42123 48687 42179
rect 39829 42122 48687 42123
rect 37852 42084 48687 42122
rect 24298 41995 34090 42068
rect 24298 41988 33817 41995
rect 24298 41932 33055 41988
rect 33111 41932 33235 41988
rect 33291 41939 33817 41988
rect 33873 41939 33997 41995
rect 34053 41939 34090 41995
rect 33291 41932 34090 41939
rect 0 41176 1706 41876
rect 24298 41866 34090 41932
rect 36640 41947 40085 41986
rect 36640 41891 36676 41947
rect 36732 41891 39992 41947
rect 40048 41891 40085 41947
rect 36640 41853 40085 41891
rect 48557 41961 48687 42084
rect 85358 42076 86372 42276
rect 48557 41905 48594 41961
rect 48650 41905 48687 41961
rect 48557 41866 48687 41905
rect 51034 41995 60825 42068
rect 51034 41939 51071 41995
rect 51127 41939 51251 41995
rect 51307 41939 51833 41995
rect 51889 41939 52013 41995
rect 52069 41939 60825 41995
rect 51034 41866 60825 41939
rect 36648 41852 40041 41853
rect 24298 41555 60825 41628
rect 24298 41499 29580 41555
rect 29636 41499 29791 41555
rect 29847 41499 30003 41555
rect 30059 41499 30214 41555
rect 30270 41499 30852 41555
rect 30908 41499 31063 41555
rect 31119 41499 31274 41555
rect 31330 41499 31484 41555
rect 31540 41499 31695 41555
rect 31751 41499 31907 41555
rect 31963 41499 32118 41555
rect 32174 41499 32328 41555
rect 32384 41499 32539 41555
rect 32595 41499 32750 41555
rect 32806 41499 35218 41555
rect 35274 41499 35428 41555
rect 35484 41499 35639 41555
rect 35695 41499 35851 41555
rect 35907 41499 36062 41555
rect 36118 41499 36272 41555
rect 36328 41499 39050 41555
rect 39106 41499 39230 41555
rect 39286 41499 44832 41555
rect 44888 41499 45043 41555
rect 45099 41499 45254 41555
rect 45310 41499 48836 41555
rect 48892 41499 49046 41555
rect 49102 41499 49257 41555
rect 49313 41499 49469 41555
rect 49525 41499 49680 41555
rect 49736 41499 49890 41555
rect 49946 41499 52314 41555
rect 52370 41499 52525 41555
rect 52581 41499 52736 41555
rect 52792 41499 52946 41555
rect 53002 41499 53157 41555
rect 53213 41499 53369 41555
rect 53425 41499 53580 41555
rect 53636 41499 53790 41555
rect 53846 41499 54001 41555
rect 54057 41499 54212 41555
rect 54268 41499 54853 41555
rect 54909 41499 55064 41555
rect 55120 41499 55276 41555
rect 55332 41499 55487 41555
rect 55543 41499 60825 41555
rect 24298 41427 60825 41499
rect 30403 41426 54622 41427
rect 36648 41201 40041 41202
rect 24298 41122 34090 41188
rect 24298 41066 33055 41122
rect 33111 41066 33235 41122
rect 33291 41115 34090 41122
rect 33291 41066 33817 41115
rect 24298 41059 33817 41066
rect 33873 41059 33997 41115
rect 34053 41059 34090 41115
rect 36640 41163 40085 41201
rect 36640 41107 36676 41163
rect 36732 41107 39992 41163
rect 40048 41107 40085 41163
rect 36640 41068 40085 41107
rect 48557 41149 48687 41188
rect 48557 41093 48594 41149
rect 48650 41093 48687 41149
rect 24298 40987 34090 41059
rect 30403 40986 34090 40987
rect 0 40776 1014 40976
rect 48557 40970 48687 41093
rect 51034 41115 60825 41188
rect 84666 41176 86372 41876
rect 51034 41059 51071 41115
rect 51127 41059 51251 41115
rect 51307 41059 51833 41115
rect 51889 41059 52013 41115
rect 52069 41059 60825 41115
rect 51034 40987 60825 41059
rect 51034 40986 54622 40987
rect 37852 40932 48687 40970
rect 37852 40876 37889 40932
rect 37945 40876 38069 40932
rect 38125 40876 39773 40932
rect 39829 40931 48687 40932
rect 39829 40876 48594 40931
rect 37852 40875 48594 40876
rect 48650 40875 48687 40931
rect 37852 40837 48687 40875
rect 85358 40776 86372 40976
rect 0 40728 27272 40776
rect 60471 40728 86372 40776
rect 0 40655 86372 40728
rect 0 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 34282 40655
rect 34338 40599 34493 40655
rect 34549 40599 34705 40655
rect 34761 40599 34916 40655
rect 34972 40599 38328 40655
rect 38384 40599 38539 40655
rect 38595 40599 38750 40655
rect 38806 40599 40251 40655
rect 40307 40599 40431 40655
rect 40487 40599 43788 40655
rect 43844 40599 43999 40655
rect 44055 40599 44211 40655
rect 44267 40599 44422 40655
rect 44478 40599 50161 40655
rect 50217 40599 50372 40655
rect 50428 40599 50584 40655
rect 50640 40599 50795 40655
rect 50851 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 86372 40655
rect 0 40527 86372 40599
rect 0 40476 27272 40527
rect 30403 40526 54622 40527
rect 60471 40476 86372 40527
rect 0 40276 1014 40476
rect 37852 40379 48687 40417
rect 37852 40378 48594 40379
rect 37852 40322 37889 40378
rect 37945 40322 38069 40378
rect 38125 40322 39773 40378
rect 39829 40323 48594 40378
rect 48650 40323 48687 40379
rect 39829 40322 48687 40323
rect 37852 40284 48687 40322
rect 24298 40195 34090 40268
rect 24298 40188 33817 40195
rect 24298 40132 33055 40188
rect 33111 40132 33235 40188
rect 33291 40139 33817 40188
rect 33873 40139 33997 40195
rect 34053 40139 34090 40195
rect 33291 40132 34090 40139
rect 0 39376 1706 40076
rect 24298 40066 34090 40132
rect 36640 40147 40085 40186
rect 36640 40091 36676 40147
rect 36732 40091 39992 40147
rect 40048 40091 40085 40147
rect 36640 40053 40085 40091
rect 48557 40161 48687 40284
rect 85358 40276 86372 40476
rect 48557 40105 48594 40161
rect 48650 40105 48687 40161
rect 48557 40066 48687 40105
rect 51034 40195 60825 40268
rect 51034 40139 51071 40195
rect 51127 40139 51251 40195
rect 51307 40139 51833 40195
rect 51889 40139 52013 40195
rect 52069 40139 60825 40195
rect 51034 40066 60825 40139
rect 36648 40052 40041 40053
rect 24298 39755 60825 39828
rect 24298 39699 29580 39755
rect 29636 39699 29791 39755
rect 29847 39699 30003 39755
rect 30059 39699 30214 39755
rect 30270 39699 30852 39755
rect 30908 39699 31063 39755
rect 31119 39699 31274 39755
rect 31330 39699 31484 39755
rect 31540 39699 31695 39755
rect 31751 39699 31907 39755
rect 31963 39699 32118 39755
rect 32174 39699 32328 39755
rect 32384 39699 32539 39755
rect 32595 39699 32750 39755
rect 32806 39699 35218 39755
rect 35274 39699 35428 39755
rect 35484 39699 35639 39755
rect 35695 39699 35851 39755
rect 35907 39699 36062 39755
rect 36118 39699 36272 39755
rect 36328 39699 39050 39755
rect 39106 39699 39230 39755
rect 39286 39699 44832 39755
rect 44888 39699 45043 39755
rect 45099 39699 45254 39755
rect 45310 39699 48836 39755
rect 48892 39699 49046 39755
rect 49102 39699 49257 39755
rect 49313 39699 49469 39755
rect 49525 39699 49680 39755
rect 49736 39699 49890 39755
rect 49946 39699 52314 39755
rect 52370 39699 52525 39755
rect 52581 39699 52736 39755
rect 52792 39699 52946 39755
rect 53002 39699 53157 39755
rect 53213 39699 53369 39755
rect 53425 39699 53580 39755
rect 53636 39699 53790 39755
rect 53846 39699 54001 39755
rect 54057 39699 54212 39755
rect 54268 39699 54853 39755
rect 54909 39699 55064 39755
rect 55120 39699 55276 39755
rect 55332 39699 55487 39755
rect 55543 39699 60825 39755
rect 24298 39627 60825 39699
rect 30403 39626 54622 39627
rect 36648 39401 40041 39402
rect 24298 39322 34090 39388
rect 24298 39266 33055 39322
rect 33111 39266 33235 39322
rect 33291 39315 34090 39322
rect 33291 39266 33817 39315
rect 24298 39259 33817 39266
rect 33873 39259 33997 39315
rect 34053 39259 34090 39315
rect 36640 39363 40085 39401
rect 36640 39307 36676 39363
rect 36732 39307 39992 39363
rect 40048 39307 40085 39363
rect 36640 39268 40085 39307
rect 48557 39349 48687 39388
rect 48557 39293 48594 39349
rect 48650 39293 48687 39349
rect 24298 39187 34090 39259
rect 30403 39186 34090 39187
rect 0 38976 1014 39176
rect 48557 39170 48687 39293
rect 51034 39315 60825 39388
rect 84666 39376 86372 40076
rect 51034 39259 51071 39315
rect 51127 39259 51251 39315
rect 51307 39259 51833 39315
rect 51889 39259 52013 39315
rect 52069 39259 60825 39315
rect 51034 39187 60825 39259
rect 51034 39186 54622 39187
rect 37852 39132 48687 39170
rect 37852 39076 37889 39132
rect 37945 39076 38069 39132
rect 38125 39076 39773 39132
rect 39829 39131 48687 39132
rect 39829 39076 48594 39131
rect 37852 39075 48594 39076
rect 48650 39075 48687 39131
rect 37852 39037 48687 39075
rect 85358 38976 86372 39176
rect 0 38928 27272 38976
rect 60471 38928 86372 38976
rect 0 38855 86372 38928
rect 0 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 34282 38855
rect 34338 38799 34493 38855
rect 34549 38799 34705 38855
rect 34761 38799 34916 38855
rect 34972 38799 38328 38855
rect 38384 38799 38539 38855
rect 38595 38799 38750 38855
rect 38806 38799 40251 38855
rect 40307 38799 40431 38855
rect 40487 38799 43788 38855
rect 43844 38799 43999 38855
rect 44055 38799 44211 38855
rect 44267 38799 44422 38855
rect 44478 38799 50161 38855
rect 50217 38799 50372 38855
rect 50428 38799 50584 38855
rect 50640 38799 50795 38855
rect 50851 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 86372 38855
rect 0 38727 86372 38799
rect 0 38676 27272 38727
rect 30403 38726 54622 38727
rect 60471 38676 86372 38727
rect 0 38476 1014 38676
rect 37852 38579 48687 38617
rect 37852 38578 48594 38579
rect 37852 38522 37889 38578
rect 37945 38522 38069 38578
rect 38125 38522 39773 38578
rect 39829 38523 48594 38578
rect 48650 38523 48687 38579
rect 39829 38522 48687 38523
rect 37852 38484 48687 38522
rect 24298 38395 34090 38468
rect 24298 38388 33817 38395
rect 24298 38332 33055 38388
rect 33111 38332 33235 38388
rect 33291 38339 33817 38388
rect 33873 38339 33997 38395
rect 34053 38339 34090 38395
rect 33291 38332 34090 38339
rect 0 37576 1706 38276
rect 24298 38266 34090 38332
rect 36640 38347 40085 38386
rect 36640 38291 36676 38347
rect 36732 38291 39992 38347
rect 40048 38291 40085 38347
rect 36640 38253 40085 38291
rect 48557 38361 48687 38484
rect 85358 38476 86372 38676
rect 48557 38305 48594 38361
rect 48650 38305 48687 38361
rect 48557 38266 48687 38305
rect 51034 38395 60825 38468
rect 51034 38339 51071 38395
rect 51127 38339 51251 38395
rect 51307 38339 51833 38395
rect 51889 38339 52013 38395
rect 52069 38339 60825 38395
rect 51034 38266 60825 38339
rect 36648 38252 40041 38253
rect 24298 37955 60825 38028
rect 24298 37899 29580 37955
rect 29636 37899 29791 37955
rect 29847 37899 30003 37955
rect 30059 37899 30214 37955
rect 30270 37899 30852 37955
rect 30908 37899 31063 37955
rect 31119 37899 31274 37955
rect 31330 37899 31484 37955
rect 31540 37899 31695 37955
rect 31751 37899 31907 37955
rect 31963 37899 32118 37955
rect 32174 37899 32328 37955
rect 32384 37899 32539 37955
rect 32595 37899 32750 37955
rect 32806 37899 35218 37955
rect 35274 37899 35428 37955
rect 35484 37899 35639 37955
rect 35695 37899 35851 37955
rect 35907 37899 36062 37955
rect 36118 37899 36272 37955
rect 36328 37899 39050 37955
rect 39106 37899 39230 37955
rect 39286 37899 44832 37955
rect 44888 37899 45043 37955
rect 45099 37899 45254 37955
rect 45310 37899 48836 37955
rect 48892 37899 49046 37955
rect 49102 37899 49257 37955
rect 49313 37899 49469 37955
rect 49525 37899 49680 37955
rect 49736 37899 49890 37955
rect 49946 37899 52314 37955
rect 52370 37899 52525 37955
rect 52581 37899 52736 37955
rect 52792 37899 52946 37955
rect 53002 37899 53157 37955
rect 53213 37899 53369 37955
rect 53425 37899 53580 37955
rect 53636 37899 53790 37955
rect 53846 37899 54001 37955
rect 54057 37899 54212 37955
rect 54268 37899 54853 37955
rect 54909 37899 55064 37955
rect 55120 37899 55276 37955
rect 55332 37899 55487 37955
rect 55543 37899 60825 37955
rect 24298 37827 60825 37899
rect 30403 37826 54622 37827
rect 36648 37601 40041 37602
rect 24298 37522 34090 37588
rect 24298 37466 33055 37522
rect 33111 37466 33235 37522
rect 33291 37515 34090 37522
rect 33291 37466 33817 37515
rect 24298 37459 33817 37466
rect 33873 37459 33997 37515
rect 34053 37459 34090 37515
rect 36640 37563 40085 37601
rect 36640 37507 36676 37563
rect 36732 37507 39992 37563
rect 40048 37507 40085 37563
rect 36640 37468 40085 37507
rect 48557 37549 48687 37588
rect 48557 37493 48594 37549
rect 48650 37493 48687 37549
rect 24298 37387 34090 37459
rect 30403 37386 34090 37387
rect 0 37176 1014 37376
rect 48557 37370 48687 37493
rect 51034 37515 60825 37588
rect 84666 37576 86372 38276
rect 51034 37459 51071 37515
rect 51127 37459 51251 37515
rect 51307 37459 51833 37515
rect 51889 37459 52013 37515
rect 52069 37459 60825 37515
rect 51034 37387 60825 37459
rect 51034 37386 54622 37387
rect 37852 37332 48687 37370
rect 37852 37276 37889 37332
rect 37945 37276 38069 37332
rect 38125 37276 39773 37332
rect 39829 37331 48687 37332
rect 39829 37276 48594 37331
rect 37852 37275 48594 37276
rect 48650 37275 48687 37331
rect 37852 37237 48687 37275
rect 85358 37176 86372 37376
rect 0 37128 27272 37176
rect 60471 37128 86372 37176
rect 0 37055 86372 37128
rect 0 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 34282 37055
rect 34338 36999 34493 37055
rect 34549 36999 34705 37055
rect 34761 36999 34916 37055
rect 34972 36999 38328 37055
rect 38384 36999 38539 37055
rect 38595 36999 38750 37055
rect 38806 36999 40251 37055
rect 40307 36999 40431 37055
rect 40487 36999 43788 37055
rect 43844 36999 43999 37055
rect 44055 36999 44211 37055
rect 44267 36999 44422 37055
rect 44478 36999 50161 37055
rect 50217 36999 50372 37055
rect 50428 36999 50584 37055
rect 50640 36999 50795 37055
rect 50851 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 86372 37055
rect 0 36927 86372 36999
rect 0 36876 27272 36927
rect 30403 36926 54622 36927
rect 60471 36876 86372 36927
rect 0 36676 1014 36876
rect 37852 36779 48687 36817
rect 37852 36778 48594 36779
rect 37852 36722 37889 36778
rect 37945 36722 38069 36778
rect 38125 36722 39773 36778
rect 39829 36723 48594 36778
rect 48650 36723 48687 36779
rect 39829 36722 48687 36723
rect 37852 36684 48687 36722
rect 24298 36595 34090 36668
rect 24298 36588 33817 36595
rect 24298 36532 33055 36588
rect 33111 36532 33235 36588
rect 33291 36539 33817 36588
rect 33873 36539 33997 36595
rect 34053 36539 34090 36595
rect 33291 36532 34090 36539
rect 0 35776 1706 36476
rect 24298 36466 34090 36532
rect 36640 36547 40085 36586
rect 36640 36491 36676 36547
rect 36732 36491 39992 36547
rect 40048 36491 40085 36547
rect 36640 36453 40085 36491
rect 48557 36561 48687 36684
rect 85358 36676 86372 36876
rect 48557 36505 48594 36561
rect 48650 36505 48687 36561
rect 48557 36466 48687 36505
rect 51034 36595 60825 36668
rect 51034 36539 51071 36595
rect 51127 36539 51251 36595
rect 51307 36539 51833 36595
rect 51889 36539 52013 36595
rect 52069 36539 60825 36595
rect 51034 36466 60825 36539
rect 36648 36452 40041 36453
rect 24298 36155 60825 36228
rect 24298 36099 29580 36155
rect 29636 36099 29791 36155
rect 29847 36099 30003 36155
rect 30059 36099 30214 36155
rect 30270 36099 30852 36155
rect 30908 36099 31063 36155
rect 31119 36099 31274 36155
rect 31330 36099 31484 36155
rect 31540 36099 31695 36155
rect 31751 36099 31907 36155
rect 31963 36099 32118 36155
rect 32174 36099 32328 36155
rect 32384 36099 32539 36155
rect 32595 36099 32750 36155
rect 32806 36099 35218 36155
rect 35274 36099 35428 36155
rect 35484 36099 35639 36155
rect 35695 36099 35851 36155
rect 35907 36099 36062 36155
rect 36118 36099 36272 36155
rect 36328 36099 39050 36155
rect 39106 36099 39230 36155
rect 39286 36099 44832 36155
rect 44888 36099 45043 36155
rect 45099 36099 45254 36155
rect 45310 36099 48836 36155
rect 48892 36099 49046 36155
rect 49102 36099 49257 36155
rect 49313 36099 49469 36155
rect 49525 36099 49680 36155
rect 49736 36099 49890 36155
rect 49946 36099 52314 36155
rect 52370 36099 52525 36155
rect 52581 36099 52736 36155
rect 52792 36099 52946 36155
rect 53002 36099 53157 36155
rect 53213 36099 53369 36155
rect 53425 36099 53580 36155
rect 53636 36099 53790 36155
rect 53846 36099 54001 36155
rect 54057 36099 54212 36155
rect 54268 36099 54853 36155
rect 54909 36099 55064 36155
rect 55120 36099 55276 36155
rect 55332 36099 55487 36155
rect 55543 36099 60825 36155
rect 24298 36027 60825 36099
rect 30403 36026 54622 36027
rect 36863 35881 37743 35920
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 0 35126 24917 35326
rect 0 35016 1014 35126
rect 27442 35024 27782 35062
rect 27442 35016 27478 35024
rect 0 34968 27478 35016
rect 27534 34968 27690 35024
rect 27746 35016 27782 35024
rect 27746 34968 27830 35016
rect 0 34961 27830 34968
rect 0 34905 25344 34961
rect 25400 34905 25468 34961
rect 25524 34905 25592 34961
rect 25648 34905 25716 34961
rect 25772 34905 25840 34961
rect 25896 34905 25964 34961
rect 26020 34905 27830 34961
rect 0 34837 27830 34905
rect 0 34781 25344 34837
rect 25400 34781 25468 34837
rect 25524 34781 25592 34837
rect 25648 34781 25716 34837
rect 25772 34781 25840 34837
rect 25896 34781 25964 34837
rect 26020 34806 27830 34837
rect 26020 34781 27478 34806
rect 0 34750 27478 34781
rect 27534 34750 27690 34806
rect 27746 34750 27830 34806
rect 0 34713 27830 34750
rect 0 34657 25344 34713
rect 25400 34657 25468 34713
rect 25524 34657 25592 34713
rect 25648 34657 25716 34713
rect 25772 34657 25840 34713
rect 25896 34657 25964 34713
rect 26020 34657 27830 34713
rect 0 34588 27830 34657
rect 0 34536 27478 34588
rect 27442 34532 27478 34536
rect 27534 34532 27690 34588
rect 27746 34536 27830 34588
rect 27746 34532 27782 34536
rect 27442 34494 27782 34532
rect 2095 34125 2188 34126
rect 0 34124 25085 34125
rect 0 34011 27214 34124
rect 0 33955 26859 34011
rect 26915 33955 27071 34011
rect 27127 33955 27214 34011
rect 0 33793 27214 33955
rect 36863 33927 37743 35825
rect 84666 35776 86372 36476
rect 60559 35298 60647 35387
rect 83360 35298 86372 35326
rect 60282 35158 86372 35298
rect 60559 35016 60647 35158
rect 83360 35126 86372 35158
rect 85358 35016 86372 35126
rect 58812 34981 59508 34991
rect 58812 34925 58822 34981
rect 58878 34925 58946 34981
rect 59002 34925 59070 34981
rect 59126 34925 59194 34981
rect 59250 34925 59318 34981
rect 59374 34925 59442 34981
rect 59498 34925 59508 34981
rect 58812 34857 59508 34925
rect 58812 34801 58822 34857
rect 58878 34801 58946 34857
rect 59002 34801 59070 34857
rect 59126 34801 59194 34857
rect 59250 34801 59318 34857
rect 59374 34801 59442 34857
rect 59498 34801 59508 34857
rect 58812 34733 59508 34801
rect 58812 34677 58822 34733
rect 58878 34677 58946 34733
rect 59002 34677 59070 34733
rect 59126 34677 59194 34733
rect 59250 34677 59318 34733
rect 59374 34677 59442 34733
rect 59498 34677 59508 34733
rect 58812 34667 59508 34677
rect 60282 34536 86372 35016
rect 61853 34124 72383 34125
rect 72653 34124 86372 34125
rect 57908 34011 86372 34124
rect 57908 33955 57996 34011
rect 58052 33955 58208 34011
rect 58264 33955 86372 34011
rect 0 33737 26859 33793
rect 26915 33737 27071 33793
rect 27127 33737 27214 33793
rect 0 33576 27214 33737
rect 0 33520 26859 33576
rect 26915 33520 27071 33576
rect 27127 33520 27214 33576
rect 0 33358 27214 33520
rect 0 33302 26859 33358
rect 26915 33302 27071 33358
rect 27127 33302 27214 33358
rect 0 33140 27214 33302
rect 57908 33793 86372 33955
rect 57908 33737 57996 33793
rect 58052 33737 58208 33793
rect 58264 33737 86372 33793
rect 57908 33576 86372 33737
rect 57908 33520 57996 33576
rect 58052 33520 58208 33576
rect 58264 33520 86372 33576
rect 57908 33358 86372 33520
rect 57908 33302 57996 33358
rect 58052 33302 58208 33358
rect 58264 33302 86372 33358
rect 0 33084 26859 33140
rect 26915 33084 27071 33140
rect 27127 33084 27214 33140
rect 0 32922 27214 33084
rect 0 32866 26859 32922
rect 26915 32866 27071 32922
rect 27127 32866 27214 32922
rect 0 32705 27214 32866
rect 0 32649 26859 32705
rect 26915 32649 27071 32705
rect 27127 32649 27214 32705
rect 0 32487 27214 32649
rect 0 32431 26859 32487
rect 26915 32431 27071 32487
rect 27127 32431 27214 32487
rect 0 32318 27214 32431
rect 27387 33141 28929 33263
rect 27387 33085 27474 33141
rect 27530 33085 27686 33141
rect 27742 33085 28929 33141
rect 27387 32923 28929 33085
rect 27387 32867 27474 32923
rect 27530 32867 27686 32923
rect 27742 32867 28929 32923
rect 27387 32705 28929 32867
rect 27387 32649 27474 32705
rect 27530 32649 27686 32705
rect 27742 32649 28929 32705
rect 27387 32487 28929 32649
rect 27387 32431 27474 32487
rect 27530 32431 27686 32487
rect 27742 32431 28929 32487
rect 0 32316 25085 32318
rect 0 32315 3011 32316
rect 0 29714 1706 32315
rect 27387 32311 28929 32431
rect 56135 33141 57736 33263
rect 56135 33085 57381 33141
rect 57437 33085 57593 33141
rect 57649 33085 57736 33141
rect 56135 32923 57736 33085
rect 56135 32867 57381 32923
rect 57437 32867 57593 32923
rect 57649 32867 57736 32923
rect 56135 32705 57736 32867
rect 56135 32649 57381 32705
rect 57437 32649 57593 32705
rect 57649 32649 57736 32705
rect 56135 32487 57736 32649
rect 56135 32431 57381 32487
rect 57437 32431 57593 32487
rect 57649 32431 57736 32487
rect 56135 32311 57736 32431
rect 57908 33140 86372 33302
rect 57908 33084 57996 33140
rect 58052 33084 58208 33140
rect 58264 33084 86372 33140
rect 57908 32922 86372 33084
rect 57908 32866 57996 32922
rect 58052 32866 58208 32922
rect 58264 32866 86372 32922
rect 57908 32705 86372 32866
rect 57908 32649 57996 32705
rect 58052 32649 58208 32705
rect 58264 32649 86372 32705
rect 57908 32487 86372 32649
rect 57908 32431 57996 32487
rect 58052 32431 58208 32487
rect 58264 32431 86372 32487
rect 57908 32315 86372 32431
rect 57908 32199 58351 32315
rect 26772 32088 58351 32199
rect 26772 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 26772 31870 58351 32032
rect 26772 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 26772 31652 58351 31814
rect 26772 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 26772 31486 58351 31596
rect 25293 31252 28929 31352
rect 25293 31248 27474 31252
rect 25293 31192 25398 31248
rect 25454 31192 25522 31248
rect 25578 31192 25646 31248
rect 25702 31192 25770 31248
rect 25826 31192 25894 31248
rect 25950 31196 27474 31248
rect 27530 31196 27686 31252
rect 27742 31196 28929 31252
rect 25950 31192 28929 31196
rect 25293 31124 28929 31192
rect 25293 31068 25398 31124
rect 25454 31068 25522 31124
rect 25578 31068 25646 31124
rect 25702 31068 25770 31124
rect 25826 31068 25894 31124
rect 25950 31068 28929 31124
rect 25293 31034 28929 31068
rect 25293 31000 27474 31034
rect 25293 30944 25398 31000
rect 25454 30944 25522 31000
rect 25578 30944 25646 31000
rect 25702 30944 25770 31000
rect 25826 30944 25894 31000
rect 25950 30978 27474 31000
rect 27530 30978 27686 31034
rect 27742 30978 28929 31034
rect 25950 30944 28929 30978
rect 25293 30816 28929 30944
rect 25293 30793 27474 30816
rect 25293 30737 25398 30793
rect 25454 30737 25522 30793
rect 25578 30737 25646 30793
rect 25702 30737 25770 30793
rect 25826 30737 25894 30793
rect 25950 30760 27474 30793
rect 27530 30760 27686 30816
rect 27742 30760 28929 30816
rect 25950 30737 28929 30760
rect 25293 30669 28929 30737
rect 25293 30613 25398 30669
rect 25454 30613 25522 30669
rect 25578 30613 25646 30669
rect 25702 30613 25770 30669
rect 25826 30613 25894 30669
rect 25950 30613 28929 30669
rect 25293 30598 28929 30613
rect 25293 30545 27474 30598
rect 25293 30489 25398 30545
rect 25454 30489 25522 30545
rect 25578 30489 25646 30545
rect 25702 30489 25770 30545
rect 25826 30489 25894 30545
rect 25950 30542 27474 30545
rect 27530 30542 27686 30598
rect 27742 30542 28929 30598
rect 25950 30489 28929 30542
rect 25293 30443 28929 30489
rect 56186 31298 59524 31352
rect 56186 31252 58873 31298
rect 56186 31196 57381 31252
rect 57437 31196 57593 31252
rect 57649 31242 58873 31252
rect 58929 31242 58997 31298
rect 59053 31242 59121 31298
rect 59177 31242 59245 31298
rect 59301 31242 59369 31298
rect 59425 31242 59524 31298
rect 57649 31196 59524 31242
rect 56186 31174 59524 31196
rect 56186 31118 58873 31174
rect 58929 31118 58997 31174
rect 59053 31118 59121 31174
rect 59177 31118 59245 31174
rect 59301 31118 59369 31174
rect 59425 31118 59524 31174
rect 56186 31050 59524 31118
rect 56186 31034 58873 31050
rect 56186 30978 57381 31034
rect 57437 30978 57593 31034
rect 57649 30994 58873 31034
rect 58929 30994 58997 31050
rect 59053 30994 59121 31050
rect 59177 30994 59245 31050
rect 59301 30994 59369 31050
rect 59425 30994 59524 31050
rect 57649 30978 59524 30994
rect 56186 30853 59524 30978
rect 56186 30816 58873 30853
rect 56186 30760 57381 30816
rect 57437 30760 57593 30816
rect 57649 30797 58873 30816
rect 58929 30797 58997 30853
rect 59053 30797 59121 30853
rect 59177 30797 59245 30853
rect 59301 30797 59369 30853
rect 59425 30797 59524 30853
rect 57649 30760 59524 30797
rect 56186 30729 59524 30760
rect 56186 30673 58873 30729
rect 58929 30673 58997 30729
rect 59053 30673 59121 30729
rect 59177 30673 59245 30729
rect 59301 30673 59369 30729
rect 59425 30673 59524 30729
rect 56186 30605 59524 30673
rect 56186 30598 58873 30605
rect 56186 30542 57381 30598
rect 57437 30542 57593 30598
rect 57649 30549 58873 30598
rect 58929 30549 58997 30605
rect 59053 30549 59121 30605
rect 59177 30549 59245 30605
rect 59301 30549 59369 30605
rect 59425 30549 59524 30605
rect 57649 30542 59524 30549
rect 56186 30443 59524 30542
rect 26772 29968 58351 30105
rect 26772 29912 26859 29968
rect 26915 29912 27071 29968
rect 27127 29912 57996 29968
rect 58052 29912 58208 29968
rect 58264 29912 58351 29968
rect 26772 29750 58351 29912
rect 26772 29714 26859 29750
rect 0 29694 26859 29714
rect 26915 29694 27071 29750
rect 27127 29694 57996 29750
rect 58052 29694 58208 29750
rect 58264 29714 58351 29750
rect 84666 29714 86372 32315
rect 58264 29694 86372 29714
rect 0 29533 86372 29694
rect 0 29477 26859 29533
rect 26915 29477 27071 29533
rect 27127 29477 57996 29533
rect 58052 29477 58208 29533
rect 58264 29477 86372 29533
rect 0 29430 86372 29477
rect 26772 29315 58351 29430
rect 26772 29259 26859 29315
rect 26915 29259 27071 29315
rect 27127 29259 57996 29315
rect 58052 29259 58208 29315
rect 58264 29259 58351 29315
rect 26772 29098 58351 29259
rect 26772 29042 26859 29098
rect 26915 29042 27071 29098
rect 27127 29042 57996 29098
rect 58052 29042 58208 29098
rect 58264 29042 58351 29098
rect 26772 28880 58351 29042
rect 26772 28824 26859 28880
rect 26915 28824 27071 28880
rect 27127 28824 57996 28880
rect 58052 28824 58208 28880
rect 58264 28824 58351 28880
rect 26772 28662 58351 28824
rect 26772 28606 26859 28662
rect 26915 28606 27071 28662
rect 27127 28606 57996 28662
rect 58052 28606 58208 28662
rect 58264 28606 58351 28662
rect 26772 28444 58351 28606
rect 1954 28416 26070 28434
rect 0 28315 26070 28416
rect 0 28259 25404 28315
rect 25460 28259 25528 28315
rect 25584 28259 25652 28315
rect 25708 28259 25776 28315
rect 25832 28259 25900 28315
rect 25956 28259 26070 28315
rect 0 28191 26070 28259
rect 0 28135 25404 28191
rect 25460 28135 25528 28191
rect 25584 28135 25652 28191
rect 25708 28135 25776 28191
rect 25832 28135 25900 28191
rect 25956 28135 26070 28191
rect 0 28067 26070 28135
rect 0 28011 25404 28067
rect 25460 28011 25528 28067
rect 25584 28011 25652 28067
rect 25708 28011 25776 28067
rect 25832 28011 25900 28067
rect 25956 28011 26070 28067
rect 0 27943 26070 28011
rect 0 27887 25404 27943
rect 25460 27887 25528 27943
rect 25584 27887 25652 27943
rect 25708 27887 25776 27943
rect 25832 27887 25900 27943
rect 25956 27887 26070 27943
rect 0 27819 26070 27887
rect 0 27763 25404 27819
rect 25460 27763 25528 27819
rect 25584 27763 25652 27819
rect 25708 27763 25776 27819
rect 25832 27763 25900 27819
rect 25956 27763 26070 27819
rect 0 27695 26070 27763
rect 0 27639 25404 27695
rect 25460 27639 25528 27695
rect 25584 27639 25652 27695
rect 25708 27639 25776 27695
rect 25832 27639 25900 27695
rect 25956 27639 26070 27695
rect 0 27571 26070 27639
rect 0 27515 25404 27571
rect 25460 27515 25528 27571
rect 25584 27515 25652 27571
rect 25708 27515 25776 27571
rect 25832 27515 25900 27571
rect 25956 27515 26070 27571
rect 0 27447 26070 27515
rect 0 27391 25404 27447
rect 25460 27391 25528 27447
rect 25584 27391 25652 27447
rect 25708 27391 25776 27447
rect 25832 27391 25900 27447
rect 25956 27391 26070 27447
rect 0 27323 26070 27391
rect 26772 28388 26859 28444
rect 26915 28388 27071 28444
rect 27127 28388 57996 28444
rect 58052 28388 58208 28444
rect 58264 28388 58351 28444
rect 26772 28227 58351 28388
rect 26772 28171 26859 28227
rect 26915 28171 27071 28227
rect 27127 28171 57996 28227
rect 58052 28171 58208 28227
rect 58264 28171 58351 28227
rect 26772 28009 58351 28171
rect 26772 27953 26859 28009
rect 26915 27953 27071 28009
rect 27127 27953 57996 28009
rect 58052 27953 58208 28009
rect 58264 27953 58351 28009
rect 26772 27792 58351 27953
rect 26772 27736 26859 27792
rect 26915 27736 27071 27792
rect 27127 27736 57996 27792
rect 58052 27736 58208 27792
rect 58264 27736 58351 27792
rect 26772 27574 58351 27736
rect 26772 27518 26859 27574
rect 26915 27518 27071 27574
rect 27127 27518 57996 27574
rect 58052 27518 58208 27574
rect 58264 27518 58351 27574
rect 26772 27382 58351 27518
rect 58785 28416 84717 28434
rect 58785 28321 86372 28416
rect 58785 28265 58859 28321
rect 58915 28265 58983 28321
rect 59039 28265 59107 28321
rect 59163 28265 59231 28321
rect 59287 28265 59355 28321
rect 59411 28265 86372 28321
rect 58785 28197 86372 28265
rect 58785 28141 58859 28197
rect 58915 28141 58983 28197
rect 59039 28141 59107 28197
rect 59163 28141 59231 28197
rect 59287 28141 59355 28197
rect 59411 28141 86372 28197
rect 58785 28073 86372 28141
rect 58785 28017 58859 28073
rect 58915 28017 58983 28073
rect 59039 28017 59107 28073
rect 59163 28017 59231 28073
rect 59287 28017 59355 28073
rect 59411 28017 86372 28073
rect 58785 27949 86372 28017
rect 58785 27893 58859 27949
rect 58915 27893 58983 27949
rect 59039 27893 59107 27949
rect 59163 27893 59231 27949
rect 59287 27893 59355 27949
rect 59411 27893 86372 27949
rect 58785 27825 86372 27893
rect 58785 27769 58859 27825
rect 58915 27769 58983 27825
rect 59039 27769 59107 27825
rect 59163 27769 59231 27825
rect 59287 27769 59355 27825
rect 59411 27769 86372 27825
rect 58785 27701 86372 27769
rect 58785 27645 58859 27701
rect 58915 27645 58983 27701
rect 59039 27645 59107 27701
rect 59163 27645 59231 27701
rect 59287 27645 59355 27701
rect 59411 27645 86372 27701
rect 58785 27577 86372 27645
rect 58785 27521 58859 27577
rect 58915 27521 58983 27577
rect 59039 27521 59107 27577
rect 59163 27521 59231 27577
rect 59287 27521 59355 27577
rect 59411 27521 86372 27577
rect 58785 27453 86372 27521
rect 58785 27397 58859 27453
rect 58915 27397 58983 27453
rect 59039 27397 59107 27453
rect 59163 27397 59231 27453
rect 59287 27397 59355 27453
rect 59411 27397 86372 27453
rect 0 27267 25404 27323
rect 25460 27267 25528 27323
rect 25584 27267 25652 27323
rect 25708 27267 25776 27323
rect 25832 27267 25900 27323
rect 25956 27267 26070 27323
rect 0 27199 26070 27267
rect 0 27143 25404 27199
rect 25460 27143 25528 27199
rect 25584 27143 25652 27199
rect 25708 27143 25776 27199
rect 25832 27143 25900 27199
rect 25956 27143 26070 27199
rect 0 27075 26070 27143
rect 0 27019 25404 27075
rect 25460 27019 25528 27075
rect 25584 27019 25652 27075
rect 25708 27019 25776 27075
rect 25832 27019 25900 27075
rect 25956 27019 26070 27075
rect 0 26951 26070 27019
rect 0 26895 25404 26951
rect 25460 26895 25528 26951
rect 25584 26895 25652 26951
rect 25708 26895 25776 26951
rect 25832 26895 25900 26951
rect 25956 26895 26070 26951
rect 0 26890 26070 26895
rect 58785 27329 86372 27397
rect 58785 27273 58859 27329
rect 58915 27273 58983 27329
rect 59039 27273 59107 27329
rect 59163 27273 59231 27329
rect 59287 27273 59355 27329
rect 59411 27273 86372 27329
rect 58785 27205 86372 27273
rect 58785 27149 58859 27205
rect 58915 27149 58983 27205
rect 59039 27149 59107 27205
rect 59163 27149 59231 27205
rect 59287 27149 59355 27205
rect 59411 27149 86372 27205
rect 58785 27081 86372 27149
rect 58785 27025 58859 27081
rect 58915 27025 58983 27081
rect 59039 27025 59107 27081
rect 59163 27025 59231 27081
rect 59287 27025 59355 27081
rect 59411 27025 86372 27081
rect 58785 26957 86372 27025
rect 58785 26901 58859 26957
rect 58915 26901 58983 26957
rect 59039 26901 59107 26957
rect 59163 26901 59231 26957
rect 59287 26901 59355 26957
rect 59411 26901 86372 26957
rect 58785 26890 86372 26901
rect 0 26827 27828 26890
rect 0 26771 25404 26827
rect 25460 26771 25528 26827
rect 25584 26771 25652 26827
rect 25708 26771 25776 26827
rect 25832 26771 25900 26827
rect 25956 26799 27828 26827
rect 25956 26771 27474 26799
rect 0 26743 27474 26771
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 0 26703 27828 26743
rect 0 26647 25404 26703
rect 25460 26647 25528 26703
rect 25584 26647 25652 26703
rect 25708 26647 25776 26703
rect 25832 26647 25900 26703
rect 25956 26647 27828 26703
rect 0 26581 27828 26647
rect 0 26579 27474 26581
rect 0 26523 25404 26579
rect 25460 26523 25528 26579
rect 25584 26523 25652 26579
rect 25708 26523 25776 26579
rect 25832 26523 25900 26579
rect 25956 26525 27474 26579
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 25956 26523 27828 26525
rect 0 26435 27828 26523
rect 57295 26833 86372 26890
rect 57295 26799 58859 26833
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26777 58859 26799
rect 58915 26777 58983 26833
rect 59039 26777 59107 26833
rect 59163 26777 59231 26833
rect 59287 26777 59355 26833
rect 59411 26777 86372 26833
rect 57649 26743 86372 26777
rect 57295 26709 86372 26743
rect 57295 26653 58859 26709
rect 58915 26653 58983 26709
rect 59039 26653 59107 26709
rect 59163 26653 59231 26709
rect 59287 26653 59355 26709
rect 59411 26653 86372 26709
rect 57295 26585 86372 26653
rect 57295 26581 58859 26585
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26529 58859 26581
rect 58915 26529 58983 26585
rect 59039 26529 59107 26585
rect 59163 26529 59231 26585
rect 59287 26529 59355 26585
rect 59411 26529 86372 26585
rect 57649 26525 86372 26529
rect 57295 26435 86372 26525
rect 23828 26286 26642 26324
rect 23828 26126 26450 26286
rect 26610 26126 26642 26286
rect 23828 26109 26642 26126
rect 23828 25967 26285 26002
rect 23828 25807 26092 25967
rect 26252 25807 26285 25967
rect 23828 25787 26285 25807
rect 23828 25647 25949 25681
rect 23828 25487 25756 25647
rect 25916 25487 25949 25647
rect 23828 25466 25949 25487
rect 23828 25328 25614 25359
rect 23828 25168 25421 25328
rect 25581 25168 25614 25328
rect 23828 25144 25614 25168
rect 27382 25028 29699 25208
rect 27382 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 29699 25028
rect 27382 24810 29699 24972
rect 27382 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 29699 24810
rect 23828 24637 25274 24667
rect 23828 24477 25081 24637
rect 25241 24477 25274 24637
rect 27382 24526 29699 24754
rect 23828 24452 25274 24477
rect 23828 24316 24935 24345
rect 23828 24156 24744 24316
rect 24904 24156 24935 24316
rect 23828 24130 24935 24156
rect 26770 24075 58348 24278
rect 23828 23995 24607 24024
rect 0 23380 1706 23938
rect 23828 23835 24416 23995
rect 24576 23835 24607 23995
rect 23828 23809 24607 23835
rect 24047 23673 24227 23683
rect 24047 23513 24057 23673
rect 24217 23513 24227 23673
rect 24047 23503 24227 23513
rect 26770 23380 26858 24075
rect 0 23187 26858 23380
rect 27122 23370 57994 24075
rect 27122 23187 27214 23370
rect 0 22938 27214 23187
rect 27387 22936 57677 23199
rect 57908 23187 57994 23370
rect 58258 23380 58348 24075
rect 84666 23380 86372 23938
rect 58258 23187 86372 23380
rect 57908 22938 86372 23187
rect 57908 22937 83763 22938
rect 27387 22282 27475 22936
rect 0 22048 27475 22282
rect 27739 22923 57677 22936
rect 27739 22291 57363 22923
rect 27739 22048 27826 22291
rect 0 21827 27826 22048
rect 0 21282 1014 21827
rect 24036 21826 27826 21827
rect 56078 22035 57363 22291
rect 57627 22282 57677 22923
rect 57627 22035 86372 22282
rect 56078 21827 86372 22035
rect 56078 21826 83763 21827
rect 44432 21707 55645 21708
rect 29521 21625 55645 21707
rect 29513 20739 55645 21625
rect 85358 21282 86372 21827
rect 0 20570 86372 20739
rect 0 20410 26924 20570
rect 27084 20410 58048 20570
rect 58208 20410 86372 20570
rect 0 20226 86372 20410
rect 0 20066 26924 20226
rect 27084 20066 58048 20226
rect 58208 20066 86372 20226
rect 0 19969 86372 20066
rect 0 18016 24250 19969
rect 26435 19692 29403 19731
rect 26435 19532 26465 19692
rect 26625 19532 29403 19692
rect 26435 19502 29403 19532
rect 55720 19502 58817 19731
rect 26077 19347 29403 19391
rect 26077 19187 26107 19347
rect 26267 19187 29403 19347
rect 26077 19162 29403 19187
rect 55720 19162 59177 19391
rect 25742 19027 29403 19051
rect 25742 18867 25771 19027
rect 25931 18867 29403 19027
rect 25742 18822 29403 18867
rect 55720 18822 59515 19051
rect 25406 18684 29403 18711
rect 25406 18524 25434 18684
rect 25594 18524 29403 18684
rect 25406 18482 29403 18524
rect 55720 18482 59846 18711
rect 25066 18350 29403 18371
rect 25066 18190 25094 18350
rect 25254 18190 29403 18350
rect 25066 18142 29403 18190
rect 55720 18142 60184 18371
rect 24730 17977 29403 18031
rect 24730 17817 24757 17977
rect 24917 17817 29403 17977
rect 24730 17802 29403 17817
rect 55720 17802 60525 18031
rect 61502 18016 86372 19969
rect 61502 18015 83763 18016
rect 0 16597 23678 17730
rect 24401 17656 29403 17691
rect 24401 17496 24429 17656
rect 24589 17496 29403 17656
rect 24401 17462 29403 17496
rect 55720 17462 60855 17691
rect 24042 17317 29403 17351
rect 24042 17157 24069 17317
rect 24229 17157 29403 17317
rect 24042 17122 29403 17157
rect 55720 17122 61205 17351
rect 61760 16784 86372 17730
rect 46982 16678 86372 16784
rect 46982 16622 57381 16678
rect 57437 16622 57593 16678
rect 57649 16622 86372 16678
rect 24111 16597 27828 16598
rect 0 16470 27828 16597
rect 0 16414 27474 16470
rect 27530 16414 27686 16470
rect 27742 16414 27828 16470
rect 0 16253 27828 16414
rect 0 16197 27474 16253
rect 27530 16197 27686 16253
rect 27742 16197 27828 16253
rect 0 16035 27828 16197
rect 0 15979 27474 16035
rect 27530 15979 27686 16035
rect 27742 15979 27828 16035
rect 0 15818 27828 15979
rect 0 15762 27474 15818
rect 27530 15762 27686 15818
rect 27742 15762 27828 15818
rect 0 15600 27828 15762
rect 0 15544 27474 15600
rect 27530 15544 27686 15600
rect 27742 15544 27828 15600
rect 0 15382 27828 15544
rect 0 15326 27474 15382
rect 27530 15326 27686 15382
rect 27742 15326 27828 15382
rect 0 15164 27828 15326
rect 0 15108 27474 15164
rect 27530 15108 27686 15164
rect 27742 15108 27828 15164
rect 0 15015 27828 15108
rect 46982 16461 86372 16622
rect 46982 16405 57381 16461
rect 57437 16405 57593 16461
rect 57649 16405 86372 16461
rect 46982 16243 86372 16405
rect 46982 16187 57381 16243
rect 57437 16187 57593 16243
rect 57649 16187 86372 16243
rect 46982 16026 86372 16187
rect 46982 15970 57381 16026
rect 57437 15970 57593 16026
rect 57649 15970 86372 16026
rect 46982 15808 86372 15970
rect 46982 15752 57381 15808
rect 57437 15752 57593 15808
rect 57649 15752 86372 15808
rect 46982 15590 86372 15752
rect 46982 15534 57381 15590
rect 57437 15534 57593 15590
rect 57649 15534 86372 15590
rect 46982 15372 86372 15534
rect 46982 15316 57381 15372
rect 57437 15316 57593 15372
rect 57649 15316 86372 15372
rect 46982 15155 86372 15316
rect 46982 15099 57381 15155
rect 57437 15099 57593 15155
rect 57649 15099 86372 15155
rect 46982 15015 86372 15099
rect 0 14968 86372 15015
rect 0 14966 55645 14968
rect 0 14947 51760 14966
rect 0 14891 27474 14947
rect 27530 14891 27686 14947
rect 27742 14936 51760 14947
rect 57295 14937 86372 14968
rect 27742 14891 47683 14936
rect 0 14729 47683 14891
rect 0 14673 27474 14729
rect 27530 14673 27686 14729
rect 27742 14673 47683 14729
rect 0 14512 47683 14673
rect 0 14456 27474 14512
rect 27530 14456 27686 14512
rect 27742 14491 47683 14512
rect 57295 14881 57381 14937
rect 57437 14881 57593 14937
rect 57649 14881 86372 14937
rect 57295 14720 86372 14881
rect 57295 14664 57381 14720
rect 57437 14664 57593 14720
rect 57649 14664 86372 14720
rect 27742 14456 45977 14491
rect 0 14329 45977 14456
rect 0 14328 24250 14329
rect 27387 14231 45977 14329
rect 57295 14328 86372 14664
rect 57295 14327 83763 14328
rect 24047 14178 27214 14179
rect 0 14119 27214 14178
rect 0 14063 26859 14119
rect 26915 14063 27071 14119
rect 27127 14063 27214 14119
rect 0 13902 27214 14063
rect 0 13846 26859 13902
rect 26915 13846 27071 13902
rect 27127 13846 27214 13902
rect 0 13684 27214 13846
rect 0 13628 26859 13684
rect 26915 13628 27071 13684
rect 27127 13628 27214 13684
rect 0 13467 27214 13628
rect 0 13461 26859 13467
rect 0 12846 1706 13461
rect 24047 13411 26859 13461
rect 26915 13411 27071 13467
rect 27127 13411 27214 13467
rect 24047 13249 27214 13411
rect 24047 13193 26859 13249
rect 26915 13193 27071 13249
rect 27127 13193 27214 13249
rect 27387 14175 27474 14231
rect 27530 14175 27686 14231
rect 27742 14175 45977 14231
rect 83169 14178 84221 14179
rect 61807 14177 72429 14178
rect 72607 14177 86372 14178
rect 27387 14014 45977 14175
rect 27387 13958 27474 14014
rect 27530 13958 27686 14014
rect 27742 13958 45977 14014
rect 27387 13796 45977 13958
rect 59826 13866 60026 14017
rect 61480 13866 86372 14177
rect 27387 13740 27474 13796
rect 27530 13740 27686 13796
rect 27742 13760 45977 13796
rect 50228 13790 86372 13866
rect 27742 13740 49775 13760
rect 27387 13578 49775 13740
rect 27387 13522 27474 13578
rect 27530 13522 27686 13578
rect 27742 13522 49775 13578
rect 27387 13361 49775 13522
rect 27387 13305 27474 13361
rect 27530 13305 27686 13361
rect 27742 13305 49775 13361
rect 27387 13245 49775 13305
rect 29478 13243 49775 13245
rect 24047 13031 27214 13193
rect 41493 13078 49775 13243
rect 50228 13734 57996 13790
rect 58052 13734 58208 13790
rect 58264 13734 86372 13790
rect 50228 13573 86372 13734
rect 50228 13517 57996 13573
rect 58052 13517 58208 13573
rect 58264 13517 86372 13573
rect 50228 13461 86372 13517
rect 50228 13355 58421 13461
rect 50228 13299 57996 13355
rect 58052 13299 58208 13355
rect 58264 13299 58421 13355
rect 50228 13138 58421 13299
rect 50228 13082 57996 13138
rect 58052 13082 58208 13138
rect 58264 13082 58421 13138
rect 24047 12975 26859 13031
rect 26915 12975 27071 13031
rect 27127 12975 27214 13031
rect 24047 12934 27214 12975
rect 24047 12847 34761 12934
rect 23821 12846 34761 12847
rect 0 12813 34761 12846
rect 0 12757 26859 12813
rect 26915 12757 27071 12813
rect 27127 12757 34761 12813
rect 0 12606 34761 12757
rect 50228 12920 58421 13082
rect 50228 12864 57996 12920
rect 58052 12864 58208 12920
rect 58264 12864 58421 12920
rect 50228 12846 58421 12864
rect 59826 12846 60026 13461
rect 83169 12846 84221 12847
rect 84666 12846 86372 13461
rect 50228 12702 86372 12846
rect 50228 12646 57996 12702
rect 58052 12646 58208 12702
rect 58264 12646 86372 12702
rect 50228 12606 86372 12646
rect 0 12596 86372 12606
rect 0 12540 26859 12596
rect 26915 12540 27071 12596
rect 27127 12540 86372 12596
rect 0 12484 86372 12540
rect 0 12428 57996 12484
rect 58052 12428 58208 12484
rect 58264 12428 86372 12484
rect 0 12378 86372 12428
rect 0 12322 26859 12378
rect 26915 12322 27071 12378
rect 27127 12322 86372 12378
rect 0 12267 86372 12322
rect 0 12211 57996 12267
rect 58052 12211 58208 12267
rect 58264 12211 86372 12267
rect 0 12161 86372 12211
rect 0 12105 26859 12161
rect 26915 12105 27071 12161
rect 27127 12105 86372 12161
rect 0 12049 86372 12105
rect 0 12046 57996 12049
rect 0 12036 24250 12046
rect 26772 11993 57996 12046
rect 58052 11993 58208 12049
rect 58264 12036 86372 12049
rect 58264 12035 84999 12036
rect 58264 11993 58351 12035
rect 26772 11844 58351 11993
rect 29478 11832 58351 11844
rect 29478 11776 57996 11832
rect 58052 11776 58208 11832
rect 58264 11776 58351 11832
rect 29478 11697 58351 11776
rect 0 11491 3011 11493
rect 24047 11491 27828 11493
rect 0 11406 27828 11491
rect 0 11350 27474 11406
rect 27530 11350 27686 11406
rect 27742 11350 27828 11406
rect 0 11189 27828 11350
rect 0 11133 27474 11189
rect 27530 11133 27686 11189
rect 27742 11133 27828 11189
rect 0 10971 27828 11133
rect 0 10915 27474 10971
rect 27530 10915 27686 10971
rect 27742 10915 27828 10971
rect 0 10753 27828 10915
rect 29478 10756 41516 11697
rect 0 10697 27474 10753
rect 27530 10697 27686 10753
rect 27742 10697 27828 10753
rect 0 10535 27828 10697
rect 0 10479 27474 10535
rect 27530 10479 27686 10535
rect 27742 10479 27828 10535
rect 0 10318 27828 10479
rect 0 10262 27474 10318
rect 27530 10262 27686 10318
rect 27742 10262 27828 10318
rect 0 10176 27828 10262
rect 2229 10175 24250 10176
rect 2249 10174 24250 10175
rect 23612 9942 29221 10030
rect 34741 9972 41516 10756
rect 42261 11491 57736 11527
rect 61825 11491 86372 11493
rect 42261 11406 86372 11491
rect 42261 11350 57381 11406
rect 57437 11350 57593 11406
rect 57649 11350 86372 11406
rect 42261 11189 86372 11350
rect 42261 11133 57381 11189
rect 57437 11133 57593 11189
rect 57649 11133 86372 11189
rect 42261 10971 86372 11133
rect 42261 10915 57381 10971
rect 57437 10915 57593 10971
rect 57649 10915 86372 10971
rect 42261 10753 86372 10915
rect 42261 10740 57381 10753
rect 57295 10697 57381 10740
rect 57437 10697 57593 10753
rect 57649 10697 86372 10753
rect 57295 10535 86372 10697
rect 57295 10479 57381 10535
rect 57437 10479 57593 10535
rect 57649 10479 86372 10535
rect 24047 9515 28729 9516
rect 0 9514 1014 9515
rect 2226 9514 28729 9515
rect 0 9407 28729 9514
rect 0 9351 26859 9407
rect 26915 9351 27071 9407
rect 27127 9351 28729 9407
rect 0 9190 28729 9351
rect 29133 9302 29221 9942
rect 41857 9502 51430 10420
rect 57295 10318 86372 10479
rect 57295 10262 57381 10318
rect 57437 10262 57593 10318
rect 57649 10262 86372 10318
rect 51750 10097 54952 10185
rect 57295 10176 86372 10262
rect 60736 10173 84482 10176
rect 51750 9971 51838 10097
rect 51750 9811 51766 9971
rect 51822 9811 51838 9971
rect 54864 10028 54952 10097
rect 54864 9940 65122 10028
rect 51750 9801 51838 9811
rect 58688 9681 66166 9777
rect 57909 9515 62278 9516
rect 57909 9514 72434 9515
rect 72602 9514 83234 9515
rect 85358 9514 86372 9515
rect 29133 9214 41656 9302
rect 0 9134 26859 9190
rect 26915 9134 27071 9190
rect 27127 9134 28729 9190
rect 0 8972 28729 9134
rect 0 8916 26859 8972
rect 26915 8916 27071 8972
rect 27127 8916 28729 8972
rect 0 8754 28729 8916
rect 41568 8972 41656 9214
rect 41857 9165 55482 9502
rect 41568 8953 50076 8972
rect 41568 8897 49906 8953
rect 50066 8897 50076 8953
rect 41568 8884 50076 8897
rect 50922 8965 55482 9165
rect 57909 9407 86372 9514
rect 57909 9351 57996 9407
rect 58052 9351 58208 9407
rect 58264 9351 86372 9407
rect 57909 9190 86372 9351
rect 57909 9134 57996 9190
rect 58052 9134 58208 9190
rect 58264 9134 86372 9190
rect 57909 8972 86372 9134
rect 0 8698 26859 8754
rect 26915 8698 27071 8754
rect 27127 8698 28729 8754
rect 0 8536 28729 8698
rect 50922 8854 57736 8965
rect 50922 8798 57381 8854
rect 57437 8798 57593 8854
rect 57649 8798 57736 8854
rect 50922 8636 57736 8798
rect 0 8480 26859 8536
rect 26915 8480 27071 8536
rect 27127 8480 28729 8536
rect 0 8319 28729 8480
rect 0 8263 26859 8319
rect 26915 8263 27071 8319
rect 27127 8263 28729 8319
rect 0 8154 28729 8263
rect 0 8153 24250 8154
rect 0 8152 3011 8153
rect 28178 7652 28729 8154
rect 29513 7900 41397 8582
rect 0 7595 3011 7596
rect 23625 7595 27828 7596
rect 0 7535 27828 7595
rect 0 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 0 7317 27828 7479
rect 0 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 0 7099 27828 7261
rect 0 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 28178 7084 34622 7652
rect 0 6982 27828 7043
rect 0 6199 1014 6982
rect 2226 6981 24250 6982
rect 2249 6980 24250 6981
rect 23625 6836 29058 6875
rect 23625 6780 28273 6836
rect 28329 6780 28484 6836
rect 28540 6780 28696 6836
rect 28752 6780 28907 6836
rect 28963 6780 29058 6836
rect 23625 6618 29058 6780
rect 29537 6744 34622 7084
rect 34860 7392 41397 7900
rect 50922 8580 57381 8636
rect 57437 8580 57593 8636
rect 57649 8580 57736 8636
rect 50922 8419 57736 8580
rect 50922 8363 57381 8419
rect 57437 8363 57593 8419
rect 57649 8363 57736 8419
rect 50922 8201 57736 8363
rect 50922 8145 57381 8201
rect 57437 8145 57593 8201
rect 57649 8145 57736 8201
rect 57909 8916 57996 8972
rect 58052 8916 58208 8972
rect 58264 8916 86372 8972
rect 57909 8754 86372 8916
rect 57909 8698 57996 8754
rect 58052 8698 58208 8754
rect 58264 8698 86372 8754
rect 57909 8536 86372 8698
rect 57909 8480 57996 8536
rect 58052 8480 58208 8536
rect 58264 8480 86372 8536
rect 57909 8319 86372 8480
rect 57909 8263 57996 8319
rect 58052 8263 58208 8319
rect 58264 8263 86372 8319
rect 57909 8154 86372 8263
rect 60736 8152 86372 8154
rect 50922 7983 57736 8145
rect 50922 7927 57381 7983
rect 57437 7927 57593 7983
rect 57649 7927 57736 7983
rect 50922 7766 57736 7927
rect 50922 7710 57381 7766
rect 57437 7710 57593 7766
rect 57649 7710 57736 7766
rect 50922 7596 57736 7710
rect 50922 7595 62747 7596
rect 83361 7595 86372 7596
rect 50922 7548 86372 7595
rect 50922 7492 57381 7548
rect 57437 7492 57593 7548
rect 57649 7492 86372 7548
rect 50922 7392 86372 7492
rect 34860 7330 86372 7392
rect 34860 7274 57381 7330
rect 57437 7274 57593 7330
rect 57649 7274 86372 7330
rect 34860 7113 86372 7274
rect 34860 7057 57381 7113
rect 57437 7057 57593 7113
rect 57649 7057 86372 7113
rect 34860 6984 86372 7057
rect 23625 6562 28273 6618
rect 28329 6562 28484 6618
rect 28540 6562 28696 6618
rect 28752 6562 28907 6618
rect 28963 6562 29058 6618
rect 34860 6592 55482 6984
rect 57295 6982 86372 6984
rect 60736 6980 84787 6982
rect 34860 6573 41397 6592
rect 23625 6400 29058 6562
rect 23625 6344 28273 6400
rect 28329 6344 28484 6400
rect 28540 6344 28696 6400
rect 28752 6344 28907 6400
rect 28963 6344 29058 6400
rect 23625 6306 29058 6344
rect 29458 6199 41397 6573
rect 0 6198 3011 6199
rect 23687 6198 41397 6199
rect 0 6177 41397 6198
rect 50922 6199 55482 6592
rect 56065 6836 62747 6875
rect 56065 6780 56160 6836
rect 56216 6780 56371 6836
rect 56427 6780 56583 6836
rect 56639 6780 56794 6836
rect 56850 6780 62747 6836
rect 56065 6618 62747 6780
rect 56065 6562 56160 6618
rect 56216 6562 56371 6618
rect 56427 6562 56583 6618
rect 56639 6562 56794 6618
rect 56850 6562 62747 6618
rect 56065 6400 62747 6562
rect 56065 6344 56160 6400
rect 56216 6344 56371 6400
rect 56427 6344 56583 6400
rect 56639 6344 56794 6400
rect 56850 6344 62747 6400
rect 56065 6306 62747 6344
rect 85358 6199 86372 6982
rect 50922 6198 62429 6199
rect 83361 6198 86372 6199
rect 0 6120 34622 6177
rect 0 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 34622 6120
rect 0 5902 34622 6064
rect 0 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 34622 5902
rect 0 5766 34622 5846
rect 29458 5665 34622 5766
rect 50922 6120 86372 6198
rect 50922 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 86372 6120
rect 50922 5902 86372 6064
rect 50922 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 86372 5902
rect 50922 5766 86372 5846
rect 23687 5629 27214 5630
rect 0 5539 27214 5629
rect 50922 5605 55482 5766
rect 57909 5629 62429 5630
rect 0 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27214 5539
rect 0 5321 27214 5483
rect 0 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27214 5321
rect 0 5175 27214 5265
rect 57909 5539 86372 5629
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 86372 5539
rect 57909 5462 86372 5483
rect 57909 5321 61287 5462
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5302 61287 5321
rect 61447 5302 86372 5462
rect 58264 5265 86372 5302
rect 57909 5175 86372 5265
rect 0 5174 24250 5175
rect 60736 5174 86372 5175
rect 0 5173 3011 5174
rect 83361 5173 86372 5174
rect 0 4515 1712 5173
rect 57909 4619 62429 4621
rect 23909 4528 62429 4619
rect 23909 4515 26859 4528
rect 0 4472 26859 4515
rect 26915 4472 27071 4528
rect 27127 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4515 62429 4528
rect 84660 4515 86372 5173
rect 58264 4472 86372 4515
rect 0 4310 86372 4472
rect 0 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 86372 4310
rect 0 4166 86372 4254
rect 0 4164 59323 4166
rect 0 4060 24341 4164
rect 60699 4060 86372 4166
rect 27438 3875 27778 3876
rect 28764 3875 28894 3876
rect 41774 3875 41904 3876
rect 42299 3875 42429 3876
rect 46873 3875 47003 3876
rect 47321 3875 47451 3876
rect 47769 3875 47899 3876
rect 48217 3875 48347 3876
rect 57345 3875 61215 3876
rect 23909 3837 61215 3875
rect 23909 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 28801 3837
rect 28857 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 61215 3837
rect 23909 3772 61215 3781
rect 0 3619 86372 3772
rect 0 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 28801 3619
rect 28857 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 86372 3619
rect 0 3524 86372 3563
rect 0 3421 24341 3524
rect 0 3420 3011 3421
rect 60699 3420 86372 3524
rect 0 2854 1014 3420
rect 24169 3044 62588 3066
rect 24169 2988 43800 3044
rect 43960 2988 62588 3044
rect 24169 2978 62588 2988
rect 85358 2854 86372 3420
rect 0 2502 86372 2854
rect 0 1232 86372 2232
rect 706 0 1706 1232
rect 2039 0 3039 1232
rect 3442 0 4442 1232
rect 4642 0 5642 932
rect 5842 0 6842 1232
rect 7042 0 8042 1232
rect 8242 0 9242 1232
rect 9442 0 10442 932
rect 10642 0 11642 1232
rect 12443 0 13443 1232
rect 14242 0 15242 1232
rect 15442 0 16442 932
rect 16642 0 17642 1232
rect 17842 0 18842 1232
rect 19042 0 20042 1232
rect 20242 0 21242 932
rect 21910 0 22910 1232
rect 23110 0 24110 1232
rect 24410 0 25410 1232
rect 25710 0 26710 1232
rect 27010 0 28010 1232
rect 28310 0 29310 1232
rect 29610 0 30610 1232
rect 31324 0 32324 932
rect 33022 0 34022 932
rect 34831 0 35831 932
rect 36031 0 37031 1232
rect 38028 0 39028 932
rect 39228 0 40228 1232
rect 41233 0 42233 932
rect 42433 0 43433 1232
rect 43633 0 44633 932
rect 44833 0 45833 1232
rect 46033 0 47033 932
rect 47233 0 48233 1232
rect 48566 0 49566 1232
rect 49876 0 50876 1232
rect 51233 0 52233 932
rect 52478 0 53478 932
rect 54458 0 55458 1232
rect 55758 0 56758 1232
rect 57058 0 58058 1232
rect 58358 0 59358 1232
rect 59658 0 60658 1232
rect 60958 0 61958 1232
rect 62295 0 63295 1232
rect 64218 0 65218 932
rect 65418 0 66418 1232
rect 66618 0 67618 1232
rect 67818 0 68818 1232
rect 69018 0 70018 932
rect 70218 0 71218 1232
rect 72017 0 73017 1232
rect 73818 0 74818 1232
rect 75018 0 76018 932
rect 76218 0 77218 1232
rect 77418 0 78418 1232
rect 78618 0 79618 1232
rect 79818 0 80818 932
rect 81018 0 82018 1232
rect 82419 0 83419 1232
rect 84666 0 85666 1232
use 256x8M8W_PWR_256x8m81  256x8M8W_PWR_256x8m81_0
timestamp 1749760379
transform 1 0 0 0 1 0
box 1912 6592 83548 35222
use control_512x8_256x8m81  control_512x8_256x8m81_0
timestamp 1749760379
transform 1 0 27533 0 1 4711
box -3624 -1833 31790 30125
use G_ring_256x8m81  G_ring_256x8m81_0
timestamp 1749760379
transform 1 0 282 0 1 0
box 0 0 85816 67902
use GF018_256x8M8WM1_lef_256x8m81  GF018_256x8M8WM1_lef_256x8m81_0
timestamp 1749760379
transform 1 0 0 0 1 0
box 0 0 86372 68176
use lcol4_256_256x8m81  lcol4_256_256x8m81_0
timestamp 1749760379
transform 1 0 2921 0 1 5019
box -1235 -3416 22164 60907
use M1_PSUB431059087816_256x8m81  M1_PSUB431059087816_256x8m81_0
timestamp 1749760379
transform 1 0 53710 0 1 2781
box 0 0 1 1
use M1_PSUB4310590878110_256x8m81  M1_PSUB4310590878110_256x8m81_0
timestamp 1749760379
transform 1 0 34404 0 1 2781
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_0
timestamp 1749760379
transform 1 0 28449 0 1 64027
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_1
timestamp 1749760379
transform 1 0 28449 0 1 62227
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_2
timestamp 1749760379
transform 1 0 28449 0 1 60427
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_3
timestamp 1749760379
transform 1 0 28449 0 1 58627
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_4
timestamp 1749760379
transform 1 0 28449 0 1 56827
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_5
timestamp 1749760379
transform 1 0 28449 0 1 55027
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_6
timestamp 1749760379
transform 1 0 28449 0 1 53227
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_7
timestamp 1749760379
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_8
timestamp 1749760379
transform 1 0 28449 0 1 49627
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_9
timestamp 1749760379
transform 1 0 28449 0 1 47827
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_10
timestamp 1749760379
transform 1 0 28449 0 1 46027
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_11
timestamp 1749760379
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_12
timestamp 1749760379
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_13
timestamp 1749760379
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_14
timestamp 1749760379
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_15
timestamp 1749760379
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_16
timestamp 1749760379
transform 1 0 28449 0 1 65827
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_17
timestamp 1749760379
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_18
timestamp 1749760379
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_19
timestamp 1749760379
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_20
timestamp 1749760379
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_21
timestamp 1749760379
transform 1 0 56674 0 1 46027
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_22
timestamp 1749760379
transform 1 0 56674 0 1 47827
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_23
timestamp 1749760379
transform 1 0 56674 0 1 49627
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_24
timestamp 1749760379
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_25
timestamp 1749760379
transform 1 0 56674 0 1 53227
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_26
timestamp 1749760379
transform 1 0 56674 0 1 55027
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_27
timestamp 1749760379
transform 1 0 56674 0 1 56827
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_28
timestamp 1749760379
transform 1 0 56674 0 1 58627
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_29
timestamp 1749760379
transform 1 0 56674 0 1 60427
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_30
timestamp 1749760379
transform 1 0 56674 0 1 62227
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_31
timestamp 1749760379
transform 1 0 56674 0 1 64027
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_32
timestamp 1749760379
transform 1 0 56674 0 1 65827
box 0 0 1 1
use M2_M1$$199747628_256x8m81  M2_M1$$199747628_256x8m81_33
timestamp 1749760379
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M2_M1$$201260076_256x8m81  M2_M1$$201260076_256x8m81_0
timestamp 1749760379
transform -1 0 57515 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_256x8m81  M2_M1$$201260076_256x8m81_1
timestamp 1749760379
transform -1 0 58130 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_256x8m81  M2_M1$$201260076_256x8m81_2
timestamp 1749760379
transform 1 0 27608 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_256x8m81  M2_M1$$201260076_256x8m81_3
timestamp 1749760379
transform 1 0 26993 0 1 19369
box 0 0 1 1
use M2_M1$$201261100_256x8m81  M2_M1$$201261100_256x8m81_0
timestamp 1749760379
transform -1 0 58130 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_256x8m81  M2_M1$$201261100_256x8m81_1
timestamp 1749760379
transform -1 0 57515 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_256x8m81  M2_M1$$201261100_256x8m81_2
timestamp 1749760379
transform 1 0 27608 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_256x8m81  M2_M1$$201261100_256x8m81_3
timestamp 1749760379
transform 1 0 26993 0 1 4126
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_0
timestamp 1749760379
transform 1 0 62227 0 1 1663
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_1
timestamp 1749760379
transform 1 0 72743 0 1 1663
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_2
timestamp 1749760379
transform 1 0 72293 0 1 1663
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_3
timestamp 1749760379
transform 1 0 82808 0 1 1663
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_4
timestamp 1749760379
transform 1 0 51732 0 1 5173
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_5
timestamp 1749760379
transform 1 0 49986 0 1 6323
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_6
timestamp 1749760379
transform 1 0 23517 0 1 1663
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_7
timestamp 1749760379
transform 1 0 13167 0 1 1663
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_8
timestamp 1749760379
transform 1 0 12717 0 1 1663
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_9
timestamp 1749760379
transform 1 0 2652 0 1 1663
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_10
timestamp 1749760379
transform 1 0 40701 0 1 3256
box 0 0 1 1
use M2_M1431059087813_256x8m81  M2_M1431059087813_256x8m81_0
timestamp 1749760379
transform 1 0 27599 0 1 34778
box 0 0 1 1
use M2_M1431059087817_256x8m81  M2_M1431059087817_256x8m81_0
timestamp 1749760379
transform 1 0 25654 0 1 65826
box 0 0 1 1
use M2_M1431059087817_256x8m81  M2_M1431059087817_256x8m81_1
timestamp 1749760379
transform 1 0 59132 0 1 65826
box 0 0 1 1
use M2_M1431059087818_256x8m81  M2_M1431059087818_256x8m81_0
timestamp 1749760379
transform 1 0 25682 0 1 34809
box 0 0 1 1
use M2_M1431059087818_256x8m81  M2_M1431059087818_256x8m81_1
timestamp 1749760379
transform 1 0 59160 0 1 34829
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_0
timestamp 1749760379
transform 1 0 29118 0 1 787
box 0 0 1 1
use M2_M14310590878112_256x8m81  M2_M14310590878112_256x8m81_0
timestamp 1749760379
transform 1 0 61367 0 1 5401
box 0 0 1 1
use m2m3_256x8m81  m2m3_256x8m81_0
timestamp 1749760379
transform 1 0 58611 0 1 17122
box 0 0 3541 9202
use M3_M2$$201248812_256x8m81  M3_M2$$201248812_256x8m81_0
timestamp 1749760379
transform -1 0 58130 0 1 12783
box 0 0 1 1
use M3_M2$$201248812_256x8m81  M3_M2$$201248812_256x8m81_1
timestamp 1749760379
transform -1 0 57515 0 1 15671
box 0 0 1 1
use M3_M2$$201248812_256x8m81  M3_M2$$201248812_256x8m81_2
timestamp 1749760379
transform 1 0 27608 0 1 15463
box 0 0 1 1
use M3_M2$$201248812_256x8m81  M3_M2$$201248812_256x8m81_3
timestamp 1749760379
transform 1 0 26993 0 1 13112
box 0 0 1 1
use M3_M2$$201249836_256x8m81  M3_M2$$201249836_256x8m81_0
timestamp 1749760379
transform -1 0 57515 0 1 10834
box 0 0 1 1
use M3_M2$$201249836_256x8m81  M3_M2$$201249836_256x8m81_1
timestamp 1749760379
transform -1 0 58130 0 1 8835
box 0 0 1 1
use M3_M2$$201249836_256x8m81  M3_M2$$201249836_256x8m81_2
timestamp 1749760379
transform 1 0 27608 0 1 10834
box 0 0 1 1
use M3_M2$$201249836_256x8m81  M3_M2$$201249836_256x8m81_3
timestamp 1749760379
transform 1 0 26993 0 1 8835
box 0 0 1 1
use M3_M2$$201250860_256x8m81  M3_M2$$201250860_256x8m81_0
timestamp 1749760379
transform -1 0 56505 0 1 6590
box 0 0 1 1
use M3_M2$$201250860_256x8m81  M3_M2$$201250860_256x8m81_1
timestamp 1749760379
transform 1 0 28618 0 1 6590
box 0 0 1 1
use M3_M2$$201251884_256x8m81  M3_M2$$201251884_256x8m81_0
timestamp 1749760379
transform 1 0 37303 0 1 35853
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_0
timestamp 1749760379
transform 1 0 28829 0 1 3700
box 0 0 1 1
use M3_M2$$201253932_256x8m81  M3_M2$$201253932_256x8m81_0
timestamp 1749760379
transform 1 0 57515 0 1 8173
box 0 0 1 1
use M3_M2$$201254956_256x8m81  M3_M2$$201254956_256x8m81_0
timestamp 1749760379
transform 1 0 27608 0 1 13768
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_0
timestamp 1749760379
transform 1 0 28449 0 1 62227
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_1
timestamp 1749760379
transform 1 0 28449 0 1 60427
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_2
timestamp 1749760379
transform 1 0 28449 0 1 58627
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_3
timestamp 1749760379
transform 1 0 28449 0 1 56827
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_4
timestamp 1749760379
transform 1 0 28449 0 1 55027
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_5
timestamp 1749760379
transform 1 0 28449 0 1 53227
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_6
timestamp 1749760379
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_7
timestamp 1749760379
transform 1 0 28449 0 1 49627
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_8
timestamp 1749760379
transform 1 0 28449 0 1 47827
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_9
timestamp 1749760379
transform 1 0 28449 0 1 46027
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_10
timestamp 1749760379
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_11
timestamp 1749760379
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_12
timestamp 1749760379
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_13
timestamp 1749760379
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_14
timestamp 1749760379
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_15
timestamp 1749760379
transform 1 0 28449 0 1 65827
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_16
timestamp 1749760379
transform 1 0 28449 0 1 64027
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_17
timestamp 1749760379
transform 1 0 56674 0 1 62227
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_18
timestamp 1749760379
transform 1 0 56674 0 1 64027
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_19
timestamp 1749760379
transform 1 0 56674 0 1 65827
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_20
timestamp 1749760379
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_21
timestamp 1749760379
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_22
timestamp 1749760379
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_23
timestamp 1749760379
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_24
timestamp 1749760379
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_25
timestamp 1749760379
transform 1 0 56674 0 1 46027
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_26
timestamp 1749760379
transform 1 0 56674 0 1 47827
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_27
timestamp 1749760379
transform 1 0 56674 0 1 49627
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_28
timestamp 1749760379
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_29
timestamp 1749760379
transform 1 0 56674 0 1 53227
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_30
timestamp 1749760379
transform 1 0 56674 0 1 55027
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_31
timestamp 1749760379
transform 1 0 56674 0 1 56827
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_32
timestamp 1749760379
transform 1 0 56674 0 1 58627
box 0 0 1 1
use M3_M2$$201258028_256x8m81  M3_M2$$201258028_256x8m81_33
timestamp 1749760379
transform 1 0 56674 0 1 60427
box 0 0 1 1
use M3_M2$$201412652_256x8m81  M3_M2$$201412652_256x8m81_0
timestamp 1749760379
transform -1 0 57515 0 1 30897
box 0 0 1 1
use M3_M2$$201412652_256x8m81  M3_M2$$201412652_256x8m81_1
timestamp 1749760379
transform -1 0 57515 0 1 32786
box 0 0 1 1
use M3_M2$$201412652_256x8m81  M3_M2$$201412652_256x8m81_2
timestamp 1749760379
transform 1 0 27608 0 1 32786
box 0 0 1 1
use M3_M2$$201412652_256x8m81  M3_M2$$201412652_256x8m81_3
timestamp 1749760379
transform 1 0 27608 0 1 30897
box 0 0 1 1
use M3_M2$$201413676_256x8m81  M3_M2$$201413676_256x8m81_0
timestamp 1749760379
transform -1 0 58130 0 1 31842
box 0 0 1 1
use M3_M2$$201413676_256x8m81  M3_M2$$201413676_256x8m81_1
timestamp 1749760379
transform 1 0 27608 0 1 7289
box 0 0 1 1
use M3_M2$$201413676_256x8m81  M3_M2$$201413676_256x8m81_2
timestamp 1749760379
transform 1 0 26993 0 1 31842
box 0 0 1 1
use M3_M2$$201413676_256x8m81  M3_M2$$201413676_256x8m81_3
timestamp 1749760379
transform 1 0 27612 0 1 34778
box 0 0 1 1
use M3_M2$$201414700_256x8m81  M3_M2$$201414700_256x8m81_0
timestamp 1749760379
transform -1 0 58130 0 1 33221
box 0 0 1 1
use M3_M2$$201414700_256x8m81  M3_M2$$201414700_256x8m81_1
timestamp 1749760379
transform 1 0 26993 0 1 33221
box 0 0 1 1
use M3_M2$$201415724_256x8m81  M3_M2$$201415724_256x8m81_0
timestamp 1749760379
transform -1 0 58130 0 1 28743
box 0 0 1 1
use M3_M2$$201415724_256x8m81  M3_M2$$201415724_256x8m81_1
timestamp 1749760379
transform 1 0 26993 0 1 28743
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_0
timestamp 1749760379
transform -1 0 57515 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_1
timestamp 1749760379
transform -1 0 57515 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_2
timestamp 1749760379
transform -1 0 58130 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_3
timestamp 1749760379
transform -1 0 57515 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_4
timestamp 1749760379
transform -1 0 58130 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_5
timestamp 1749760379
transform 1 0 27608 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_6
timestamp 1749760379
transform 1 0 26993 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_7
timestamp 1749760379
transform 1 0 27608 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_8
timestamp 1749760379
transform 1 0 26993 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_9
timestamp 1749760379
transform 1 0 27608 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_10
timestamp 1749760379
transform 1 0 27608 0 1 24891
box 0 0 1 1
use M3_M2431059087811_256x8m81  M3_M2431059087811_256x8m81_0
timestamp 1749760379
transform 0 -1 49986 1 0 8925
box 0 0 1 1
use M3_M2431059087811_256x8m81  M3_M2431059087811_256x8m81_1
timestamp 1749760379
transform 1 0 51794 0 1 9891
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_0
timestamp 1749760379
transform 1 0 58128 0 1 20490
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_1
timestamp 1749760379
transform 1 0 58128 0 1 20146
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_2
timestamp 1749760379
transform 1 0 61367 0 1 5382
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_3
timestamp 1749760379
transform 1 0 26187 0 1 19267
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_4
timestamp 1749760379
transform 1 0 26530 0 1 26206
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_5
timestamp 1749760379
transform 1 0 26545 0 1 19612
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_6
timestamp 1749760379
transform 1 0 27004 0 1 20490
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_7
timestamp 1749760379
transform 1 0 27004 0 1 20146
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_8
timestamp 1749760379
transform 1 0 24137 0 1 23593
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_9
timestamp 1749760379
transform 1 0 24149 0 1 17237
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_10
timestamp 1749760379
transform 1 0 24496 0 1 23915
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_11
timestamp 1749760379
transform 1 0 24509 0 1 17576
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_12
timestamp 1749760379
transform 1 0 24824 0 1 24236
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_13
timestamp 1749760379
transform 1 0 24837 0 1 17897
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_14
timestamp 1749760379
transform 1 0 25161 0 1 24557
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_15
timestamp 1749760379
transform 1 0 25174 0 1 18270
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_16
timestamp 1749760379
transform 1 0 25501 0 1 25248
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_17
timestamp 1749760379
transform 1 0 25514 0 1 18604
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_18
timestamp 1749760379
transform 1 0 25836 0 1 25567
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_19
timestamp 1749760379
transform 1 0 25851 0 1 18947
box 0 0 1 1
use M3_M2431059087812_256x8m81  M3_M2431059087812_256x8m81_20
timestamp 1749760379
transform 1 0 26172 0 1 25887
box 0 0 1 1
use M3_M2431059087814_256x8m81  M3_M2431059087814_256x8m81_0
timestamp 1749760379
transform 1 0 43880 0 1 3016
box 0 0 1 1
use M3_M2431059087814_256x8m81  M3_M2431059087814_256x8m81_1
timestamp 1749760379
transform 1 0 41961 0 1 64926
box 0 0 1 1
use M3_M2431059087815_256x8m81  M3_M2431059087815_256x8m81_0
timestamp 1749760379
transform 1 0 59149 0 1 31146
box 0 0 1 1
use M3_M2431059087815_256x8m81  M3_M2431059087815_256x8m81_1
timestamp 1749760379
transform 1 0 59149 0 1 30701
box 0 0 1 1
use M3_M2431059087815_256x8m81  M3_M2431059087815_256x8m81_2
timestamp 1749760379
transform 1 0 25674 0 1 30641
box 0 0 1 1
use M3_M2431059087815_256x8m81  M3_M2431059087815_256x8m81_3
timestamp 1749760379
transform 1 0 25674 0 1 31096
box 0 0 1 1
use M3_M2431059087819_256x8m81  M3_M2431059087819_256x8m81_0
timestamp 1749760379
transform 1 0 58126 0 1 23631
box 0 0 1 1
use M3_M2431059087819_256x8m81  M3_M2431059087819_256x8m81_1
timestamp 1749760379
transform 1 0 57495 0 1 22479
box 0 0 1 1
use M3_M2431059087819_256x8m81  M3_M2431059087819_256x8m81_2
timestamp 1749760379
transform 1 0 26990 0 1 23631
box 0 0 1 1
use M3_M2431059087819_256x8m81  M3_M2431059087819_256x8m81_3
timestamp 1749760379
transform 1 0 27607 0 1 22492
box 0 0 1 1
use M3_M24310590878113_256x8m81  M3_M24310590878113_256x8m81_0
timestamp 1749760379
transform 1 0 59135 0 1 27425
box 0 0 1 1
use M3_M24310590878113_256x8m81  M3_M24310590878113_256x8m81_1
timestamp 1749760379
transform 1 0 25680 0 1 27419
box 0 0 1 1
use M3_M24310590878114_256x8m81  M3_M24310590878114_256x8m81_0
timestamp 1749760379
transform 1 0 25682 0 1 34809
box 0 0 1 1
use M3_M24310590878114_256x8m81  M3_M24310590878114_256x8m81_1
timestamp 1749760379
transform 1 0 59160 0 1 34829
box 0 0 1 1
use M3_M24310590878115_256x8m81  M3_M24310590878115_256x8m81_0
timestamp 1749760379
transform 1 0 25654 0 1 65826
box 0 0 1 1
use M3_M24310590878115_256x8m81  M3_M24310590878115_256x8m81_1
timestamp 1749760379
transform 1 0 59132 0 1 65826
box 0 0 1 1
use power_a_256x8m81  power_a_256x8m81_0
timestamp 1749760379
transform -1 0 80818 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_1
timestamp 1749760379
transform -1 0 70018 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_2
timestamp 1749760379
transform 1 0 64218 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_3
timestamp 1749760379
transform 1 0 52478 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_4
timestamp 1749760379
transform 1 0 46033 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_5
timestamp 1749760379
transform 1 0 43633 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_6
timestamp 1749760379
transform 1 0 51233 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_7
timestamp 1749760379
transform 1 0 75018 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_8
timestamp 1749760379
transform -1 0 32324 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_9
timestamp 1749760379
transform -1 0 21242 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_10
timestamp 1749760379
transform -1 0 10442 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_11
timestamp 1749760379
transform -1 0 34022 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_12
timestamp 1749760379
transform 1 0 41233 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_13
timestamp 1749760379
transform 1 0 38028 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_14
timestamp 1749760379
transform 1 0 34831 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_15
timestamp 1749760379
transform 1 0 15442 0 1 282
box 0 -282 1000 1000
use power_a_256x8m81  power_a_256x8m81_16
timestamp 1749760379
transform 1 0 4642 0 1 282
box 0 -282 1000 1000
use power_route_01_a_256x8m81  power_route_01_a_256x8m81_0
timestamp 1749760379
transform 1 0 4648 0 1 65746
box -511 630 1714 2430
use power_route_01_a_256x8m81  power_route_01_a_256x8m81_1
timestamp 1749760379
transform 1 0 10048 0 1 65746
box -511 630 1714 2430
use power_route_01_a_256x8m81  power_route_01_a_256x8m81_2
timestamp 1749760379
transform 1 0 15448 0 1 65746
box -511 630 1714 2430
use power_route_01_a_256x8m81  power_route_01_a_256x8m81_3
timestamp 1749760379
transform 1 0 69624 0 1 65746
box -511 630 1714 2430
use power_route_01_a_256x8m81  power_route_01_a_256x8m81_4
timestamp 1749760379
transform 1 0 64224 0 1 65746
box -511 630 1714 2430
use power_route_01_a_256x8m81  power_route_01_a_256x8m81_5
timestamp 1749760379
transform 1 0 46824 0 1 65746
box -511 630 1714 2430
use power_route_01_a_256x8m81  power_route_01_a_256x8m81_6
timestamp 1749760379
transform 1 0 75024 0 1 65746
box -511 630 1714 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_0
timestamp 1749760379
transform -1 0 31199 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_1
timestamp 1749760379
transform -1 0 35904 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_2
timestamp 1749760379
transform -1 0 39074 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_3
timestamp 1749760379
transform -1 0 41719 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_4
timestamp 1749760379
transform -1 0 21142 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_5
timestamp 1749760379
transform -1 0 27061 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_6
timestamp 1749760379
transform -1 0 83548 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_7
timestamp 1749760379
transform -1 0 85155 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_8
timestamp 1749760379
transform -1 0 80718 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_9
timestamp 1749760379
transform -1 0 53058 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_10
timestamp 1749760379
transform -1 0 54751 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_11
timestamp 1749760379
transform -1 0 49390 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_12
timestamp 1749760379
transform -1 0 58036 0 1 65746
box -511 630 489 2430
use power_route_01_b_256x8m81  power_route_01_b_256x8m81_13
timestamp 1749760379
transform -1 0 45558 0 1 65746
box -511 630 489 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_0
timestamp 1749760379
transform -1 0 35738 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_1
timestamp 1749760379
transform -1 0 38662 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_2
timestamp 1749760379
transform -1 0 41596 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_3
timestamp 1749760379
transform -1 0 26872 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_4
timestamp 1749760379
transform -1 0 29591 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_5
timestamp 1749760379
transform -1 0 30987 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_6
timestamp 1749760379
transform -1 0 34095 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_7
timestamp 1749760379
transform -1 0 45427 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_8
timestamp 1749760379
transform -1 0 83548 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_9
timestamp 1749760379
transform -1 0 52179 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_10
timestamp 1749760379
transform -1 0 57704 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_11
timestamp 1749760379
transform -1 0 60505 0 1 65746
box 714 1822 1714 2430
use power_route_01_c_256x8m81  power_route_01_c_256x8m81_12
timestamp 1749760379
transform -1 0 44144 0 1 65746
box 714 1822 1714 2430
use power_route_256_256x8m81  power_route_256_256x8m81_0
timestamp 1749760379
transform 1 0 -1921 0 1 -2063
box 1921 2345 88293 70239
use rcol4_256_256x8m81  rcol4_256_256x8m81_0
timestamp 1749760379
transform 1 0 60511 0 1 5019
box -493 -3398 24936 60907
use xdec32_256_256x8m81  xdec32_256_256x8m81_0
timestamp 1749760379
transform 1 0 28677 0 1 36127
box 155 -1 27614 29760
<< labels >>
flabel metal3 s 2626 67568 3626 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 64576 1706 65276 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 4642 0 5642 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 5362 67568 6362 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 62776 1706 63476 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 60976 1706 61676 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 59176 1706 59876 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 8026 67568 9026 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 9442 0 10442 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 10762 67568 11762 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 13426 67568 14426 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 57376 1706 58076 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 55576 1706 56276 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 53776 1706 54476 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 51976 1706 52676 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 50176 1706 50876 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 48376 1706 49076 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 46576 1706 47276 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 44776 1706 45476 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 15442 0 16442 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 16162 67568 17162 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 18826 67568 19826 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 20242 0 21242 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 22258 67568 23258 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 25158 67568 26158 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 26435 26070 28416 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 42976 1706 43676 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 41176 1706 41876 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 39376 1706 40076 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 1954 26435 26070 28434 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 26435 27828 26890 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 10176 3011 11493 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 2249 10174 24250 11491 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 2229 10175 24250 11491 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 24047 10176 27828 11493 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 34536 1014 35326 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 35126 24917 35326 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 37576 1706 38276 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 35776 1706 36476 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 8152 1014 9515 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 8152 3011 9514 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 2226 8154 28729 9515 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 8153 24250 9514 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 28178 7084 28729 9516 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 24047 8154 28729 9516 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 29537 6744 34622 7652 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 27442 34494 27782 35062 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 28178 7084 34622 7652 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 34536 27830 35016 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 1401 66376 2401 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 27877 67568 28877 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 4137 66376 5137 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 6801 66376 7801 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 29273 67568 30273 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 9537 66376 10537 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 31324 0 32324 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 12201 66376 13201 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 32381 67568 33381 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 14937 66376 15937 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 17601 66376 18601 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 33022 0 34022 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 34024 67568 35024 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 20653 66376 21653 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 34831 0 35831 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 23483 66376 24483 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 36948 67568 37948 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 38028 0 39028 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 39882 67568 40882 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 41233 0 42233 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 42430 67568 43430 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 43633 0 44633 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 43713 67568 44713 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 46033 0 47033 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 47538 67568 48538 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 26572 66376 27572 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 50465 67568 51465 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 30710 66376 31710 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 51233 0 52233 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 35415 66376 36415 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 38585 66376 39585 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 41230 66376 42230 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 45069 66376 46069 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 46313 66376 47313 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 48901 66376 49901 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 52569 66376 53569 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 54262 66376 55262 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 52478 0 53478 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 55990 67568 56990 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 58791 67568 59791 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 62202 67568 63202 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 64218 0 65218 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 64938 67568 65938 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 67602 67568 68603 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 69018 0 70018 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 57547 66376 58547 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 70338 67568 71338 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 60977 66376 61977 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 73002 67568 74002 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 63713 66376 64713 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 75018 0 76018 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 66378 66376 67378 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 75738 67568 76738 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 66377 67568 67378 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 69113 66376 70113 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 71777 66376 72777 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 74513 66376 75513 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 77177 66376 78177 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 80229 66376 81229 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 83059 66376 84059 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 84666 66376 85666 68176 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 66376 86372 67376 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 84666 64576 86372 65276 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 78402 67568 79402 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 62776 86372 63476 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 79818 0 80818 932 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 60976 86372 61676 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 81834 67568 82834 68176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 59176 86372 59876 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 65476 1014 66176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 57376 86372 58076 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 65676 27272 65976 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 55576 86372 56276 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 65726 27779 65928 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 53776 86372 54476 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 30402 65726 54622 65928 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 65727 57494 65928 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 51976 86372 52676 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 57410 65726 86372 65926 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 60471 65676 86372 65976 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 50176 86372 50876 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 85358 65476 86372 66176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 63676 1014 64376 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 48376 86372 49076 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 84666 46576 86372 47276 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 84666 44776 86372 45476 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 84666 42976 86372 43676 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 84666 41176 86372 41876 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 84666 39376 86372 40076 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 84666 37576 86372 38276 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 84666 35776 86372 36476 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 29430 1706 34125 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 63876 27272 64176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 2095 32315 2188 34126 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 30403 63926 54622 64128 0 FreeSans 448 180 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 63927 86372 64128 0 FreeSans 448 180 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 32315 3011 34125 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 32316 25085 34125 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 32318 27214 34124 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 26772 31486 58351 32199 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 26772 27382 58351 30105 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 60471 63876 86372 64176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 57908 31486 58351 34124 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 61853 32315 72383 34125 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 57908 32315 86372 34124 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 85358 63676 86372 64376 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 29430 86372 29714 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 61876 1014 62576 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 29430 86372 34125 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 62076 27272 62376 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 72653 32315 86372 34125 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 30403 62126 54622 62328 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 22938 1706 23938 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 62127 86372 62328 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 22938 27214 23380 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 60471 62076 86372 62376 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 26770 23370 58348 24278 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 57908 22937 83763 23380 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 57908 22938 86372 23380 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 84666 22938 86372 23938 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 18016 24250 20739 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 85358 61876 86372 62576 0 FreeSans 448 180 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 60076 1014 60776 0 FreeSans 448 180 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 60276 27272 60576 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 30403 60326 54622 60528 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 60327 86372 60528 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 29513 19969 55645 21625 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 29521 19969 55645 21707 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 44432 19969 55645 21708 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 61502 18015 83763 20739 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 60471 60276 86372 60576 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 61502 18016 86372 20739 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 19969 86372 20739 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 12036 1706 14178 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 23821 12046 34761 12847 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 13461 27214 14178 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 85358 60076 86372 60776 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 58276 1014 58976 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 12036 24250 12846 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 24047 12046 27214 14179 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 24047 12046 34761 12934 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 58476 27272 58776 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 34741 9972 41516 12606 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 29478 10756 41516 12606 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 29478 11697 58351 12606 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 26772 11844 58351 12606 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 30403 58526 54622 58728 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 50228 12035 58421 13866 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 59826 12035 60026 14017 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 58527 86372 58728 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 60471 58476 86372 58776 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 85358 58276 86372 58976 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 0 56476 1014 57176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 50228 13461 86372 13866 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 61807 13461 72429 14178 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 61480 13461 86372 14177 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 83169 12035 84221 12847 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 83169 13461 84221 14179 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 50228 12036 86372 12846 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 56676 27272 56976 0 FreeSans 448 180 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 30403 56726 54622 56928 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 26772 12035 84999 12606 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 0 56727 86372 56928 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 60471 56676 86372 56976 0 FreeSans 448 180 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 85358 56476 86372 57176 0 FreeSans 448 0 0 0 VSS
port 29 nsew ground bidirectional
flabel metal3 s 84666 12036 86372 14178 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 72607 13461 86372 14178 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 57909 8154 62278 9516 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 57909 8154 72434 9515 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 72602 8152 83234 9515 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 60736 8152 86372 9514 0 FreeSans 448 180 0 0 VDD
port 28 nsew power bidirectional
flabel metal3 s 85358 8152 86372 9515 0 FreeSans 448 0 0 0 VDD
port 28 nsew power bidirectional
flabel metal2 s 27936 0 28160 200 0 FreeSans 1600 0 0 0 CLK
port 10 nsew signal input
flabel metal2 s 1864 0 2088 200 0 FreeSans 1000 0 0 0 D[0]
port 18 nsew signal input
flabel metal2 s 29705 0 29929 200 0 FreeSans 1600 0 0 0 A[7]
port 1 nsew signal input
flabel metal2 s 30859 0 31083 200 0 FreeSans 1600 0 0 0 A[2]
port 6 nsew signal input
flabel metal2 s 32552 0 32776 200 0 FreeSans 1600 0 0 0 A[1]
port 7 nsew signal input
flabel metal2 s 34243 0 34467 200 0 FreeSans 1600 0 0 0 A[0]
port 8 nsew signal input
flabel metal2 s 14127 0 14351 200 0 FreeSans 1000 180 0 0 Q[2]
port 25 nsew signal output
flabel metal2 s 22279 0 22503 200 0 FreeSans 1000 180 0 0 Q[3]
port 24 nsew signal output
flabel metal2 s 50342 0 50566 200 0 FreeSans 1600 0 0 0 CEN
port 9 nsew signal input
flabel metal2 s 54417 0 54641 200 0 FreeSans 1600 0 0 0 A[5]
port 3 nsew signal input
flabel metal2 s 53772 0 53996 200 0 FreeSans 1600 0 0 0 A[6]
port 2 nsew signal input
flabel metal2 s 55164 0 55388 200 0 FreeSans 1600 0 0 0 A[4]
port 4 nsew signal input
flabel metal2 s 23404 0 23628 200 0 FreeSans 1000 180 0 0 WEN[3]
port 34 nsew signal input
flabel metal2 s 23795 0 24019 200 0 FreeSans 1000 180 0 0 D[3]
port 15 nsew signal input
flabel metal2 s 12206 0 12430 200 0 FreeSans 1000 180 0 0 D[1]
port 17 nsew signal input
flabel metal2 s 13454 0 13678 200 0 FreeSans 1000 180 0 0 D[2]
port 16 nsew signal input
flabel metal2 s 56265 0 56489 200 0 FreeSans 1600 0 0 0 A[3]
port 5 nsew signal input
flabel metal2 s 11533 0 11757 200 0 FreeSans 1000 180 0 0 Q[1]
port 26 nsew signal output
flabel metal2 s 73703 0 73927 200 0 FreeSans 1000 180 0 0 Q[6]
port 21 nsew signal output
flabel metal2 s 71782 0 72006 200 0 FreeSans 1000 180 0 0 D[5]
port 13 nsew signal input
flabel metal2 s 62958 0 63182 200 0 FreeSans 1000 180 0 0 Q[4]
port 23 nsew signal output
flabel metal2 s 72180 0 72404 200 0 FreeSans 1000 180 0 0 WEN[5]
port 32 nsew signal input
flabel metal2 s 13054 0 13278 200 0 FreeSans 1000 180 0 0 WEN[2]
port 35 nsew signal input
flabel metal2 s 12604 0 12828 200 0 FreeSans 1000 180 0 0 WEN[1]
port 36 nsew signal input
flabel metal2 s 62115 0 62339 200 0 FreeSans 1000 180 0 0 WEN[4]
port 33 nsew signal input
flabel metal2 s 82695 0 82919 200 0 FreeSans 1000 180 0 0 WEN[7]
port 30 nsew signal input
flabel metal2 s 72630 0 72854 200 0 FreeSans 1000 180 0 0 WEN[6]
port 31 nsew signal input
flabel metal2 s 73030 0 73254 200 0 FreeSans 1000 180 0 0 D[6]
port 12 nsew signal input
flabel metal2 s 71109 0 71333 200 0 FreeSans 1000 180 0 0 Q[5]
port 22 nsew signal output
flabel metal2 s 3380 0 3604 200 0 FreeSans 1000 0 0 0 Q[0]
port 27 nsew signal output
flabel metal2 s 40588 0 40812 200 0 FreeSans 1600 0 0 0 GWEN
port 19 nsew signal input
flabel metal2 s 2539 0 2763 200 0 FreeSans 1000 0 0 0 WEN[0]
port 37 nsew signal input
flabel metal2 s 61447 0 61671 200 0 FreeSans 1000 180 0 0 D[4]
port 14 nsew signal input
flabel metal2 s 83372 0 83596 200 0 FreeSans 1000 180 0 0 D[7]
port 11 nsew signal input
flabel metal2 s 81855 0 82079 200 0 FreeSans 1000 180 0 0 Q[7]
port 20 nsew signal output
rlabel metal3 s 0 4060 1712 5629 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 5173 3011 5629 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 5174 24250 5629 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 4060 24341 4515 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 23687 5175 27214 5630 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 23909 4166 62429 4619 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 4164 59323 4515 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 57909 4166 62429 4621 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 57909 5175 62429 5630 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 60699 4060 86372 4515 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 83361 5173 86372 5629 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 60736 5174 86372 5629 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 84660 4060 86372 5629 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 706 0 1706 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 2039 0 3039 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 3442 0 4442 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 5842 0 6842 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 7042 0 8042 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 8242 0 9242 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 10642 0 11642 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 12443 0 13443 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 14242 0 15242 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 16642 0 17642 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 17842 0 18842 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 19042 0 20042 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 21910 0 22910 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 23110 0 24110 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 24410 0 25410 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 25710 0 26710 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 27010 0 28010 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 28310 0 29310 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 29610 0 30610 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 36031 0 37031 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 39228 0 40228 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 42433 0 43433 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 44833 0 45833 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 47233 0 48233 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 48566 0 49566 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 49876 0 50876 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 54458 0 55458 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 55758 0 56758 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 57058 0 58058 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 58358 0 59358 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 59658 0 60658 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 60958 0 61958 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 62295 0 63295 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 65418 0 66418 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 66618 0 67618 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 67818 0 68818 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 70218 0 71218 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 72017 0 73017 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 73818 0 74818 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 76218 0 77218 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 77418 0 78418 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 78618 0 79618 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 81018 0 82018 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 82419 0 83419 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 84666 0 85666 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 1232 86372 2232 1 VDD
port 28 nsew power bidirectional
rlabel metal3 s 0 54676 1014 55376 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 54876 27272 55176 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 54926 54622 55128 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 54927 86372 55128 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 54876 86372 55176 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 54676 86372 55376 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 52876 1014 53576 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 53076 27272 53376 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 53126 54622 53328 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 53127 86372 53328 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 53076 86372 53376 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 52876 86372 53576 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 51076 1014 51776 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 51276 27272 51576 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 51326 54622 51528 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 51327 86372 51528 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 51276 86372 51576 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 51076 86372 51776 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 49276 1014 49976 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 49476 27272 49776 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 49526 54622 49728 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 49527 86372 49728 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 49476 86372 49776 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 49276 86372 49976 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 47476 1014 48176 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 47676 27272 47976 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 47726 54622 47928 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 47727 86372 47928 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 47676 86372 47976 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 47476 86372 48176 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 45676 1014 46376 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 45876 27272 46176 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 45926 54622 46128 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 45927 86372 46128 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 45876 86372 46176 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 45676 86372 46376 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 43876 1014 44576 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 44076 27272 44376 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 44126 54622 44328 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 44127 86372 44328 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 44076 86372 44376 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 43876 86372 44576 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 42076 1014 42776 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 42276 27272 42576 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 42326 54622 42528 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 42327 86372 42528 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 42276 86372 42576 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 42076 86372 42776 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 40276 1014 40976 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 40476 27272 40776 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 40526 54622 40728 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 40527 86372 40728 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 40476 86372 40776 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 40276 86372 40976 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 38476 1014 39176 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 38676 27272 38976 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 38726 54622 38928 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 38727 86372 38928 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 38676 86372 38976 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 38476 86372 39176 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 36676 1014 37376 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 36876 27272 37176 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 30403 36926 54622 37128 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 36927 86372 37128 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60471 36876 86372 37176 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 36676 86372 37376 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60559 34536 60647 35387 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60282 35158 86372 35298 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60282 34536 86372 35016 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 34536 86372 35326 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 83360 35126 86372 35326 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 57295 26435 86372 26890 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 58785 26435 84717 28434 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 58785 26435 86372 28416 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 21282 1014 22282 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 24036 21826 27826 22282 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 21827 27826 22282 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 27387 21826 27826 23199 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 56078 21826 57677 23199 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 27387 22291 57677 23199 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 56078 21826 83763 22282 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 21282 86372 22282 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 56078 21827 86372 22282 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 14328 23678 17730 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 14328 24250 16597 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 24111 14329 27828 16598 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 29478 13243 45977 15015 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 27387 13245 45977 15015 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 14491 47683 15015 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 41493 13078 49775 13760 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 14936 51760 15015 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 14966 55645 15015 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 46982 14968 86372 16784 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 57295 14327 83763 16784 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 61760 14328 86372 17730 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 42261 10740 57736 11527 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 57295 10176 86372 11491 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60736 10173 84482 11491 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 61825 10176 86372 11493 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 5766 1014 7596 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 5766 3011 6199 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 6982 3011 7596 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 2249 6980 24250 7595 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 2226 6981 24250 7595 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 23625 6982 27828 7596 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 23687 6177 41397 6199 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 29458 5665 34622 6573 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 5766 34622 6198 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 29458 6177 41397 6573 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 34860 6177 41397 8582 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 29513 7900 41397 8582 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 34860 6592 55482 7392 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 41857 9165 51430 10420 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 50922 5605 55482 9502 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 50922 6984 57736 8965 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 57295 6982 86372 7595 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 50922 5766 62429 6199 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 50922 6984 62747 7596 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 50922 5766 86372 6198 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60736 6980 84787 7595 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 83361 5766 86372 6199 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 5766 86372 7596 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 83361 6982 86372 7596 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 2502 1014 3772 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 3420 3011 3772 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 3421 24341 3772 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 27438 3524 27778 3876 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 28764 3524 28894 3876 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 41774 3524 41904 3876 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 42299 3524 42429 3876 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 46873 3524 47003 3876 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 47321 3524 47451 3876 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 47769 3524 47899 3876 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 48217 3524 48347 3876 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 23909 3524 61215 3875 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 57345 3524 61215 3876 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 0 2502 86372 2854 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 60699 3420 86372 3772 1 VSS
port 29 nsew ground bidirectional
rlabel metal3 s 85358 2502 86372 3772 1 VSS
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 86372 68176
string GDS_END 2452518
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2396452
string LEFclass BLOCK
string LEFsymmetry X Y R90
string path 287.790 11.160 287.790 0.000 
<< end >>
