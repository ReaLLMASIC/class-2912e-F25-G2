magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
use via1_x2_R90_128x8m81  via1_x2_R90_128x8m81_0
timestamp 1749760379
transform 1 0 0 0 1 0
box 0 0 1 1
use via2_x2_R90_128x8m81  via2_x2_R90_128x8m81_0
timestamp 1749760379
transform 1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 308936
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 308844
<< end >>
