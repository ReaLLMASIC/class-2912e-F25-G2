magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< deepnwell >>
rect -680 -680 1680 1680
<< pbase >>
rect -180 -180 1180 1180
<< ndiff >>
rect 0 943 1000 1000
rect 0 897 57 943
rect 103 897 177 943
rect 223 897 297 943
rect 343 897 417 943
rect 463 897 537 943
rect 583 897 657 943
rect 703 897 777 943
rect 823 897 897 943
rect 943 897 1000 943
rect 0 823 1000 897
rect 0 777 57 823
rect 103 777 177 823
rect 223 777 297 823
rect 343 777 417 823
rect 463 777 537 823
rect 583 777 657 823
rect 703 777 777 823
rect 823 777 897 823
rect 943 777 1000 823
rect 0 703 1000 777
rect 0 657 57 703
rect 103 657 177 703
rect 223 657 297 703
rect 343 657 417 703
rect 463 657 537 703
rect 583 657 657 703
rect 703 657 777 703
rect 823 657 897 703
rect 943 657 1000 703
rect 0 583 1000 657
rect 0 537 57 583
rect 103 537 177 583
rect 223 537 297 583
rect 343 537 417 583
rect 463 537 537 583
rect 583 537 657 583
rect 703 537 777 583
rect 823 537 897 583
rect 943 537 1000 583
rect 0 463 1000 537
rect 0 417 57 463
rect 103 417 177 463
rect 223 417 297 463
rect 343 417 417 463
rect 463 417 537 463
rect 583 417 657 463
rect 703 417 777 463
rect 823 417 897 463
rect 943 417 1000 463
rect 0 343 1000 417
rect 0 297 57 343
rect 103 297 177 343
rect 223 297 297 343
rect 343 297 417 343
rect 463 297 537 343
rect 583 297 657 343
rect 703 297 777 343
rect 823 297 897 343
rect 943 297 1000 343
rect 0 223 1000 297
rect 0 177 57 223
rect 103 177 177 223
rect 223 177 297 223
rect 343 177 417 223
rect 463 177 537 223
rect 583 177 657 223
rect 703 177 777 223
rect 823 177 897 223
rect 943 177 1000 223
rect 0 103 1000 177
rect 0 57 57 103
rect 103 57 177 103
rect 223 57 297 103
rect 343 57 417 103
rect 463 57 537 103
rect 583 57 657 103
rect 703 57 777 103
rect 823 57 897 103
rect 943 57 1000 103
rect 0 0 1000 57
<< ndiffc >>
rect 57 897 103 943
rect 177 897 223 943
rect 297 897 343 943
rect 417 897 463 943
rect 537 897 583 943
rect 657 897 703 943
rect 777 897 823 943
rect 897 897 943 943
rect 57 777 103 823
rect 177 777 223 823
rect 297 777 343 823
rect 417 777 463 823
rect 537 777 583 823
rect 657 777 703 823
rect 777 777 823 823
rect 897 777 943 823
rect 57 657 103 703
rect 177 657 223 703
rect 297 657 343 703
rect 417 657 463 703
rect 537 657 583 703
rect 657 657 703 703
rect 777 657 823 703
rect 897 657 943 703
rect 57 537 103 583
rect 177 537 223 583
rect 297 537 343 583
rect 417 537 463 583
rect 537 537 583 583
rect 657 537 703 583
rect 777 537 823 583
rect 897 537 943 583
rect 57 417 103 463
rect 177 417 223 463
rect 297 417 343 463
rect 417 417 463 463
rect 537 417 583 463
rect 657 417 703 463
rect 777 417 823 463
rect 897 417 943 463
rect 57 297 103 343
rect 177 297 223 343
rect 297 297 343 343
rect 417 297 463 343
rect 537 297 583 343
rect 657 297 703 343
rect 777 297 823 343
rect 897 297 943 343
rect 57 177 103 223
rect 177 177 223 223
rect 297 177 343 223
rect 417 177 463 223
rect 537 177 583 223
rect 657 177 703 223
rect 777 177 823 223
rect 897 177 943 223
rect 57 57 103 103
rect 177 57 223 103
rect 297 57 343 103
rect 417 57 463 103
rect 537 57 583 103
rect 657 57 703 103
rect 777 57 823 103
rect 897 57 943 103
<< psubdiff >>
rect -1264 2245 2264 2264
rect -1264 2199 -1074 2245
rect 2074 2199 2264 2245
rect -1264 2180 2264 2199
rect -1264 2074 -1180 2180
rect -1264 -1074 -1245 2074
rect -1199 -1074 -1180 2074
rect 2180 2074 2264 2180
rect -148 1129 1148 1148
rect -148 1083 -87 1129
rect 1087 1083 1148 1129
rect -148 1064 1148 1083
rect -148 999 -64 1064
rect -148 -81 -129 999
rect -83 -64 -64 999
rect 1064 999 1148 1064
rect 1064 -64 1083 999
rect -83 -81 1083 -64
rect 1129 -81 1148 999
rect -148 -148 1148 -81
rect -1264 -1180 -1180 -1074
rect 2180 -1074 2199 2074
rect 2245 -1074 2264 2074
rect 2180 -1180 2264 -1074
rect -1264 -1199 2264 -1180
rect -1264 -1245 -1074 -1199
rect -746 -1245 1746 -1199
rect 2074 -1245 2264 -1199
rect -1264 -1264 2264 -1245
<< nsubdiff >>
rect -296 1277 1296 1296
rect -296 1231 -229 1277
rect 1227 1231 1296 1277
rect -296 1212 1296 1231
rect -296 1181 -212 1212
rect -296 -275 -277 1181
rect -231 -212 -212 1181
rect 1212 1181 1296 1212
rect 1212 -212 1231 1181
rect -231 -275 1231 -212
rect 1277 -275 1296 1181
rect -296 -296 1296 -275
<< psubdiffcont >>
rect -1074 2199 2074 2245
rect -1245 -1074 -1199 2074
rect -87 1083 1087 1129
rect -129 -81 -83 999
rect 1083 -81 1129 999
rect 2199 -1074 2245 2074
rect -1074 -1245 -746 -1199
rect 1746 -1245 2074 -1199
<< nsubdiffcont >>
rect -229 1231 1227 1277
rect -277 -275 -231 1181
rect 1231 -275 1277 1181
<< metal1 >>
rect -1264 2245 2264 2264
rect -1264 2199 -1074 2245
rect 2074 2199 2264 2245
rect -1264 2180 2264 2199
rect -1264 2074 -1180 2180
rect -1264 -1074 -1245 2074
rect -1199 -1074 -1180 2074
rect 2180 2074 2264 2180
rect -296 1277 1296 1296
rect -296 1231 -229 1277
rect 1227 1231 1296 1277
rect -296 1212 1296 1231
rect -296 1181 -212 1212
rect -296 -275 -277 1181
rect -231 -275 -212 1181
rect 1212 1181 1296 1212
rect -148 1129 1148 1148
rect -148 1083 -87 1129
rect 1087 1083 1148 1129
rect -148 1064 1148 1083
rect -148 999 -64 1064
rect -148 -81 -129 999
rect -83 -81 -64 999
rect 0 943 1000 1000
rect 0 897 57 943
rect 103 897 177 943
rect 223 897 297 943
rect 343 897 417 943
rect 463 897 537 943
rect 583 897 657 943
rect 703 897 777 943
rect 823 897 897 943
rect 943 897 1000 943
rect 0 823 1000 897
rect 0 777 57 823
rect 103 777 177 823
rect 223 777 297 823
rect 343 777 417 823
rect 463 777 537 823
rect 583 777 657 823
rect 703 777 777 823
rect 823 777 897 823
rect 943 777 1000 823
rect 0 703 1000 777
rect 0 657 57 703
rect 103 657 177 703
rect 223 657 297 703
rect 343 657 417 703
rect 463 657 537 703
rect 583 657 657 703
rect 703 657 777 703
rect 823 657 897 703
rect 943 657 1000 703
rect 0 583 1000 657
rect 0 537 57 583
rect 103 537 177 583
rect 223 537 297 583
rect 343 537 417 583
rect 463 537 537 583
rect 583 537 657 583
rect 703 537 777 583
rect 823 537 897 583
rect 943 537 1000 583
rect 0 463 1000 537
rect 0 417 57 463
rect 103 417 177 463
rect 223 417 297 463
rect 343 417 417 463
rect 463 417 537 463
rect 583 417 657 463
rect 703 417 777 463
rect 823 417 897 463
rect 943 417 1000 463
rect 0 343 1000 417
rect 0 297 57 343
rect 103 297 177 343
rect 223 297 297 343
rect 343 297 417 343
rect 463 297 537 343
rect 583 297 657 343
rect 703 297 777 343
rect 823 297 897 343
rect 943 297 1000 343
rect 0 223 1000 297
rect 0 177 57 223
rect 103 177 177 223
rect 223 177 297 223
rect 343 177 417 223
rect 463 177 537 223
rect 583 177 657 223
rect 703 177 777 223
rect 823 177 897 223
rect 943 177 1000 223
rect 0 103 1000 177
rect 0 57 57 103
rect 103 57 177 103
rect 223 57 297 103
rect 343 57 417 103
rect 463 57 537 103
rect 583 57 657 103
rect 703 57 777 103
rect 823 57 897 103
rect 943 57 1000 103
rect 0 0 1000 57
rect 1064 999 1148 1064
rect -148 -148 -64 -81
rect 1064 -81 1083 999
rect 1129 -81 1148 999
rect 1064 -148 1148 -81
rect -296 -296 -212 -275
rect 1212 -275 1231 1181
rect 1277 -275 1296 1181
rect 1212 -296 1296 -275
rect -1264 -1180 -1180 -1074
rect 2180 -1074 2199 2074
rect 2245 -1074 2264 2074
rect 2180 -1180 2264 -1074
rect -1264 -1199 -680 -1180
rect -1264 -1245 -1074 -1199
rect -746 -1245 -680 -1199
rect -1264 -1264 -680 -1245
rect 1680 -1199 2264 -1180
rect 1680 -1245 1746 -1199
rect 2074 -1245 2264 -1199
rect 1680 -1264 2264 -1245
<< labels >>
flabel metal1 -1215 -1215 -1215 -1215 0 FreeSans 400 0 0 0 S
flabel metal1 -1215 -1215 -1215 -1215 0 FreeSans 400 0 0 0 S
flabel metal1 2221 -1216 2221 -1216 0 FreeSans 400 0 0 0 S
flabel metal1 2221 -1216 2221 -1216 0 FreeSans 400 0 0 0 S
flabel metal1 2224 2224 2224 2224 0 FreeSans 400 0 0 0 S
flabel metal1 497 545 497 545 0 FreeSans 400 0 0 0 E
flabel metal1 1107 -97 1107 -97 0 FreeSans 400 0 0 0 B
flabel metal1 1107 1108 1107 1108 0 FreeSans 400 0 0 0 B
flabel metal1 -103 -86 -103 -86 0 FreeSans 400 0 0 0 B
flabel metal1 -255 1248 -255 1248 0 FreeSans 400 0 0 0 C
flabel nsubdiffcont 1256 -248 1256 -248 0 FreeSans 400 0 0 0 C
flabel metal1 1259 1253 1259 1253 0 FreeSans 400 0 0 0 C
<< properties >>
string GDS_END 19692
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/npn_05p00x05p00.gds
string GDS_START 112
string gencell npn_05p00x05p00
string library gf180mcu
string parameter m=1
<< end >>
