magic
tech gf180mcuD
timestamp 1749760379
<< properties >>
string GDS_END 3641678
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 3640010
<< end >>
