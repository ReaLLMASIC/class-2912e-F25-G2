magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
use xdec_512x8m81  xdec_512x8m81_0
timestamp 1749760379
transform 1 0 1 0 -1 6300
box 1425 0 22888 901
use xdec_512x8m81  xdec_512x8m81_1
timestamp 1749760379
transform 1 0 1 0 -1 4500
box 1425 0 22888 901
use xdec_512x8m81  xdec_512x8m81_2
timestamp 1749760379
transform 1 0 1 0 -1 2700
box 1425 0 22888 901
use xdec_512x8m81  xdec_512x8m81_3
timestamp 1749760379
transform 1 0 1 0 -1 900
box 1425 0 22888 901
use xdec_512x8m81  xdec_512x8m81_4
timestamp 1749760379
transform 1 0 1 0 1 6300
box 1425 0 22888 901
use xdec_512x8m81  xdec_512x8m81_5
timestamp 1749760379
transform 1 0 1 0 1 4500
box 1425 0 22888 901
use xdec_512x8m81  xdec_512x8m81_6
timestamp 1749760379
transform 1 0 1 0 1 2700
box 1425 0 22888 901
use xdec_512x8m81  xdec_512x8m81_7
timestamp 1749760379
transform 1 0 1 0 1 900
box 1425 0 22888 901
<< properties >>
string GDS_END 789880
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 785124
<< end >>
