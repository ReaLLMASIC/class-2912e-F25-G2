magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< pwell >>
rect 559 6633 2735 11633
rect 2995 6633 5171 11633
rect 5431 6633 7607 11633
rect 7867 6633 10043 11633
rect 5431 621 7607 5621
rect 7867 621 10043 5621
<< mvndiff >>
rect 559 11596 647 11633
rect 559 6670 572 11596
rect 618 6670 647 11596
rect 559 6633 647 6670
rect 2647 11596 2735 11633
rect 2647 6670 2676 11596
rect 2722 6670 2735 11596
rect 2647 6633 2735 6670
rect 2995 11596 3083 11633
rect 2995 6670 3008 11596
rect 3054 6670 3083 11596
rect 2995 6633 3083 6670
rect 5083 11596 5171 11633
rect 5083 6670 5112 11596
rect 5158 6670 5171 11596
rect 5083 6633 5171 6670
rect 5431 11596 5519 11633
rect 5431 6670 5444 11596
rect 5490 6670 5519 11596
rect 5431 6633 5519 6670
rect 7519 11596 7607 11633
rect 7519 6670 7548 11596
rect 7594 6670 7607 11596
rect 7519 6633 7607 6670
rect 7867 11596 7955 11633
rect 7867 6670 7880 11596
rect 7926 6670 7955 11596
rect 7867 6633 7955 6670
rect 9955 11596 10043 11633
rect 9955 6670 9984 11596
rect 10030 6670 10043 11596
rect 9955 6633 10043 6670
rect 5431 5584 5519 5621
rect 5431 658 5444 5584
rect 5490 658 5519 5584
rect 5431 621 5519 658
rect 7519 5584 7607 5621
rect 7519 658 7548 5584
rect 7594 658 7607 5584
rect 7519 621 7607 658
rect 7867 5584 7955 5621
rect 7867 658 7880 5584
rect 7926 658 7955 5584
rect 7867 621 7955 658
rect 9955 5584 10043 5621
rect 9955 658 9984 5584
rect 10030 658 10043 5584
rect 9955 621 10043 658
<< mvndiffc >>
rect 572 6670 618 11596
rect 2676 6670 2722 11596
rect 3008 6670 3054 11596
rect 5112 6670 5158 11596
rect 5444 6670 5490 11596
rect 7548 6670 7594 11596
rect 7880 6670 7926 11596
rect 9984 6670 10030 11596
rect 5444 658 5490 5584
rect 7548 658 7594 5584
rect 7880 658 7926 5584
rect 9984 658 10030 5584
<< psubdiff >>
rect 32 12298 10576 12320
rect 32 12252 54 12298
rect 100 12252 168 12298
rect 214 12252 322 12298
rect 368 12252 436 12298
rect 482 12252 550 12298
rect 596 12252 664 12298
rect 710 12252 778 12298
rect 824 12252 892 12298
rect 938 12252 1006 12298
rect 1052 12252 1120 12298
rect 1166 12252 1234 12298
rect 1280 12252 1348 12298
rect 1394 12252 1462 12298
rect 1508 12252 1576 12298
rect 1622 12252 1690 12298
rect 1736 12252 1804 12298
rect 1850 12252 1918 12298
rect 1964 12252 2032 12298
rect 2078 12252 2146 12298
rect 2192 12252 2260 12298
rect 2306 12252 2374 12298
rect 2420 12252 2488 12298
rect 2534 12252 2602 12298
rect 2648 12252 2716 12298
rect 2762 12252 2830 12298
rect 2876 12252 2944 12298
rect 2990 12252 3058 12298
rect 3104 12252 3172 12298
rect 3218 12252 3286 12298
rect 3332 12252 3400 12298
rect 3446 12252 3514 12298
rect 3560 12252 3628 12298
rect 3674 12252 3742 12298
rect 3788 12252 3856 12298
rect 3902 12252 3970 12298
rect 4016 12252 4084 12298
rect 4130 12252 4198 12298
rect 4244 12252 4312 12298
rect 4358 12252 4426 12298
rect 4472 12252 4540 12298
rect 4586 12252 4654 12298
rect 4700 12252 4768 12298
rect 4814 12252 4882 12298
rect 4928 12252 4996 12298
rect 5042 12252 5110 12298
rect 5156 12252 5224 12298
rect 5270 12252 5338 12298
rect 5384 12252 5452 12298
rect 5498 12252 5566 12298
rect 5612 12252 5680 12298
rect 5726 12252 5794 12298
rect 5840 12252 5908 12298
rect 5954 12252 6022 12298
rect 6068 12252 6136 12298
rect 6182 12252 6250 12298
rect 6296 12252 6364 12298
rect 6410 12252 6478 12298
rect 6524 12252 6592 12298
rect 6638 12252 6706 12298
rect 6752 12252 6820 12298
rect 6866 12252 6934 12298
rect 6980 12252 7048 12298
rect 7094 12252 7162 12298
rect 7208 12252 7276 12298
rect 7322 12252 7390 12298
rect 7436 12252 7504 12298
rect 7550 12252 7618 12298
rect 7664 12252 7732 12298
rect 7778 12252 7846 12298
rect 7892 12252 7960 12298
rect 8006 12252 8074 12298
rect 8120 12252 8188 12298
rect 8234 12252 8302 12298
rect 8348 12252 8416 12298
rect 8462 12252 8530 12298
rect 8576 12252 8644 12298
rect 8690 12252 8758 12298
rect 8804 12252 8872 12298
rect 8918 12252 8986 12298
rect 9032 12252 9100 12298
rect 9146 12252 9214 12298
rect 9260 12252 9328 12298
rect 9374 12252 9442 12298
rect 9488 12252 9556 12298
rect 9602 12252 9670 12298
rect 9716 12252 9784 12298
rect 9830 12252 9898 12298
rect 9944 12252 10012 12298
rect 10058 12252 10126 12298
rect 10172 12252 10240 12298
rect 10286 12252 10394 12298
rect 10440 12252 10508 12298
rect 10554 12252 10576 12298
rect 32 12184 10576 12252
rect 32 12138 54 12184
rect 100 12138 168 12184
rect 214 12138 322 12184
rect 368 12138 436 12184
rect 482 12138 550 12184
rect 596 12138 664 12184
rect 710 12138 778 12184
rect 824 12138 892 12184
rect 938 12138 1006 12184
rect 1052 12138 1120 12184
rect 1166 12138 1234 12184
rect 1280 12138 1348 12184
rect 1394 12138 1462 12184
rect 1508 12138 1576 12184
rect 1622 12138 1690 12184
rect 1736 12138 1804 12184
rect 1850 12138 1918 12184
rect 1964 12138 2032 12184
rect 2078 12138 2146 12184
rect 2192 12138 2260 12184
rect 2306 12138 2374 12184
rect 2420 12138 2488 12184
rect 2534 12138 2602 12184
rect 2648 12138 2716 12184
rect 2762 12138 2830 12184
rect 2876 12138 2944 12184
rect 2990 12138 3058 12184
rect 3104 12138 3172 12184
rect 3218 12138 3286 12184
rect 3332 12138 3400 12184
rect 3446 12138 3514 12184
rect 3560 12138 3628 12184
rect 3674 12138 3742 12184
rect 3788 12138 3856 12184
rect 3902 12138 3970 12184
rect 4016 12138 4084 12184
rect 4130 12138 4198 12184
rect 4244 12138 4312 12184
rect 4358 12138 4426 12184
rect 4472 12138 4540 12184
rect 4586 12138 4654 12184
rect 4700 12138 4768 12184
rect 4814 12138 4882 12184
rect 4928 12138 4996 12184
rect 5042 12138 5110 12184
rect 5156 12138 5224 12184
rect 5270 12138 5338 12184
rect 5384 12138 5452 12184
rect 5498 12138 5566 12184
rect 5612 12138 5680 12184
rect 5726 12138 5794 12184
rect 5840 12138 5908 12184
rect 5954 12138 6022 12184
rect 6068 12138 6136 12184
rect 6182 12138 6250 12184
rect 6296 12138 6364 12184
rect 6410 12138 6478 12184
rect 6524 12138 6592 12184
rect 6638 12138 6706 12184
rect 6752 12138 6820 12184
rect 6866 12138 6934 12184
rect 6980 12138 7048 12184
rect 7094 12138 7162 12184
rect 7208 12138 7276 12184
rect 7322 12138 7390 12184
rect 7436 12138 7504 12184
rect 7550 12138 7618 12184
rect 7664 12138 7732 12184
rect 7778 12138 7846 12184
rect 7892 12138 7960 12184
rect 8006 12138 8074 12184
rect 8120 12138 8188 12184
rect 8234 12138 8302 12184
rect 8348 12138 8416 12184
rect 8462 12138 8530 12184
rect 8576 12138 8644 12184
rect 8690 12138 8758 12184
rect 8804 12138 8872 12184
rect 8918 12138 8986 12184
rect 9032 12138 9100 12184
rect 9146 12138 9214 12184
rect 9260 12138 9328 12184
rect 9374 12138 9442 12184
rect 9488 12138 9556 12184
rect 9602 12138 9670 12184
rect 9716 12138 9784 12184
rect 9830 12138 9898 12184
rect 9944 12138 10012 12184
rect 10058 12138 10126 12184
rect 10172 12138 10240 12184
rect 10286 12138 10394 12184
rect 10440 12138 10508 12184
rect 10554 12138 10576 12184
rect 32 12116 10576 12138
rect 32 12070 236 12116
rect 32 12024 54 12070
rect 100 12024 168 12070
rect 214 12024 236 12070
rect 32 11500 236 12024
rect 10372 12070 10576 12116
rect 10372 12024 10394 12070
rect 10440 12024 10508 12070
rect 10554 12024 10576 12070
rect 10372 11956 10576 12024
rect 10372 11910 10394 11956
rect 10440 11910 10508 11956
rect 10554 11910 10576 11956
rect 10372 11842 10576 11910
rect 10372 11796 10394 11842
rect 10440 11796 10508 11842
rect 10554 11796 10576 11842
rect 10372 11728 10576 11796
rect 10372 11682 10394 11728
rect 10440 11682 10508 11728
rect 10554 11682 10576 11728
rect 32 11454 54 11500
rect 100 11454 168 11500
rect 214 11454 236 11500
rect 32 11386 236 11454
rect 32 11340 54 11386
rect 100 11340 168 11386
rect 214 11340 236 11386
rect 32 11272 236 11340
rect 32 11226 54 11272
rect 100 11226 168 11272
rect 214 11226 236 11272
rect 32 11158 236 11226
rect 32 11112 54 11158
rect 100 11112 168 11158
rect 214 11112 236 11158
rect 32 11044 236 11112
rect 32 10998 54 11044
rect 100 10998 168 11044
rect 214 10998 236 11044
rect 32 10930 236 10998
rect 32 10884 54 10930
rect 100 10884 168 10930
rect 214 10884 236 10930
rect 32 10816 236 10884
rect 32 10770 54 10816
rect 100 10770 168 10816
rect 214 10770 236 10816
rect 32 10702 236 10770
rect 32 10656 54 10702
rect 100 10656 168 10702
rect 214 10656 236 10702
rect 32 10588 236 10656
rect 32 10542 54 10588
rect 100 10542 168 10588
rect 214 10542 236 10588
rect 32 10474 236 10542
rect 32 10428 54 10474
rect 100 10428 168 10474
rect 214 10428 236 10474
rect 32 10360 236 10428
rect 32 10314 54 10360
rect 100 10314 168 10360
rect 214 10314 236 10360
rect 32 10246 236 10314
rect 32 10200 54 10246
rect 100 10200 168 10246
rect 214 10200 236 10246
rect 32 10132 236 10200
rect 32 10086 54 10132
rect 100 10086 168 10132
rect 214 10086 236 10132
rect 32 10018 236 10086
rect 32 9972 54 10018
rect 100 9972 168 10018
rect 214 9972 236 10018
rect 32 9904 236 9972
rect 32 9858 54 9904
rect 100 9858 168 9904
rect 214 9858 236 9904
rect 32 9790 236 9858
rect 32 9744 54 9790
rect 100 9744 168 9790
rect 214 9744 236 9790
rect 32 9676 236 9744
rect 32 9630 54 9676
rect 100 9630 168 9676
rect 214 9630 236 9676
rect 32 9562 236 9630
rect 32 9516 54 9562
rect 100 9516 168 9562
rect 214 9516 236 9562
rect 32 9448 236 9516
rect 32 9402 54 9448
rect 100 9402 168 9448
rect 214 9402 236 9448
rect 32 9334 236 9402
rect 32 9288 54 9334
rect 100 9288 168 9334
rect 214 9288 236 9334
rect 32 9220 236 9288
rect 32 9174 54 9220
rect 100 9174 168 9220
rect 214 9174 236 9220
rect 32 9106 236 9174
rect 32 9060 54 9106
rect 100 9060 168 9106
rect 214 9060 236 9106
rect 32 8992 236 9060
rect 32 8946 54 8992
rect 100 8946 168 8992
rect 214 8946 236 8992
rect 32 8878 236 8946
rect 32 8832 54 8878
rect 100 8832 168 8878
rect 214 8832 236 8878
rect 32 8764 236 8832
rect 32 8718 54 8764
rect 100 8718 168 8764
rect 214 8718 236 8764
rect 32 8650 236 8718
rect 32 8604 54 8650
rect 100 8604 168 8650
rect 214 8604 236 8650
rect 32 8536 236 8604
rect 32 8490 54 8536
rect 100 8490 168 8536
rect 214 8490 236 8536
rect 32 8422 236 8490
rect 32 8376 54 8422
rect 100 8376 168 8422
rect 214 8376 236 8422
rect 32 8308 236 8376
rect 32 8262 54 8308
rect 100 8262 168 8308
rect 214 8262 236 8308
rect 32 8194 236 8262
rect 32 8148 54 8194
rect 100 8148 168 8194
rect 214 8148 236 8194
rect 32 8080 236 8148
rect 32 8034 54 8080
rect 100 8034 168 8080
rect 214 8034 236 8080
rect 32 7966 236 8034
rect 32 7920 54 7966
rect 100 7920 168 7966
rect 214 7920 236 7966
rect 32 7852 236 7920
rect 32 7806 54 7852
rect 100 7806 168 7852
rect 214 7806 236 7852
rect 32 7738 236 7806
rect 32 7692 54 7738
rect 100 7692 168 7738
rect 214 7692 236 7738
rect 32 7624 236 7692
rect 32 7578 54 7624
rect 100 7578 168 7624
rect 214 7578 236 7624
rect 32 7510 236 7578
rect 32 7464 54 7510
rect 100 7464 168 7510
rect 214 7464 236 7510
rect 32 7396 236 7464
rect 32 7350 54 7396
rect 100 7350 168 7396
rect 214 7350 236 7396
rect 32 7282 236 7350
rect 32 7236 54 7282
rect 100 7236 168 7282
rect 214 7236 236 7282
rect 32 7168 236 7236
rect 32 7122 54 7168
rect 100 7122 168 7168
rect 214 7122 236 7168
rect 32 7054 236 7122
rect 32 7008 54 7054
rect 100 7008 168 7054
rect 214 7008 236 7054
rect 32 6940 236 7008
rect 32 6894 54 6940
rect 100 6894 168 6940
rect 214 6894 236 6940
rect 32 6826 236 6894
rect 32 6780 54 6826
rect 100 6780 168 6826
rect 214 6780 236 6826
rect 32 6712 236 6780
rect 32 6666 54 6712
rect 100 6666 168 6712
rect 214 6666 236 6712
rect 32 6598 236 6666
rect 10372 11614 10576 11682
rect 10372 11568 10394 11614
rect 10440 11568 10508 11614
rect 10554 11568 10576 11614
rect 10372 11500 10576 11568
rect 10372 11454 10394 11500
rect 10440 11454 10508 11500
rect 10554 11454 10576 11500
rect 10372 11386 10576 11454
rect 10372 11340 10394 11386
rect 10440 11340 10508 11386
rect 10554 11340 10576 11386
rect 10372 11272 10576 11340
rect 10372 11226 10394 11272
rect 10440 11226 10508 11272
rect 10554 11226 10576 11272
rect 10372 11158 10576 11226
rect 10372 11112 10394 11158
rect 10440 11112 10508 11158
rect 10554 11112 10576 11158
rect 10372 11044 10576 11112
rect 10372 10998 10394 11044
rect 10440 10998 10508 11044
rect 10554 10998 10576 11044
rect 10372 10930 10576 10998
rect 10372 10884 10394 10930
rect 10440 10884 10508 10930
rect 10554 10884 10576 10930
rect 10372 10816 10576 10884
rect 10372 10770 10394 10816
rect 10440 10770 10508 10816
rect 10554 10770 10576 10816
rect 10372 10702 10576 10770
rect 10372 10656 10394 10702
rect 10440 10656 10508 10702
rect 10554 10656 10576 10702
rect 10372 10588 10576 10656
rect 10372 10542 10394 10588
rect 10440 10542 10508 10588
rect 10554 10542 10576 10588
rect 10372 10474 10576 10542
rect 10372 10428 10394 10474
rect 10440 10428 10508 10474
rect 10554 10428 10576 10474
rect 10372 10360 10576 10428
rect 10372 10314 10394 10360
rect 10440 10314 10508 10360
rect 10554 10314 10576 10360
rect 10372 10246 10576 10314
rect 10372 10200 10394 10246
rect 10440 10200 10508 10246
rect 10554 10200 10576 10246
rect 10372 10132 10576 10200
rect 10372 10086 10394 10132
rect 10440 10086 10508 10132
rect 10554 10086 10576 10132
rect 10372 10018 10576 10086
rect 10372 9972 10394 10018
rect 10440 9972 10508 10018
rect 10554 9972 10576 10018
rect 10372 9904 10576 9972
rect 10372 9858 10394 9904
rect 10440 9858 10508 9904
rect 10554 9858 10576 9904
rect 10372 9790 10576 9858
rect 10372 9744 10394 9790
rect 10440 9744 10508 9790
rect 10554 9744 10576 9790
rect 10372 9676 10576 9744
rect 10372 9630 10394 9676
rect 10440 9630 10508 9676
rect 10554 9630 10576 9676
rect 10372 9562 10576 9630
rect 10372 9516 10394 9562
rect 10440 9516 10508 9562
rect 10554 9516 10576 9562
rect 10372 9448 10576 9516
rect 10372 9402 10394 9448
rect 10440 9402 10508 9448
rect 10554 9402 10576 9448
rect 10372 9334 10576 9402
rect 10372 9288 10394 9334
rect 10440 9288 10508 9334
rect 10554 9288 10576 9334
rect 10372 9220 10576 9288
rect 10372 9174 10394 9220
rect 10440 9174 10508 9220
rect 10554 9174 10576 9220
rect 10372 9106 10576 9174
rect 10372 9060 10394 9106
rect 10440 9060 10508 9106
rect 10554 9060 10576 9106
rect 10372 8992 10576 9060
rect 10372 8946 10394 8992
rect 10440 8946 10508 8992
rect 10554 8946 10576 8992
rect 10372 8878 10576 8946
rect 10372 8832 10394 8878
rect 10440 8832 10508 8878
rect 10554 8832 10576 8878
rect 10372 8764 10576 8832
rect 10372 8718 10394 8764
rect 10440 8718 10508 8764
rect 10554 8718 10576 8764
rect 10372 8650 10576 8718
rect 10372 8604 10394 8650
rect 10440 8604 10508 8650
rect 10554 8604 10576 8650
rect 10372 8536 10576 8604
rect 10372 8490 10394 8536
rect 10440 8490 10508 8536
rect 10554 8490 10576 8536
rect 10372 8422 10576 8490
rect 10372 8376 10394 8422
rect 10440 8376 10508 8422
rect 10554 8376 10576 8422
rect 10372 8308 10576 8376
rect 10372 8262 10394 8308
rect 10440 8262 10508 8308
rect 10554 8262 10576 8308
rect 10372 8194 10576 8262
rect 10372 8148 10394 8194
rect 10440 8148 10508 8194
rect 10554 8148 10576 8194
rect 10372 8080 10576 8148
rect 10372 8034 10394 8080
rect 10440 8034 10508 8080
rect 10554 8034 10576 8080
rect 10372 7966 10576 8034
rect 10372 7920 10394 7966
rect 10440 7920 10508 7966
rect 10554 7920 10576 7966
rect 10372 7852 10576 7920
rect 10372 7806 10394 7852
rect 10440 7806 10508 7852
rect 10554 7806 10576 7852
rect 10372 7738 10576 7806
rect 10372 7692 10394 7738
rect 10440 7692 10508 7738
rect 10554 7692 10576 7738
rect 10372 7624 10576 7692
rect 10372 7578 10394 7624
rect 10440 7578 10508 7624
rect 10554 7578 10576 7624
rect 10372 7510 10576 7578
rect 10372 7464 10394 7510
rect 10440 7464 10508 7510
rect 10554 7464 10576 7510
rect 10372 7396 10576 7464
rect 10372 7350 10394 7396
rect 10440 7350 10508 7396
rect 10554 7350 10576 7396
rect 10372 7282 10576 7350
rect 10372 7236 10394 7282
rect 10440 7236 10508 7282
rect 10554 7236 10576 7282
rect 10372 7168 10576 7236
rect 10372 7122 10394 7168
rect 10440 7122 10508 7168
rect 10554 7122 10576 7168
rect 10372 7054 10576 7122
rect 10372 7008 10394 7054
rect 10440 7008 10508 7054
rect 10554 7008 10576 7054
rect 10372 6940 10576 7008
rect 10372 6894 10394 6940
rect 10440 6894 10508 6940
rect 10554 6894 10576 6940
rect 10372 6826 10576 6894
rect 10372 6780 10394 6826
rect 10440 6780 10508 6826
rect 10554 6780 10576 6826
rect 10372 6712 10576 6780
rect 10372 6666 10394 6712
rect 10440 6666 10508 6712
rect 10554 6666 10576 6712
rect 32 6552 54 6598
rect 100 6552 168 6598
rect 214 6552 236 6598
rect 32 6484 236 6552
rect 10372 6598 10576 6666
rect 10372 6552 10394 6598
rect 10440 6552 10508 6598
rect 10554 6552 10576 6598
rect 32 6438 54 6484
rect 100 6438 168 6484
rect 214 6438 236 6484
rect 32 6370 236 6438
rect 32 6324 54 6370
rect 100 6324 168 6370
rect 214 6324 236 6370
rect 32 6229 236 6324
rect 10372 6484 10576 6552
rect 10372 6438 10394 6484
rect 10440 6438 10508 6484
rect 10554 6438 10576 6484
rect 10372 6370 10576 6438
rect 10372 6324 10394 6370
rect 10440 6324 10508 6370
rect 10554 6324 10576 6370
rect 10372 6256 10576 6324
rect 10372 6229 10394 6256
rect 32 6210 10394 6229
rect 10440 6210 10508 6256
rect 10554 6210 10576 6256
rect 32 6207 10576 6210
rect 32 6161 322 6207
rect 368 6161 436 6207
rect 482 6161 550 6207
rect 596 6161 664 6207
rect 710 6161 778 6207
rect 824 6161 892 6207
rect 938 6161 1006 6207
rect 1052 6161 1120 6207
rect 1166 6161 1234 6207
rect 1280 6161 1348 6207
rect 1394 6161 1462 6207
rect 1508 6161 1576 6207
rect 1622 6161 1690 6207
rect 1736 6161 1804 6207
rect 1850 6161 1918 6207
rect 1964 6161 2032 6207
rect 2078 6161 2146 6207
rect 2192 6161 2260 6207
rect 2306 6161 2374 6207
rect 2420 6161 2488 6207
rect 2534 6161 2602 6207
rect 2648 6161 2716 6207
rect 2762 6161 2830 6207
rect 2876 6161 2944 6207
rect 2990 6161 3058 6207
rect 3104 6161 3172 6207
rect 3218 6161 3286 6207
rect 3332 6161 3400 6207
rect 3446 6161 3514 6207
rect 3560 6161 3628 6207
rect 3674 6161 3742 6207
rect 3788 6161 3856 6207
rect 3902 6161 3970 6207
rect 4016 6161 4084 6207
rect 4130 6161 4198 6207
rect 4244 6161 4312 6207
rect 4358 6161 4426 6207
rect 4472 6161 4540 6207
rect 4586 6161 4654 6207
rect 4700 6161 4768 6207
rect 4814 6161 4882 6207
rect 4928 6161 4996 6207
rect 5042 6161 5110 6207
rect 5156 6161 5224 6207
rect 5270 6161 5338 6207
rect 5384 6161 5452 6207
rect 5498 6161 5566 6207
rect 5612 6161 5680 6207
rect 5726 6161 5794 6207
rect 5840 6161 5908 6207
rect 5954 6161 6022 6207
rect 6068 6161 6136 6207
rect 6182 6161 6250 6207
rect 6296 6161 6364 6207
rect 6410 6161 6478 6207
rect 6524 6161 6592 6207
rect 6638 6161 6706 6207
rect 6752 6161 6820 6207
rect 6866 6161 6934 6207
rect 6980 6161 7048 6207
rect 7094 6161 7162 6207
rect 7208 6161 7276 6207
rect 7322 6161 7390 6207
rect 7436 6161 7504 6207
rect 7550 6161 7618 6207
rect 7664 6161 7732 6207
rect 7778 6161 7846 6207
rect 7892 6161 7960 6207
rect 8006 6161 8074 6207
rect 8120 6161 8188 6207
rect 8234 6161 8302 6207
rect 8348 6161 8416 6207
rect 8462 6161 8530 6207
rect 8576 6161 8644 6207
rect 8690 6161 8758 6207
rect 8804 6161 8872 6207
rect 8918 6161 8986 6207
rect 9032 6161 9100 6207
rect 9146 6161 9214 6207
rect 9260 6161 9328 6207
rect 9374 6161 9442 6207
rect 9488 6161 9556 6207
rect 9602 6161 9670 6207
rect 9716 6161 9784 6207
rect 9830 6161 9898 6207
rect 9944 6161 10012 6207
rect 10058 6161 10126 6207
rect 10172 6161 10240 6207
rect 10286 6161 10576 6207
rect 32 6142 10576 6161
rect 32 6096 10394 6142
rect 10440 6096 10508 6142
rect 10554 6096 10576 6142
rect 32 6093 10576 6096
rect 32 6047 322 6093
rect 368 6047 436 6093
rect 482 6047 550 6093
rect 596 6047 664 6093
rect 710 6047 778 6093
rect 824 6047 892 6093
rect 938 6047 1006 6093
rect 1052 6047 1120 6093
rect 1166 6047 1234 6093
rect 1280 6047 1348 6093
rect 1394 6047 1462 6093
rect 1508 6047 1576 6093
rect 1622 6047 1690 6093
rect 1736 6047 1804 6093
rect 1850 6047 1918 6093
rect 1964 6047 2032 6093
rect 2078 6047 2146 6093
rect 2192 6047 2260 6093
rect 2306 6047 2374 6093
rect 2420 6047 2488 6093
rect 2534 6047 2602 6093
rect 2648 6047 2716 6093
rect 2762 6047 2830 6093
rect 2876 6047 2944 6093
rect 2990 6047 3058 6093
rect 3104 6047 3172 6093
rect 3218 6047 3286 6093
rect 3332 6047 3400 6093
rect 3446 6047 3514 6093
rect 3560 6047 3628 6093
rect 3674 6047 3742 6093
rect 3788 6047 3856 6093
rect 3902 6047 3970 6093
rect 4016 6047 4084 6093
rect 4130 6047 4198 6093
rect 4244 6047 4312 6093
rect 4358 6047 4426 6093
rect 4472 6047 4540 6093
rect 4586 6047 4654 6093
rect 4700 6047 4768 6093
rect 4814 6047 4882 6093
rect 4928 6047 4996 6093
rect 5042 6047 5110 6093
rect 5156 6047 5224 6093
rect 5270 6047 5338 6093
rect 5384 6047 5452 6093
rect 5498 6047 5566 6093
rect 5612 6047 5680 6093
rect 5726 6047 5794 6093
rect 5840 6047 5908 6093
rect 5954 6047 6022 6093
rect 6068 6047 6136 6093
rect 6182 6047 6250 6093
rect 6296 6047 6364 6093
rect 6410 6047 6478 6093
rect 6524 6047 6592 6093
rect 6638 6047 6706 6093
rect 6752 6047 6820 6093
rect 6866 6047 6934 6093
rect 6980 6047 7048 6093
rect 7094 6047 7162 6093
rect 7208 6047 7276 6093
rect 7322 6047 7390 6093
rect 7436 6047 7504 6093
rect 7550 6047 7618 6093
rect 7664 6047 7732 6093
rect 7778 6047 7846 6093
rect 7892 6047 7960 6093
rect 8006 6047 8074 6093
rect 8120 6047 8188 6093
rect 8234 6047 8302 6093
rect 8348 6047 8416 6093
rect 8462 6047 8530 6093
rect 8576 6047 8644 6093
rect 8690 6047 8758 6093
rect 8804 6047 8872 6093
rect 8918 6047 8986 6093
rect 9032 6047 9100 6093
rect 9146 6047 9214 6093
rect 9260 6047 9328 6093
rect 9374 6047 9442 6093
rect 9488 6047 9556 6093
rect 9602 6047 9670 6093
rect 9716 6047 9784 6093
rect 9830 6047 9898 6093
rect 9944 6047 10012 6093
rect 10058 6047 10126 6093
rect 10172 6047 10240 6093
rect 10286 6047 10576 6093
rect 32 6028 10576 6047
rect 32 6025 10394 6028
rect 4998 5951 5088 6025
rect 4998 5905 5020 5951
rect 5066 5905 5088 5951
rect 4998 5827 5088 5905
rect 4998 5781 5020 5827
rect 5066 5781 5088 5827
rect 4998 5703 5088 5781
rect 10372 5982 10394 6025
rect 10440 5982 10508 6028
rect 10554 5982 10576 6028
rect 10372 5914 10576 5982
rect 10372 5868 10394 5914
rect 10440 5868 10508 5914
rect 10554 5868 10576 5914
rect 10372 5800 10576 5868
rect 10372 5754 10394 5800
rect 10440 5754 10508 5800
rect 10554 5754 10576 5800
rect 4998 5657 5020 5703
rect 5066 5657 5088 5703
rect 4998 5579 5088 5657
rect 10372 5686 10576 5754
rect 10372 5640 10394 5686
rect 10440 5640 10508 5686
rect 10554 5640 10576 5686
rect 4998 5533 5020 5579
rect 5066 5533 5088 5579
rect 4998 5455 5088 5533
rect 4998 5409 5020 5455
rect 5066 5409 5088 5455
rect 4998 5331 5088 5409
rect 4998 5285 5020 5331
rect 5066 5285 5088 5331
rect 4998 5207 5088 5285
rect 4998 5161 5020 5207
rect 5066 5161 5088 5207
rect 4998 5083 5088 5161
rect 4998 5037 5020 5083
rect 5066 5037 5088 5083
rect 4998 4959 5088 5037
rect 4998 4913 5020 4959
rect 5066 4913 5088 4959
rect 4998 4835 5088 4913
rect 4998 4789 5020 4835
rect 5066 4789 5088 4835
rect 4998 4711 5088 4789
rect 4998 4665 5020 4711
rect 5066 4665 5088 4711
rect 4998 4587 5088 4665
rect 4998 4541 5020 4587
rect 5066 4541 5088 4587
rect 4998 4463 5088 4541
rect 4998 4417 5020 4463
rect 5066 4417 5088 4463
rect 4998 4339 5088 4417
rect 4998 4293 5020 4339
rect 5066 4293 5088 4339
rect 4998 4215 5088 4293
rect 4998 4169 5020 4215
rect 5066 4169 5088 4215
rect 4998 4091 5088 4169
rect 4998 4045 5020 4091
rect 5066 4045 5088 4091
rect 4998 3967 5088 4045
rect 4998 3921 5020 3967
rect 5066 3921 5088 3967
rect 4998 3843 5088 3921
rect 4998 3797 5020 3843
rect 5066 3797 5088 3843
rect 4998 3719 5088 3797
rect 4998 3673 5020 3719
rect 5066 3673 5088 3719
rect 4998 3595 5088 3673
rect 4998 3549 5020 3595
rect 5066 3549 5088 3595
rect 4998 3471 5088 3549
rect 4998 3425 5020 3471
rect 5066 3425 5088 3471
rect 4998 3347 5088 3425
rect 4998 3301 5020 3347
rect 5066 3301 5088 3347
rect 4998 3223 5088 3301
rect 4998 3177 5020 3223
rect 5066 3177 5088 3223
rect 4998 3099 5088 3177
rect 4998 3053 5020 3099
rect 5066 3053 5088 3099
rect 4998 2975 5088 3053
rect 4998 2929 5020 2975
rect 5066 2929 5088 2975
rect 4998 2851 5088 2929
rect 4998 2805 5020 2851
rect 5066 2805 5088 2851
rect 4998 2727 5088 2805
rect 4998 2681 5020 2727
rect 5066 2681 5088 2727
rect 4998 2603 5088 2681
rect 4998 2557 5020 2603
rect 5066 2557 5088 2603
rect 4998 2479 5088 2557
rect 4998 2433 5020 2479
rect 5066 2433 5088 2479
rect 4998 2355 5088 2433
rect 4998 2309 5020 2355
rect 5066 2309 5088 2355
rect 4998 2231 5088 2309
rect 4998 2185 5020 2231
rect 5066 2185 5088 2231
rect 4998 2107 5088 2185
rect 4998 2061 5020 2107
rect 5066 2061 5088 2107
rect 4998 1983 5088 2061
rect 4998 1937 5020 1983
rect 5066 1937 5088 1983
rect 4998 1859 5088 1937
rect 4998 1813 5020 1859
rect 5066 1813 5088 1859
rect 4998 1735 5088 1813
rect 4998 1689 5020 1735
rect 5066 1689 5088 1735
rect 4998 1611 5088 1689
rect 4998 1565 5020 1611
rect 5066 1565 5088 1611
rect 4998 1487 5088 1565
rect 4998 1441 5020 1487
rect 5066 1441 5088 1487
rect 4998 1363 5088 1441
rect 4998 1317 5020 1363
rect 5066 1317 5088 1363
rect 4998 1239 5088 1317
rect 4998 1193 5020 1239
rect 5066 1193 5088 1239
rect 4998 1115 5088 1193
rect 4998 1069 5020 1115
rect 5066 1069 5088 1115
rect 4998 991 5088 1069
rect 4998 945 5020 991
rect 5066 945 5088 991
rect 4998 867 5088 945
rect 4998 821 5020 867
rect 5066 821 5088 867
rect 4998 743 5088 821
rect 4998 697 5020 743
rect 5066 697 5088 743
rect 4998 619 5088 697
rect 10372 5572 10576 5640
rect 10372 5526 10394 5572
rect 10440 5526 10508 5572
rect 10554 5526 10576 5572
rect 10372 5458 10576 5526
rect 10372 5412 10394 5458
rect 10440 5412 10508 5458
rect 10554 5412 10576 5458
rect 10372 5344 10576 5412
rect 10372 5298 10394 5344
rect 10440 5298 10508 5344
rect 10554 5298 10576 5344
rect 10372 5230 10576 5298
rect 10372 5184 10394 5230
rect 10440 5184 10508 5230
rect 10554 5184 10576 5230
rect 10372 5116 10576 5184
rect 10372 5070 10394 5116
rect 10440 5070 10508 5116
rect 10554 5070 10576 5116
rect 10372 5002 10576 5070
rect 10372 4956 10394 5002
rect 10440 4956 10508 5002
rect 10554 4956 10576 5002
rect 10372 4888 10576 4956
rect 10372 4842 10394 4888
rect 10440 4842 10508 4888
rect 10554 4842 10576 4888
rect 10372 4774 10576 4842
rect 10372 4728 10394 4774
rect 10440 4728 10508 4774
rect 10554 4728 10576 4774
rect 10372 4660 10576 4728
rect 10372 4614 10394 4660
rect 10440 4614 10508 4660
rect 10554 4614 10576 4660
rect 10372 4546 10576 4614
rect 10372 4500 10394 4546
rect 10440 4500 10508 4546
rect 10554 4500 10576 4546
rect 10372 4432 10576 4500
rect 10372 4386 10394 4432
rect 10440 4386 10508 4432
rect 10554 4386 10576 4432
rect 10372 4318 10576 4386
rect 10372 4272 10394 4318
rect 10440 4272 10508 4318
rect 10554 4272 10576 4318
rect 10372 4204 10576 4272
rect 10372 4158 10394 4204
rect 10440 4158 10508 4204
rect 10554 4158 10576 4204
rect 10372 4090 10576 4158
rect 10372 4044 10394 4090
rect 10440 4044 10508 4090
rect 10554 4044 10576 4090
rect 10372 3976 10576 4044
rect 10372 3930 10394 3976
rect 10440 3930 10508 3976
rect 10554 3930 10576 3976
rect 10372 3862 10576 3930
rect 10372 3816 10394 3862
rect 10440 3816 10508 3862
rect 10554 3816 10576 3862
rect 10372 3748 10576 3816
rect 10372 3702 10394 3748
rect 10440 3702 10508 3748
rect 10554 3702 10576 3748
rect 10372 3634 10576 3702
rect 10372 3588 10394 3634
rect 10440 3588 10508 3634
rect 10554 3588 10576 3634
rect 10372 3520 10576 3588
rect 10372 3474 10394 3520
rect 10440 3474 10508 3520
rect 10554 3474 10576 3520
rect 10372 3406 10576 3474
rect 10372 3360 10394 3406
rect 10440 3360 10508 3406
rect 10554 3360 10576 3406
rect 10372 3292 10576 3360
rect 10372 3246 10394 3292
rect 10440 3246 10508 3292
rect 10554 3246 10576 3292
rect 10372 3178 10576 3246
rect 10372 3132 10394 3178
rect 10440 3132 10508 3178
rect 10554 3132 10576 3178
rect 10372 3064 10576 3132
rect 10372 3018 10394 3064
rect 10440 3018 10508 3064
rect 10554 3018 10576 3064
rect 10372 2950 10576 3018
rect 10372 2904 10394 2950
rect 10440 2904 10508 2950
rect 10554 2904 10576 2950
rect 10372 2836 10576 2904
rect 10372 2790 10394 2836
rect 10440 2790 10508 2836
rect 10554 2790 10576 2836
rect 10372 2722 10576 2790
rect 10372 2676 10394 2722
rect 10440 2676 10508 2722
rect 10554 2676 10576 2722
rect 10372 2608 10576 2676
rect 10372 2562 10394 2608
rect 10440 2562 10508 2608
rect 10554 2562 10576 2608
rect 10372 2494 10576 2562
rect 10372 2448 10394 2494
rect 10440 2448 10508 2494
rect 10554 2448 10576 2494
rect 10372 2380 10576 2448
rect 10372 2334 10394 2380
rect 10440 2334 10508 2380
rect 10554 2334 10576 2380
rect 10372 2266 10576 2334
rect 10372 2220 10394 2266
rect 10440 2220 10508 2266
rect 10554 2220 10576 2266
rect 10372 2152 10576 2220
rect 10372 2106 10394 2152
rect 10440 2106 10508 2152
rect 10554 2106 10576 2152
rect 10372 2038 10576 2106
rect 10372 1992 10394 2038
rect 10440 1992 10508 2038
rect 10554 1992 10576 2038
rect 10372 1924 10576 1992
rect 10372 1878 10394 1924
rect 10440 1878 10508 1924
rect 10554 1878 10576 1924
rect 10372 1810 10576 1878
rect 10372 1764 10394 1810
rect 10440 1764 10508 1810
rect 10554 1764 10576 1810
rect 10372 1696 10576 1764
rect 10372 1650 10394 1696
rect 10440 1650 10508 1696
rect 10554 1650 10576 1696
rect 10372 1582 10576 1650
rect 10372 1536 10394 1582
rect 10440 1536 10508 1582
rect 10554 1536 10576 1582
rect 10372 1468 10576 1536
rect 10372 1422 10394 1468
rect 10440 1422 10508 1468
rect 10554 1422 10576 1468
rect 10372 1354 10576 1422
rect 10372 1308 10394 1354
rect 10440 1308 10508 1354
rect 10554 1308 10576 1354
rect 10372 1240 10576 1308
rect 10372 1194 10394 1240
rect 10440 1194 10508 1240
rect 10554 1194 10576 1240
rect 10372 1126 10576 1194
rect 10372 1080 10394 1126
rect 10440 1080 10508 1126
rect 10554 1080 10576 1126
rect 10372 1012 10576 1080
rect 10372 966 10394 1012
rect 10440 966 10508 1012
rect 10554 966 10576 1012
rect 10372 898 10576 966
rect 10372 852 10394 898
rect 10440 852 10508 898
rect 10554 852 10576 898
rect 10372 784 10576 852
rect 10372 738 10394 784
rect 10440 738 10508 784
rect 10554 738 10576 784
rect 10372 670 10576 738
rect 10372 624 10394 670
rect 10440 624 10508 670
rect 10554 624 10576 670
rect 4998 573 5020 619
rect 5066 573 5088 619
rect 4998 495 5088 573
rect 10372 556 10576 624
rect 4998 449 5020 495
rect 5066 449 5088 495
rect 4998 371 5088 449
rect 4998 325 5020 371
rect 5066 325 5088 371
rect 4998 247 5088 325
rect 4998 201 5020 247
rect 5066 236 5088 247
rect 10372 510 10394 556
rect 10440 510 10508 556
rect 10554 510 10576 556
rect 10372 442 10576 510
rect 10372 396 10394 442
rect 10440 396 10508 442
rect 10554 396 10576 442
rect 10372 328 10576 396
rect 10372 282 10394 328
rect 10440 282 10508 328
rect 10554 282 10576 328
rect 10372 236 10576 282
rect 5066 214 10576 236
rect 5066 201 5354 214
rect 4998 168 5354 201
rect 5400 168 5468 214
rect 5514 168 5582 214
rect 5628 168 5696 214
rect 5742 168 5810 214
rect 5856 168 5924 214
rect 5970 168 6038 214
rect 6084 168 6152 214
rect 6198 168 6266 214
rect 6312 168 6380 214
rect 6426 168 6494 214
rect 6540 168 6608 214
rect 6654 168 6722 214
rect 6768 168 6836 214
rect 6882 168 6950 214
rect 6996 168 7064 214
rect 7110 168 7178 214
rect 7224 168 7292 214
rect 7338 168 7406 214
rect 7452 168 7520 214
rect 7566 168 7634 214
rect 7680 168 7748 214
rect 7794 168 7862 214
rect 7908 168 7976 214
rect 8022 168 8090 214
rect 8136 168 8204 214
rect 8250 168 8318 214
rect 8364 168 8432 214
rect 8478 168 8546 214
rect 8592 168 8660 214
rect 8706 168 8774 214
rect 8820 168 8888 214
rect 8934 168 9002 214
rect 9048 168 9116 214
rect 9162 168 9230 214
rect 9276 168 9344 214
rect 9390 168 9458 214
rect 9504 168 9572 214
rect 9618 168 9686 214
rect 9732 168 9800 214
rect 9846 168 9914 214
rect 9960 168 10028 214
rect 10074 168 10142 214
rect 10188 168 10256 214
rect 10302 168 10394 214
rect 10440 168 10508 214
rect 10554 168 10576 214
rect 4998 123 10576 168
rect 4998 77 5020 123
rect 5066 100 10576 123
rect 5066 77 5354 100
rect 4998 54 5354 77
rect 5400 54 5468 100
rect 5514 54 5582 100
rect 5628 54 5696 100
rect 5742 54 5810 100
rect 5856 54 5924 100
rect 5970 54 6038 100
rect 6084 54 6152 100
rect 6198 54 6266 100
rect 6312 54 6380 100
rect 6426 54 6494 100
rect 6540 54 6608 100
rect 6654 54 6722 100
rect 6768 54 6836 100
rect 6882 54 6950 100
rect 6996 54 7064 100
rect 7110 54 7178 100
rect 7224 54 7292 100
rect 7338 54 7406 100
rect 7452 54 7520 100
rect 7566 54 7634 100
rect 7680 54 7748 100
rect 7794 54 7862 100
rect 7908 54 7976 100
rect 8022 54 8090 100
rect 8136 54 8204 100
rect 8250 54 8318 100
rect 8364 54 8432 100
rect 8478 54 8546 100
rect 8592 54 8660 100
rect 8706 54 8774 100
rect 8820 54 8888 100
rect 8934 54 9002 100
rect 9048 54 9116 100
rect 9162 54 9230 100
rect 9276 54 9344 100
rect 9390 54 9458 100
rect 9504 54 9572 100
rect 9618 54 9686 100
rect 9732 54 9800 100
rect 9846 54 9914 100
rect 9960 54 10028 100
rect 10074 54 10142 100
rect 10188 54 10256 100
rect 10302 54 10394 100
rect 10440 54 10508 100
rect 10554 54 10576 100
rect 4998 32 10576 54
<< psubdiffcont >>
rect 54 12252 100 12298
rect 168 12252 214 12298
rect 322 12252 368 12298
rect 436 12252 482 12298
rect 550 12252 596 12298
rect 664 12252 710 12298
rect 778 12252 824 12298
rect 892 12252 938 12298
rect 1006 12252 1052 12298
rect 1120 12252 1166 12298
rect 1234 12252 1280 12298
rect 1348 12252 1394 12298
rect 1462 12252 1508 12298
rect 1576 12252 1622 12298
rect 1690 12252 1736 12298
rect 1804 12252 1850 12298
rect 1918 12252 1964 12298
rect 2032 12252 2078 12298
rect 2146 12252 2192 12298
rect 2260 12252 2306 12298
rect 2374 12252 2420 12298
rect 2488 12252 2534 12298
rect 2602 12252 2648 12298
rect 2716 12252 2762 12298
rect 2830 12252 2876 12298
rect 2944 12252 2990 12298
rect 3058 12252 3104 12298
rect 3172 12252 3218 12298
rect 3286 12252 3332 12298
rect 3400 12252 3446 12298
rect 3514 12252 3560 12298
rect 3628 12252 3674 12298
rect 3742 12252 3788 12298
rect 3856 12252 3902 12298
rect 3970 12252 4016 12298
rect 4084 12252 4130 12298
rect 4198 12252 4244 12298
rect 4312 12252 4358 12298
rect 4426 12252 4472 12298
rect 4540 12252 4586 12298
rect 4654 12252 4700 12298
rect 4768 12252 4814 12298
rect 4882 12252 4928 12298
rect 4996 12252 5042 12298
rect 5110 12252 5156 12298
rect 5224 12252 5270 12298
rect 5338 12252 5384 12298
rect 5452 12252 5498 12298
rect 5566 12252 5612 12298
rect 5680 12252 5726 12298
rect 5794 12252 5840 12298
rect 5908 12252 5954 12298
rect 6022 12252 6068 12298
rect 6136 12252 6182 12298
rect 6250 12252 6296 12298
rect 6364 12252 6410 12298
rect 6478 12252 6524 12298
rect 6592 12252 6638 12298
rect 6706 12252 6752 12298
rect 6820 12252 6866 12298
rect 6934 12252 6980 12298
rect 7048 12252 7094 12298
rect 7162 12252 7208 12298
rect 7276 12252 7322 12298
rect 7390 12252 7436 12298
rect 7504 12252 7550 12298
rect 7618 12252 7664 12298
rect 7732 12252 7778 12298
rect 7846 12252 7892 12298
rect 7960 12252 8006 12298
rect 8074 12252 8120 12298
rect 8188 12252 8234 12298
rect 8302 12252 8348 12298
rect 8416 12252 8462 12298
rect 8530 12252 8576 12298
rect 8644 12252 8690 12298
rect 8758 12252 8804 12298
rect 8872 12252 8918 12298
rect 8986 12252 9032 12298
rect 9100 12252 9146 12298
rect 9214 12252 9260 12298
rect 9328 12252 9374 12298
rect 9442 12252 9488 12298
rect 9556 12252 9602 12298
rect 9670 12252 9716 12298
rect 9784 12252 9830 12298
rect 9898 12252 9944 12298
rect 10012 12252 10058 12298
rect 10126 12252 10172 12298
rect 10240 12252 10286 12298
rect 10394 12252 10440 12298
rect 10508 12252 10554 12298
rect 54 12138 100 12184
rect 168 12138 214 12184
rect 322 12138 368 12184
rect 436 12138 482 12184
rect 550 12138 596 12184
rect 664 12138 710 12184
rect 778 12138 824 12184
rect 892 12138 938 12184
rect 1006 12138 1052 12184
rect 1120 12138 1166 12184
rect 1234 12138 1280 12184
rect 1348 12138 1394 12184
rect 1462 12138 1508 12184
rect 1576 12138 1622 12184
rect 1690 12138 1736 12184
rect 1804 12138 1850 12184
rect 1918 12138 1964 12184
rect 2032 12138 2078 12184
rect 2146 12138 2192 12184
rect 2260 12138 2306 12184
rect 2374 12138 2420 12184
rect 2488 12138 2534 12184
rect 2602 12138 2648 12184
rect 2716 12138 2762 12184
rect 2830 12138 2876 12184
rect 2944 12138 2990 12184
rect 3058 12138 3104 12184
rect 3172 12138 3218 12184
rect 3286 12138 3332 12184
rect 3400 12138 3446 12184
rect 3514 12138 3560 12184
rect 3628 12138 3674 12184
rect 3742 12138 3788 12184
rect 3856 12138 3902 12184
rect 3970 12138 4016 12184
rect 4084 12138 4130 12184
rect 4198 12138 4244 12184
rect 4312 12138 4358 12184
rect 4426 12138 4472 12184
rect 4540 12138 4586 12184
rect 4654 12138 4700 12184
rect 4768 12138 4814 12184
rect 4882 12138 4928 12184
rect 4996 12138 5042 12184
rect 5110 12138 5156 12184
rect 5224 12138 5270 12184
rect 5338 12138 5384 12184
rect 5452 12138 5498 12184
rect 5566 12138 5612 12184
rect 5680 12138 5726 12184
rect 5794 12138 5840 12184
rect 5908 12138 5954 12184
rect 6022 12138 6068 12184
rect 6136 12138 6182 12184
rect 6250 12138 6296 12184
rect 6364 12138 6410 12184
rect 6478 12138 6524 12184
rect 6592 12138 6638 12184
rect 6706 12138 6752 12184
rect 6820 12138 6866 12184
rect 6934 12138 6980 12184
rect 7048 12138 7094 12184
rect 7162 12138 7208 12184
rect 7276 12138 7322 12184
rect 7390 12138 7436 12184
rect 7504 12138 7550 12184
rect 7618 12138 7664 12184
rect 7732 12138 7778 12184
rect 7846 12138 7892 12184
rect 7960 12138 8006 12184
rect 8074 12138 8120 12184
rect 8188 12138 8234 12184
rect 8302 12138 8348 12184
rect 8416 12138 8462 12184
rect 8530 12138 8576 12184
rect 8644 12138 8690 12184
rect 8758 12138 8804 12184
rect 8872 12138 8918 12184
rect 8986 12138 9032 12184
rect 9100 12138 9146 12184
rect 9214 12138 9260 12184
rect 9328 12138 9374 12184
rect 9442 12138 9488 12184
rect 9556 12138 9602 12184
rect 9670 12138 9716 12184
rect 9784 12138 9830 12184
rect 9898 12138 9944 12184
rect 10012 12138 10058 12184
rect 10126 12138 10172 12184
rect 10240 12138 10286 12184
rect 10394 12138 10440 12184
rect 10508 12138 10554 12184
rect 54 12024 100 12070
rect 168 12024 214 12070
rect 10394 12024 10440 12070
rect 10508 12024 10554 12070
rect 10394 11910 10440 11956
rect 10508 11910 10554 11956
rect 10394 11796 10440 11842
rect 10508 11796 10554 11842
rect 10394 11682 10440 11728
rect 10508 11682 10554 11728
rect 54 11454 100 11500
rect 168 11454 214 11500
rect 54 11340 100 11386
rect 168 11340 214 11386
rect 54 11226 100 11272
rect 168 11226 214 11272
rect 54 11112 100 11158
rect 168 11112 214 11158
rect 54 10998 100 11044
rect 168 10998 214 11044
rect 54 10884 100 10930
rect 168 10884 214 10930
rect 54 10770 100 10816
rect 168 10770 214 10816
rect 54 10656 100 10702
rect 168 10656 214 10702
rect 54 10542 100 10588
rect 168 10542 214 10588
rect 54 10428 100 10474
rect 168 10428 214 10474
rect 54 10314 100 10360
rect 168 10314 214 10360
rect 54 10200 100 10246
rect 168 10200 214 10246
rect 54 10086 100 10132
rect 168 10086 214 10132
rect 54 9972 100 10018
rect 168 9972 214 10018
rect 54 9858 100 9904
rect 168 9858 214 9904
rect 54 9744 100 9790
rect 168 9744 214 9790
rect 54 9630 100 9676
rect 168 9630 214 9676
rect 54 9516 100 9562
rect 168 9516 214 9562
rect 54 9402 100 9448
rect 168 9402 214 9448
rect 54 9288 100 9334
rect 168 9288 214 9334
rect 54 9174 100 9220
rect 168 9174 214 9220
rect 54 9060 100 9106
rect 168 9060 214 9106
rect 54 8946 100 8992
rect 168 8946 214 8992
rect 54 8832 100 8878
rect 168 8832 214 8878
rect 54 8718 100 8764
rect 168 8718 214 8764
rect 54 8604 100 8650
rect 168 8604 214 8650
rect 54 8490 100 8536
rect 168 8490 214 8536
rect 54 8376 100 8422
rect 168 8376 214 8422
rect 54 8262 100 8308
rect 168 8262 214 8308
rect 54 8148 100 8194
rect 168 8148 214 8194
rect 54 8034 100 8080
rect 168 8034 214 8080
rect 54 7920 100 7966
rect 168 7920 214 7966
rect 54 7806 100 7852
rect 168 7806 214 7852
rect 54 7692 100 7738
rect 168 7692 214 7738
rect 54 7578 100 7624
rect 168 7578 214 7624
rect 54 7464 100 7510
rect 168 7464 214 7510
rect 54 7350 100 7396
rect 168 7350 214 7396
rect 54 7236 100 7282
rect 168 7236 214 7282
rect 54 7122 100 7168
rect 168 7122 214 7168
rect 54 7008 100 7054
rect 168 7008 214 7054
rect 54 6894 100 6940
rect 168 6894 214 6940
rect 54 6780 100 6826
rect 168 6780 214 6826
rect 54 6666 100 6712
rect 168 6666 214 6712
rect 10394 11568 10440 11614
rect 10508 11568 10554 11614
rect 10394 11454 10440 11500
rect 10508 11454 10554 11500
rect 10394 11340 10440 11386
rect 10508 11340 10554 11386
rect 10394 11226 10440 11272
rect 10508 11226 10554 11272
rect 10394 11112 10440 11158
rect 10508 11112 10554 11158
rect 10394 10998 10440 11044
rect 10508 10998 10554 11044
rect 10394 10884 10440 10930
rect 10508 10884 10554 10930
rect 10394 10770 10440 10816
rect 10508 10770 10554 10816
rect 10394 10656 10440 10702
rect 10508 10656 10554 10702
rect 10394 10542 10440 10588
rect 10508 10542 10554 10588
rect 10394 10428 10440 10474
rect 10508 10428 10554 10474
rect 10394 10314 10440 10360
rect 10508 10314 10554 10360
rect 10394 10200 10440 10246
rect 10508 10200 10554 10246
rect 10394 10086 10440 10132
rect 10508 10086 10554 10132
rect 10394 9972 10440 10018
rect 10508 9972 10554 10018
rect 10394 9858 10440 9904
rect 10508 9858 10554 9904
rect 10394 9744 10440 9790
rect 10508 9744 10554 9790
rect 10394 9630 10440 9676
rect 10508 9630 10554 9676
rect 10394 9516 10440 9562
rect 10508 9516 10554 9562
rect 10394 9402 10440 9448
rect 10508 9402 10554 9448
rect 10394 9288 10440 9334
rect 10508 9288 10554 9334
rect 10394 9174 10440 9220
rect 10508 9174 10554 9220
rect 10394 9060 10440 9106
rect 10508 9060 10554 9106
rect 10394 8946 10440 8992
rect 10508 8946 10554 8992
rect 10394 8832 10440 8878
rect 10508 8832 10554 8878
rect 10394 8718 10440 8764
rect 10508 8718 10554 8764
rect 10394 8604 10440 8650
rect 10508 8604 10554 8650
rect 10394 8490 10440 8536
rect 10508 8490 10554 8536
rect 10394 8376 10440 8422
rect 10508 8376 10554 8422
rect 10394 8262 10440 8308
rect 10508 8262 10554 8308
rect 10394 8148 10440 8194
rect 10508 8148 10554 8194
rect 10394 8034 10440 8080
rect 10508 8034 10554 8080
rect 10394 7920 10440 7966
rect 10508 7920 10554 7966
rect 10394 7806 10440 7852
rect 10508 7806 10554 7852
rect 10394 7692 10440 7738
rect 10508 7692 10554 7738
rect 10394 7578 10440 7624
rect 10508 7578 10554 7624
rect 10394 7464 10440 7510
rect 10508 7464 10554 7510
rect 10394 7350 10440 7396
rect 10508 7350 10554 7396
rect 10394 7236 10440 7282
rect 10508 7236 10554 7282
rect 10394 7122 10440 7168
rect 10508 7122 10554 7168
rect 10394 7008 10440 7054
rect 10508 7008 10554 7054
rect 10394 6894 10440 6940
rect 10508 6894 10554 6940
rect 10394 6780 10440 6826
rect 10508 6780 10554 6826
rect 10394 6666 10440 6712
rect 10508 6666 10554 6712
rect 54 6552 100 6598
rect 168 6552 214 6598
rect 10394 6552 10440 6598
rect 10508 6552 10554 6598
rect 54 6438 100 6484
rect 168 6438 214 6484
rect 54 6324 100 6370
rect 168 6324 214 6370
rect 10394 6438 10440 6484
rect 10508 6438 10554 6484
rect 10394 6324 10440 6370
rect 10508 6324 10554 6370
rect 10394 6210 10440 6256
rect 10508 6210 10554 6256
rect 322 6161 368 6207
rect 436 6161 482 6207
rect 550 6161 596 6207
rect 664 6161 710 6207
rect 778 6161 824 6207
rect 892 6161 938 6207
rect 1006 6161 1052 6207
rect 1120 6161 1166 6207
rect 1234 6161 1280 6207
rect 1348 6161 1394 6207
rect 1462 6161 1508 6207
rect 1576 6161 1622 6207
rect 1690 6161 1736 6207
rect 1804 6161 1850 6207
rect 1918 6161 1964 6207
rect 2032 6161 2078 6207
rect 2146 6161 2192 6207
rect 2260 6161 2306 6207
rect 2374 6161 2420 6207
rect 2488 6161 2534 6207
rect 2602 6161 2648 6207
rect 2716 6161 2762 6207
rect 2830 6161 2876 6207
rect 2944 6161 2990 6207
rect 3058 6161 3104 6207
rect 3172 6161 3218 6207
rect 3286 6161 3332 6207
rect 3400 6161 3446 6207
rect 3514 6161 3560 6207
rect 3628 6161 3674 6207
rect 3742 6161 3788 6207
rect 3856 6161 3902 6207
rect 3970 6161 4016 6207
rect 4084 6161 4130 6207
rect 4198 6161 4244 6207
rect 4312 6161 4358 6207
rect 4426 6161 4472 6207
rect 4540 6161 4586 6207
rect 4654 6161 4700 6207
rect 4768 6161 4814 6207
rect 4882 6161 4928 6207
rect 4996 6161 5042 6207
rect 5110 6161 5156 6207
rect 5224 6161 5270 6207
rect 5338 6161 5384 6207
rect 5452 6161 5498 6207
rect 5566 6161 5612 6207
rect 5680 6161 5726 6207
rect 5794 6161 5840 6207
rect 5908 6161 5954 6207
rect 6022 6161 6068 6207
rect 6136 6161 6182 6207
rect 6250 6161 6296 6207
rect 6364 6161 6410 6207
rect 6478 6161 6524 6207
rect 6592 6161 6638 6207
rect 6706 6161 6752 6207
rect 6820 6161 6866 6207
rect 6934 6161 6980 6207
rect 7048 6161 7094 6207
rect 7162 6161 7208 6207
rect 7276 6161 7322 6207
rect 7390 6161 7436 6207
rect 7504 6161 7550 6207
rect 7618 6161 7664 6207
rect 7732 6161 7778 6207
rect 7846 6161 7892 6207
rect 7960 6161 8006 6207
rect 8074 6161 8120 6207
rect 8188 6161 8234 6207
rect 8302 6161 8348 6207
rect 8416 6161 8462 6207
rect 8530 6161 8576 6207
rect 8644 6161 8690 6207
rect 8758 6161 8804 6207
rect 8872 6161 8918 6207
rect 8986 6161 9032 6207
rect 9100 6161 9146 6207
rect 9214 6161 9260 6207
rect 9328 6161 9374 6207
rect 9442 6161 9488 6207
rect 9556 6161 9602 6207
rect 9670 6161 9716 6207
rect 9784 6161 9830 6207
rect 9898 6161 9944 6207
rect 10012 6161 10058 6207
rect 10126 6161 10172 6207
rect 10240 6161 10286 6207
rect 10394 6096 10440 6142
rect 10508 6096 10554 6142
rect 322 6047 368 6093
rect 436 6047 482 6093
rect 550 6047 596 6093
rect 664 6047 710 6093
rect 778 6047 824 6093
rect 892 6047 938 6093
rect 1006 6047 1052 6093
rect 1120 6047 1166 6093
rect 1234 6047 1280 6093
rect 1348 6047 1394 6093
rect 1462 6047 1508 6093
rect 1576 6047 1622 6093
rect 1690 6047 1736 6093
rect 1804 6047 1850 6093
rect 1918 6047 1964 6093
rect 2032 6047 2078 6093
rect 2146 6047 2192 6093
rect 2260 6047 2306 6093
rect 2374 6047 2420 6093
rect 2488 6047 2534 6093
rect 2602 6047 2648 6093
rect 2716 6047 2762 6093
rect 2830 6047 2876 6093
rect 2944 6047 2990 6093
rect 3058 6047 3104 6093
rect 3172 6047 3218 6093
rect 3286 6047 3332 6093
rect 3400 6047 3446 6093
rect 3514 6047 3560 6093
rect 3628 6047 3674 6093
rect 3742 6047 3788 6093
rect 3856 6047 3902 6093
rect 3970 6047 4016 6093
rect 4084 6047 4130 6093
rect 4198 6047 4244 6093
rect 4312 6047 4358 6093
rect 4426 6047 4472 6093
rect 4540 6047 4586 6093
rect 4654 6047 4700 6093
rect 4768 6047 4814 6093
rect 4882 6047 4928 6093
rect 4996 6047 5042 6093
rect 5110 6047 5156 6093
rect 5224 6047 5270 6093
rect 5338 6047 5384 6093
rect 5452 6047 5498 6093
rect 5566 6047 5612 6093
rect 5680 6047 5726 6093
rect 5794 6047 5840 6093
rect 5908 6047 5954 6093
rect 6022 6047 6068 6093
rect 6136 6047 6182 6093
rect 6250 6047 6296 6093
rect 6364 6047 6410 6093
rect 6478 6047 6524 6093
rect 6592 6047 6638 6093
rect 6706 6047 6752 6093
rect 6820 6047 6866 6093
rect 6934 6047 6980 6093
rect 7048 6047 7094 6093
rect 7162 6047 7208 6093
rect 7276 6047 7322 6093
rect 7390 6047 7436 6093
rect 7504 6047 7550 6093
rect 7618 6047 7664 6093
rect 7732 6047 7778 6093
rect 7846 6047 7892 6093
rect 7960 6047 8006 6093
rect 8074 6047 8120 6093
rect 8188 6047 8234 6093
rect 8302 6047 8348 6093
rect 8416 6047 8462 6093
rect 8530 6047 8576 6093
rect 8644 6047 8690 6093
rect 8758 6047 8804 6093
rect 8872 6047 8918 6093
rect 8986 6047 9032 6093
rect 9100 6047 9146 6093
rect 9214 6047 9260 6093
rect 9328 6047 9374 6093
rect 9442 6047 9488 6093
rect 9556 6047 9602 6093
rect 9670 6047 9716 6093
rect 9784 6047 9830 6093
rect 9898 6047 9944 6093
rect 10012 6047 10058 6093
rect 10126 6047 10172 6093
rect 10240 6047 10286 6093
rect 5020 5905 5066 5951
rect 5020 5781 5066 5827
rect 10394 5982 10440 6028
rect 10508 5982 10554 6028
rect 10394 5868 10440 5914
rect 10508 5868 10554 5914
rect 10394 5754 10440 5800
rect 10508 5754 10554 5800
rect 5020 5657 5066 5703
rect 10394 5640 10440 5686
rect 10508 5640 10554 5686
rect 5020 5533 5066 5579
rect 5020 5409 5066 5455
rect 5020 5285 5066 5331
rect 5020 5161 5066 5207
rect 5020 5037 5066 5083
rect 5020 4913 5066 4959
rect 5020 4789 5066 4835
rect 5020 4665 5066 4711
rect 5020 4541 5066 4587
rect 5020 4417 5066 4463
rect 5020 4293 5066 4339
rect 5020 4169 5066 4215
rect 5020 4045 5066 4091
rect 5020 3921 5066 3967
rect 5020 3797 5066 3843
rect 5020 3673 5066 3719
rect 5020 3549 5066 3595
rect 5020 3425 5066 3471
rect 5020 3301 5066 3347
rect 5020 3177 5066 3223
rect 5020 3053 5066 3099
rect 5020 2929 5066 2975
rect 5020 2805 5066 2851
rect 5020 2681 5066 2727
rect 5020 2557 5066 2603
rect 5020 2433 5066 2479
rect 5020 2309 5066 2355
rect 5020 2185 5066 2231
rect 5020 2061 5066 2107
rect 5020 1937 5066 1983
rect 5020 1813 5066 1859
rect 5020 1689 5066 1735
rect 5020 1565 5066 1611
rect 5020 1441 5066 1487
rect 5020 1317 5066 1363
rect 5020 1193 5066 1239
rect 5020 1069 5066 1115
rect 5020 945 5066 991
rect 5020 821 5066 867
rect 5020 697 5066 743
rect 10394 5526 10440 5572
rect 10508 5526 10554 5572
rect 10394 5412 10440 5458
rect 10508 5412 10554 5458
rect 10394 5298 10440 5344
rect 10508 5298 10554 5344
rect 10394 5184 10440 5230
rect 10508 5184 10554 5230
rect 10394 5070 10440 5116
rect 10508 5070 10554 5116
rect 10394 4956 10440 5002
rect 10508 4956 10554 5002
rect 10394 4842 10440 4888
rect 10508 4842 10554 4888
rect 10394 4728 10440 4774
rect 10508 4728 10554 4774
rect 10394 4614 10440 4660
rect 10508 4614 10554 4660
rect 10394 4500 10440 4546
rect 10508 4500 10554 4546
rect 10394 4386 10440 4432
rect 10508 4386 10554 4432
rect 10394 4272 10440 4318
rect 10508 4272 10554 4318
rect 10394 4158 10440 4204
rect 10508 4158 10554 4204
rect 10394 4044 10440 4090
rect 10508 4044 10554 4090
rect 10394 3930 10440 3976
rect 10508 3930 10554 3976
rect 10394 3816 10440 3862
rect 10508 3816 10554 3862
rect 10394 3702 10440 3748
rect 10508 3702 10554 3748
rect 10394 3588 10440 3634
rect 10508 3588 10554 3634
rect 10394 3474 10440 3520
rect 10508 3474 10554 3520
rect 10394 3360 10440 3406
rect 10508 3360 10554 3406
rect 10394 3246 10440 3292
rect 10508 3246 10554 3292
rect 10394 3132 10440 3178
rect 10508 3132 10554 3178
rect 10394 3018 10440 3064
rect 10508 3018 10554 3064
rect 10394 2904 10440 2950
rect 10508 2904 10554 2950
rect 10394 2790 10440 2836
rect 10508 2790 10554 2836
rect 10394 2676 10440 2722
rect 10508 2676 10554 2722
rect 10394 2562 10440 2608
rect 10508 2562 10554 2608
rect 10394 2448 10440 2494
rect 10508 2448 10554 2494
rect 10394 2334 10440 2380
rect 10508 2334 10554 2380
rect 10394 2220 10440 2266
rect 10508 2220 10554 2266
rect 10394 2106 10440 2152
rect 10508 2106 10554 2152
rect 10394 1992 10440 2038
rect 10508 1992 10554 2038
rect 10394 1878 10440 1924
rect 10508 1878 10554 1924
rect 10394 1764 10440 1810
rect 10508 1764 10554 1810
rect 10394 1650 10440 1696
rect 10508 1650 10554 1696
rect 10394 1536 10440 1582
rect 10508 1536 10554 1582
rect 10394 1422 10440 1468
rect 10508 1422 10554 1468
rect 10394 1308 10440 1354
rect 10508 1308 10554 1354
rect 10394 1194 10440 1240
rect 10508 1194 10554 1240
rect 10394 1080 10440 1126
rect 10508 1080 10554 1126
rect 10394 966 10440 1012
rect 10508 966 10554 1012
rect 10394 852 10440 898
rect 10508 852 10554 898
rect 10394 738 10440 784
rect 10508 738 10554 784
rect 10394 624 10440 670
rect 10508 624 10554 670
rect 5020 573 5066 619
rect 5020 449 5066 495
rect 5020 325 5066 371
rect 5020 201 5066 247
rect 10394 510 10440 556
rect 10508 510 10554 556
rect 10394 396 10440 442
rect 10508 396 10554 442
rect 10394 282 10440 328
rect 10508 282 10554 328
rect 5354 168 5400 214
rect 5468 168 5514 214
rect 5582 168 5628 214
rect 5696 168 5742 214
rect 5810 168 5856 214
rect 5924 168 5970 214
rect 6038 168 6084 214
rect 6152 168 6198 214
rect 6266 168 6312 214
rect 6380 168 6426 214
rect 6494 168 6540 214
rect 6608 168 6654 214
rect 6722 168 6768 214
rect 6836 168 6882 214
rect 6950 168 6996 214
rect 7064 168 7110 214
rect 7178 168 7224 214
rect 7292 168 7338 214
rect 7406 168 7452 214
rect 7520 168 7566 214
rect 7634 168 7680 214
rect 7748 168 7794 214
rect 7862 168 7908 214
rect 7976 168 8022 214
rect 8090 168 8136 214
rect 8204 168 8250 214
rect 8318 168 8364 214
rect 8432 168 8478 214
rect 8546 168 8592 214
rect 8660 168 8706 214
rect 8774 168 8820 214
rect 8888 168 8934 214
rect 9002 168 9048 214
rect 9116 168 9162 214
rect 9230 168 9276 214
rect 9344 168 9390 214
rect 9458 168 9504 214
rect 9572 168 9618 214
rect 9686 168 9732 214
rect 9800 168 9846 214
rect 9914 168 9960 214
rect 10028 168 10074 214
rect 10142 168 10188 214
rect 10256 168 10302 214
rect 10394 168 10440 214
rect 10508 168 10554 214
rect 5020 77 5066 123
rect 5354 54 5400 100
rect 5468 54 5514 100
rect 5582 54 5628 100
rect 5696 54 5742 100
rect 5810 54 5856 100
rect 5924 54 5970 100
rect 6038 54 6084 100
rect 6152 54 6198 100
rect 6266 54 6312 100
rect 6380 54 6426 100
rect 6494 54 6540 100
rect 6608 54 6654 100
rect 6722 54 6768 100
rect 6836 54 6882 100
rect 6950 54 6996 100
rect 7064 54 7110 100
rect 7178 54 7224 100
rect 7292 54 7338 100
rect 7406 54 7452 100
rect 7520 54 7566 100
rect 7634 54 7680 100
rect 7748 54 7794 100
rect 7862 54 7908 100
rect 7976 54 8022 100
rect 8090 54 8136 100
rect 8204 54 8250 100
rect 8318 54 8364 100
rect 8432 54 8478 100
rect 8546 54 8592 100
rect 8660 54 8706 100
rect 8774 54 8820 100
rect 8888 54 8934 100
rect 9002 54 9048 100
rect 9116 54 9162 100
rect 9230 54 9276 100
rect 9344 54 9390 100
rect 9458 54 9504 100
rect 9572 54 9618 100
rect 9686 54 9732 100
rect 9800 54 9846 100
rect 9914 54 9960 100
rect 10028 54 10074 100
rect 10142 54 10188 100
rect 10256 54 10302 100
rect 10394 54 10440 100
rect 10508 54 10554 100
<< mvnmoscap >>
rect 647 6633 2647 11633
rect 3083 6633 5083 11633
rect 5519 6633 7519 11633
rect 7955 6633 9955 11633
rect 5519 621 7519 5621
rect 7955 621 9955 5621
<< polysilicon >>
rect 647 11712 2647 11725
rect 647 11666 700 11712
rect 2594 11666 2647 11712
rect 647 11633 2647 11666
rect 3083 11712 5083 11725
rect 3083 11666 3136 11712
rect 5030 11666 5083 11712
rect 3083 11633 5083 11666
rect 5519 11712 7519 11725
rect 5519 11666 5572 11712
rect 7466 11666 7519 11712
rect 5519 11633 7519 11666
rect 7955 11712 9955 11725
rect 7955 11666 8008 11712
rect 9902 11666 9955 11712
rect 7955 11633 9955 11666
rect 647 6600 2647 6633
rect 647 6554 700 6600
rect 2594 6554 2647 6600
rect 647 6541 2647 6554
rect 3083 6600 5083 6633
rect 3083 6554 3136 6600
rect 5030 6554 5083 6600
rect 3083 6541 5083 6554
rect 5519 6600 7519 6633
rect 5519 6554 5572 6600
rect 7466 6554 7519 6600
rect 5519 6541 7519 6554
rect 7955 6600 9955 6633
rect 7955 6554 8008 6600
rect 9902 6554 9955 6600
rect 7955 6541 9955 6554
rect 5519 5700 7519 5713
rect 5519 5654 5572 5700
rect 7466 5654 7519 5700
rect 5519 5621 7519 5654
rect 7955 5700 9955 5713
rect 7955 5654 8008 5700
rect 9902 5654 9955 5700
rect 7955 5621 9955 5654
rect 5519 588 7519 621
rect 5519 542 5572 588
rect 7466 542 7519 588
rect 5519 529 7519 542
rect 7955 588 9955 621
rect 7955 542 8008 588
rect 9902 542 9955 588
rect 7955 529 9955 542
<< polycontact >>
rect 700 11666 2594 11712
rect 3136 11666 5030 11712
rect 5572 11666 7466 11712
rect 8008 11666 9902 11712
rect 700 6554 2594 6600
rect 3136 6554 5030 6600
rect 5572 6554 7466 6600
rect 8008 6554 9902 6600
rect 5572 5654 7466 5700
rect 8008 5654 9902 5700
rect 5572 542 7466 588
rect 8008 542 9902 588
<< metal1 >>
rect 43 12298 10565 12310
rect 43 12252 54 12298
rect 100 12252 168 12298
rect 214 12252 322 12298
rect 368 12252 436 12298
rect 482 12252 550 12298
rect 596 12252 664 12298
rect 710 12252 778 12298
rect 824 12252 892 12298
rect 938 12252 1006 12298
rect 1052 12252 1120 12298
rect 1166 12252 1234 12298
rect 1280 12252 1348 12298
rect 1394 12252 1462 12298
rect 1508 12252 1576 12298
rect 1622 12252 1690 12298
rect 1736 12252 1804 12298
rect 1850 12252 1918 12298
rect 1964 12252 2032 12298
rect 2078 12252 2146 12298
rect 2192 12252 2260 12298
rect 2306 12252 2374 12298
rect 2420 12252 2488 12298
rect 2534 12252 2602 12298
rect 2648 12252 2716 12298
rect 2762 12252 2830 12298
rect 2876 12252 2944 12298
rect 2990 12252 3058 12298
rect 3104 12252 3172 12298
rect 3218 12252 3286 12298
rect 3332 12252 3400 12298
rect 3446 12252 3514 12298
rect 3560 12252 3628 12298
rect 3674 12252 3742 12298
rect 3788 12252 3856 12298
rect 3902 12252 3970 12298
rect 4016 12252 4084 12298
rect 4130 12252 4198 12298
rect 4244 12252 4312 12298
rect 4358 12252 4426 12298
rect 4472 12252 4540 12298
rect 4586 12252 4654 12298
rect 4700 12252 4768 12298
rect 4814 12252 4882 12298
rect 4928 12252 4996 12298
rect 5042 12252 5110 12298
rect 5156 12252 5224 12298
rect 5270 12252 5338 12298
rect 5384 12252 5452 12298
rect 5498 12252 5566 12298
rect 5612 12252 5680 12298
rect 5726 12252 5794 12298
rect 5840 12252 5908 12298
rect 5954 12252 6022 12298
rect 6068 12252 6136 12298
rect 6182 12252 6250 12298
rect 6296 12252 6364 12298
rect 6410 12252 6478 12298
rect 6524 12252 6592 12298
rect 6638 12252 6706 12298
rect 6752 12252 6820 12298
rect 6866 12252 6934 12298
rect 6980 12252 7048 12298
rect 7094 12252 7162 12298
rect 7208 12252 7276 12298
rect 7322 12252 7390 12298
rect 7436 12252 7504 12298
rect 7550 12252 7618 12298
rect 7664 12252 7732 12298
rect 7778 12252 7846 12298
rect 7892 12252 7960 12298
rect 8006 12252 8074 12298
rect 8120 12252 8188 12298
rect 8234 12252 8302 12298
rect 8348 12252 8416 12298
rect 8462 12252 8530 12298
rect 8576 12252 8644 12298
rect 8690 12252 8758 12298
rect 8804 12252 8872 12298
rect 8918 12252 8986 12298
rect 9032 12252 9100 12298
rect 9146 12252 9214 12298
rect 9260 12252 9328 12298
rect 9374 12252 9442 12298
rect 9488 12252 9556 12298
rect 9602 12252 9670 12298
rect 9716 12252 9784 12298
rect 9830 12252 9898 12298
rect 9944 12252 10012 12298
rect 10058 12252 10126 12298
rect 10172 12252 10240 12298
rect 10286 12252 10394 12298
rect 10440 12252 10508 12298
rect 10554 12252 10565 12298
rect 43 12184 10565 12252
rect 43 12138 54 12184
rect 100 12138 168 12184
rect 214 12138 322 12184
rect 368 12138 436 12184
rect 482 12138 550 12184
rect 596 12138 664 12184
rect 710 12138 778 12184
rect 824 12138 892 12184
rect 938 12138 1006 12184
rect 1052 12138 1120 12184
rect 1166 12138 1234 12184
rect 1280 12138 1348 12184
rect 1394 12138 1462 12184
rect 1508 12138 1576 12184
rect 1622 12138 1690 12184
rect 1736 12138 1804 12184
rect 1850 12138 1918 12184
rect 1964 12138 2032 12184
rect 2078 12138 2146 12184
rect 2192 12138 2260 12184
rect 2306 12138 2374 12184
rect 2420 12138 2488 12184
rect 2534 12138 2602 12184
rect 2648 12138 2716 12184
rect 2762 12138 2830 12184
rect 2876 12138 2944 12184
rect 2990 12138 3058 12184
rect 3104 12138 3172 12184
rect 3218 12138 3286 12184
rect 3332 12138 3400 12184
rect 3446 12138 3514 12184
rect 3560 12138 3628 12184
rect 3674 12138 3742 12184
rect 3788 12138 3856 12184
rect 3902 12138 3970 12184
rect 4016 12138 4084 12184
rect 4130 12138 4198 12184
rect 4244 12138 4312 12184
rect 4358 12138 4426 12184
rect 4472 12138 4540 12184
rect 4586 12138 4654 12184
rect 4700 12138 4768 12184
rect 4814 12138 4882 12184
rect 4928 12138 4996 12184
rect 5042 12138 5110 12184
rect 5156 12138 5224 12184
rect 5270 12138 5338 12184
rect 5384 12138 5452 12184
rect 5498 12138 5566 12184
rect 5612 12138 5680 12184
rect 5726 12138 5794 12184
rect 5840 12138 5908 12184
rect 5954 12138 6022 12184
rect 6068 12138 6136 12184
rect 6182 12138 6250 12184
rect 6296 12138 6364 12184
rect 6410 12138 6478 12184
rect 6524 12138 6592 12184
rect 6638 12138 6706 12184
rect 6752 12138 6820 12184
rect 6866 12138 6934 12184
rect 6980 12138 7048 12184
rect 7094 12138 7162 12184
rect 7208 12138 7276 12184
rect 7322 12138 7390 12184
rect 7436 12138 7504 12184
rect 7550 12138 7618 12184
rect 7664 12138 7732 12184
rect 7778 12138 7846 12184
rect 7892 12138 7960 12184
rect 8006 12138 8074 12184
rect 8120 12138 8188 12184
rect 8234 12138 8302 12184
rect 8348 12138 8416 12184
rect 8462 12138 8530 12184
rect 8576 12138 8644 12184
rect 8690 12138 8758 12184
rect 8804 12138 8872 12184
rect 8918 12138 8986 12184
rect 9032 12138 9100 12184
rect 9146 12138 9214 12184
rect 9260 12138 9328 12184
rect 9374 12138 9442 12184
rect 9488 12138 9556 12184
rect 9602 12138 9670 12184
rect 9716 12138 9784 12184
rect 9830 12138 9898 12184
rect 9944 12138 10012 12184
rect 10058 12138 10126 12184
rect 10172 12138 10240 12184
rect 10286 12138 10394 12184
rect 10440 12138 10508 12184
rect 10554 12138 10565 12184
rect 43 12126 10565 12138
rect 43 12070 225 12126
rect 43 12024 54 12070
rect 100 12024 168 12070
rect 214 12024 225 12070
rect 43 11633 225 12024
rect 10383 12070 10565 12126
rect 10383 12024 10394 12070
rect 10440 12024 10508 12070
rect 10554 12024 10565 12070
rect 10383 11956 10565 12024
rect 10383 11910 10394 11956
rect 10440 11910 10508 11956
rect 10554 11910 10565 11956
rect 689 11723 9913 11855
rect 689 11712 2605 11723
rect 689 11666 700 11712
rect 2594 11666 2605 11712
rect 689 11655 2605 11666
rect 3125 11712 5041 11723
rect 3125 11666 3136 11712
rect 5030 11666 5041 11712
rect 3125 11655 5041 11666
rect 5561 11712 7477 11723
rect 5561 11666 5572 11712
rect 7466 11666 7477 11712
rect 5561 11655 7477 11666
rect 7997 11712 9913 11723
rect 7997 11666 8008 11712
rect 9902 11666 9913 11712
rect 7997 11655 9913 11666
rect 10383 11842 10565 11910
rect 10383 11796 10394 11842
rect 10440 11796 10508 11842
rect 10554 11796 10565 11842
rect 10383 11728 10565 11796
rect 10383 11682 10394 11728
rect 10440 11682 10508 11728
rect 10554 11682 10565 11728
rect 43 11596 629 11633
rect 43 11500 572 11596
rect 43 11454 54 11500
rect 100 11454 168 11500
rect 214 11454 572 11500
rect 43 11386 572 11454
rect 43 11340 54 11386
rect 100 11340 168 11386
rect 214 11340 572 11386
rect 43 11272 572 11340
rect 43 11226 54 11272
rect 100 11226 168 11272
rect 214 11226 572 11272
rect 43 11158 572 11226
rect 43 11112 54 11158
rect 100 11112 168 11158
rect 214 11112 572 11158
rect 43 11044 572 11112
rect 43 10998 54 11044
rect 100 10998 168 11044
rect 214 10998 572 11044
rect 43 10930 572 10998
rect 43 10884 54 10930
rect 100 10884 168 10930
rect 214 10884 572 10930
rect 43 10816 572 10884
rect 43 10770 54 10816
rect 100 10770 168 10816
rect 214 10770 572 10816
rect 43 10702 572 10770
rect 43 10656 54 10702
rect 100 10656 168 10702
rect 214 10656 572 10702
rect 43 10588 572 10656
rect 43 10542 54 10588
rect 100 10542 168 10588
rect 214 10542 572 10588
rect 43 10474 572 10542
rect 43 10428 54 10474
rect 100 10428 168 10474
rect 214 10428 572 10474
rect 43 10360 572 10428
rect 43 10314 54 10360
rect 100 10314 168 10360
rect 214 10314 572 10360
rect 43 10246 572 10314
rect 43 10200 54 10246
rect 100 10200 168 10246
rect 214 10200 572 10246
rect 43 10132 572 10200
rect 43 10086 54 10132
rect 100 10086 168 10132
rect 214 10086 572 10132
rect 43 10018 572 10086
rect 43 9972 54 10018
rect 100 9972 168 10018
rect 214 9972 572 10018
rect 43 9904 572 9972
rect 43 9858 54 9904
rect 100 9858 168 9904
rect 214 9858 572 9904
rect 43 9790 572 9858
rect 43 9744 54 9790
rect 100 9744 168 9790
rect 214 9744 572 9790
rect 43 9676 572 9744
rect 43 9630 54 9676
rect 100 9630 168 9676
rect 214 9630 572 9676
rect 43 9562 572 9630
rect 43 9516 54 9562
rect 100 9516 168 9562
rect 214 9516 572 9562
rect 43 9448 572 9516
rect 43 9402 54 9448
rect 100 9402 168 9448
rect 214 9402 572 9448
rect 43 9334 572 9402
rect 43 9288 54 9334
rect 100 9288 168 9334
rect 214 9288 572 9334
rect 43 9220 572 9288
rect 43 9174 54 9220
rect 100 9174 168 9220
rect 214 9174 572 9220
rect 43 9106 572 9174
rect 43 9060 54 9106
rect 100 9060 168 9106
rect 214 9060 572 9106
rect 43 8992 572 9060
rect 43 8946 54 8992
rect 100 8946 168 8992
rect 214 8946 572 8992
rect 43 8878 572 8946
rect 43 8832 54 8878
rect 100 8832 168 8878
rect 214 8832 572 8878
rect 43 8764 572 8832
rect 43 8718 54 8764
rect 100 8718 168 8764
rect 214 8718 572 8764
rect 43 8650 572 8718
rect 43 8604 54 8650
rect 100 8604 168 8650
rect 214 8604 572 8650
rect 43 8536 572 8604
rect 43 8490 54 8536
rect 100 8490 168 8536
rect 214 8490 572 8536
rect 43 8422 572 8490
rect 43 8376 54 8422
rect 100 8376 168 8422
rect 214 8376 572 8422
rect 43 8308 572 8376
rect 43 8262 54 8308
rect 100 8262 168 8308
rect 214 8262 572 8308
rect 43 8194 572 8262
rect 43 8148 54 8194
rect 100 8148 168 8194
rect 214 8148 572 8194
rect 43 8080 572 8148
rect 43 8034 54 8080
rect 100 8034 168 8080
rect 214 8034 572 8080
rect 43 7966 572 8034
rect 43 7920 54 7966
rect 100 7920 168 7966
rect 214 7920 572 7966
rect 43 7852 572 7920
rect 43 7806 54 7852
rect 100 7806 168 7852
rect 214 7806 572 7852
rect 43 7738 572 7806
rect 43 7692 54 7738
rect 100 7692 168 7738
rect 214 7692 572 7738
rect 43 7624 572 7692
rect 43 7578 54 7624
rect 100 7578 168 7624
rect 214 7578 572 7624
rect 43 7510 572 7578
rect 43 7464 54 7510
rect 100 7464 168 7510
rect 214 7464 572 7510
rect 43 7396 572 7464
rect 43 7350 54 7396
rect 100 7350 168 7396
rect 214 7350 572 7396
rect 43 7282 572 7350
rect 43 7236 54 7282
rect 100 7236 168 7282
rect 214 7236 572 7282
rect 43 7168 572 7236
rect 43 7122 54 7168
rect 100 7122 168 7168
rect 214 7122 572 7168
rect 43 7054 572 7122
rect 43 7008 54 7054
rect 100 7008 168 7054
rect 214 7008 572 7054
rect 43 6940 572 7008
rect 43 6894 54 6940
rect 100 6894 168 6940
rect 214 6894 572 6940
rect 43 6826 572 6894
rect 43 6780 54 6826
rect 100 6780 168 6826
rect 214 6780 572 6826
rect 43 6712 572 6780
rect 43 6666 54 6712
rect 100 6666 168 6712
rect 214 6670 572 6712
rect 618 6670 629 11596
rect 214 6666 629 6670
rect 43 6598 629 6666
rect 1147 6611 2147 11655
rect 2665 11596 3065 11633
rect 2665 6670 2676 11596
rect 2722 6670 3008 11596
rect 3054 6670 3065 11596
rect 43 6552 54 6598
rect 100 6552 168 6598
rect 214 6552 629 6598
rect 43 6484 629 6552
rect 689 6600 2605 6611
rect 689 6554 700 6600
rect 2594 6554 2605 6600
rect 689 6543 2605 6554
rect 43 6438 54 6484
rect 100 6438 168 6484
rect 214 6483 629 6484
rect 2665 6483 3065 6670
rect 3583 6611 4583 11655
rect 5101 11596 5501 11633
rect 5101 6670 5112 11596
rect 5158 6670 5444 11596
rect 5490 6670 5501 11596
rect 3125 6600 5041 6611
rect 3125 6554 3136 6600
rect 5030 6554 5041 6600
rect 3125 6543 5041 6554
rect 5101 6483 5501 6670
rect 6019 6611 7019 11655
rect 7537 11596 7937 11633
rect 7537 6670 7548 11596
rect 7594 6670 7880 11596
rect 7926 6670 7937 11596
rect 5561 6600 7477 6611
rect 5561 6554 5572 6600
rect 7466 6554 7477 6600
rect 5561 6543 7477 6554
rect 7537 6483 7937 6670
rect 8455 6611 9455 11655
rect 10383 11633 10565 11682
rect 9973 11614 10565 11633
rect 9973 11596 10394 11614
rect 9973 6670 9984 11596
rect 10030 11568 10394 11596
rect 10440 11568 10508 11614
rect 10554 11568 10565 11614
rect 10030 11500 10565 11568
rect 10030 11454 10394 11500
rect 10440 11454 10508 11500
rect 10554 11454 10565 11500
rect 10030 11386 10565 11454
rect 10030 11340 10394 11386
rect 10440 11340 10508 11386
rect 10554 11340 10565 11386
rect 10030 11272 10565 11340
rect 10030 11226 10394 11272
rect 10440 11226 10508 11272
rect 10554 11226 10565 11272
rect 10030 11158 10565 11226
rect 10030 11112 10394 11158
rect 10440 11112 10508 11158
rect 10554 11112 10565 11158
rect 10030 11044 10565 11112
rect 10030 10998 10394 11044
rect 10440 10998 10508 11044
rect 10554 10998 10565 11044
rect 10030 10930 10565 10998
rect 10030 10884 10394 10930
rect 10440 10884 10508 10930
rect 10554 10884 10565 10930
rect 10030 10816 10565 10884
rect 10030 10770 10394 10816
rect 10440 10770 10508 10816
rect 10554 10770 10565 10816
rect 10030 10702 10565 10770
rect 10030 10656 10394 10702
rect 10440 10656 10508 10702
rect 10554 10656 10565 10702
rect 10030 10588 10565 10656
rect 10030 10542 10394 10588
rect 10440 10542 10508 10588
rect 10554 10542 10565 10588
rect 10030 10474 10565 10542
rect 10030 10428 10394 10474
rect 10440 10428 10508 10474
rect 10554 10428 10565 10474
rect 10030 10360 10565 10428
rect 10030 10314 10394 10360
rect 10440 10314 10508 10360
rect 10554 10314 10565 10360
rect 10030 10246 10565 10314
rect 10030 10200 10394 10246
rect 10440 10200 10508 10246
rect 10554 10200 10565 10246
rect 10030 10132 10565 10200
rect 10030 10086 10394 10132
rect 10440 10086 10508 10132
rect 10554 10086 10565 10132
rect 10030 10018 10565 10086
rect 10030 9972 10394 10018
rect 10440 9972 10508 10018
rect 10554 9972 10565 10018
rect 10030 9904 10565 9972
rect 10030 9858 10394 9904
rect 10440 9858 10508 9904
rect 10554 9858 10565 9904
rect 10030 9790 10565 9858
rect 10030 9744 10394 9790
rect 10440 9744 10508 9790
rect 10554 9744 10565 9790
rect 10030 9676 10565 9744
rect 10030 9630 10394 9676
rect 10440 9630 10508 9676
rect 10554 9630 10565 9676
rect 10030 9562 10565 9630
rect 10030 9516 10394 9562
rect 10440 9516 10508 9562
rect 10554 9516 10565 9562
rect 10030 9448 10565 9516
rect 10030 9402 10394 9448
rect 10440 9402 10508 9448
rect 10554 9402 10565 9448
rect 10030 9334 10565 9402
rect 10030 9288 10394 9334
rect 10440 9288 10508 9334
rect 10554 9288 10565 9334
rect 10030 9220 10565 9288
rect 10030 9174 10394 9220
rect 10440 9174 10508 9220
rect 10554 9174 10565 9220
rect 10030 9106 10565 9174
rect 10030 9060 10394 9106
rect 10440 9060 10508 9106
rect 10554 9060 10565 9106
rect 10030 8992 10565 9060
rect 10030 8946 10394 8992
rect 10440 8946 10508 8992
rect 10554 8946 10565 8992
rect 10030 8878 10565 8946
rect 10030 8832 10394 8878
rect 10440 8832 10508 8878
rect 10554 8832 10565 8878
rect 10030 8764 10565 8832
rect 10030 8718 10394 8764
rect 10440 8718 10508 8764
rect 10554 8718 10565 8764
rect 10030 8650 10565 8718
rect 10030 8604 10394 8650
rect 10440 8604 10508 8650
rect 10554 8604 10565 8650
rect 10030 8536 10565 8604
rect 10030 8490 10394 8536
rect 10440 8490 10508 8536
rect 10554 8490 10565 8536
rect 10030 8422 10565 8490
rect 10030 8376 10394 8422
rect 10440 8376 10508 8422
rect 10554 8376 10565 8422
rect 10030 8308 10565 8376
rect 10030 8262 10394 8308
rect 10440 8262 10508 8308
rect 10554 8262 10565 8308
rect 10030 8194 10565 8262
rect 10030 8148 10394 8194
rect 10440 8148 10508 8194
rect 10554 8148 10565 8194
rect 10030 8080 10565 8148
rect 10030 8034 10394 8080
rect 10440 8034 10508 8080
rect 10554 8034 10565 8080
rect 10030 7966 10565 8034
rect 10030 7920 10394 7966
rect 10440 7920 10508 7966
rect 10554 7920 10565 7966
rect 10030 7852 10565 7920
rect 10030 7806 10394 7852
rect 10440 7806 10508 7852
rect 10554 7806 10565 7852
rect 10030 7738 10565 7806
rect 10030 7692 10394 7738
rect 10440 7692 10508 7738
rect 10554 7692 10565 7738
rect 10030 7624 10565 7692
rect 10030 7578 10394 7624
rect 10440 7578 10508 7624
rect 10554 7578 10565 7624
rect 10030 7510 10565 7578
rect 10030 7464 10394 7510
rect 10440 7464 10508 7510
rect 10554 7464 10565 7510
rect 10030 7396 10565 7464
rect 10030 7350 10394 7396
rect 10440 7350 10508 7396
rect 10554 7350 10565 7396
rect 10030 7282 10565 7350
rect 10030 7236 10394 7282
rect 10440 7236 10508 7282
rect 10554 7236 10565 7282
rect 10030 7168 10565 7236
rect 10030 7122 10394 7168
rect 10440 7122 10508 7168
rect 10554 7122 10565 7168
rect 10030 7054 10565 7122
rect 10030 7008 10394 7054
rect 10440 7008 10508 7054
rect 10554 7008 10565 7054
rect 10030 6940 10565 7008
rect 10030 6894 10394 6940
rect 10440 6894 10508 6940
rect 10554 6894 10565 6940
rect 10030 6826 10565 6894
rect 10030 6780 10394 6826
rect 10440 6780 10508 6826
rect 10554 6780 10565 6826
rect 10030 6712 10565 6780
rect 10030 6670 10394 6712
rect 9973 6666 10394 6670
rect 10440 6666 10508 6712
rect 10554 6666 10565 6712
rect 7997 6600 9913 6611
rect 7997 6554 8008 6600
rect 9902 6554 9913 6600
rect 7997 6543 9913 6554
rect 9973 6598 10565 6666
rect 9973 6552 10394 6598
rect 10440 6552 10508 6598
rect 10554 6552 10565 6598
rect 9973 6484 10565 6552
rect 9973 6483 10394 6484
rect 214 6438 10394 6483
rect 10440 6438 10508 6484
rect 10554 6438 10565 6484
rect 43 6370 10565 6438
rect 43 6324 54 6370
rect 100 6324 168 6370
rect 214 6324 10394 6370
rect 10440 6324 10508 6370
rect 10554 6324 10565 6370
rect 43 6256 10565 6324
rect 43 6210 10394 6256
rect 10440 6210 10508 6256
rect 10554 6210 10565 6256
rect 43 6207 10565 6210
rect 43 6161 322 6207
rect 368 6161 436 6207
rect 482 6161 550 6207
rect 596 6161 664 6207
rect 710 6161 778 6207
rect 824 6161 892 6207
rect 938 6161 1006 6207
rect 1052 6161 1120 6207
rect 1166 6161 1234 6207
rect 1280 6161 1348 6207
rect 1394 6161 1462 6207
rect 1508 6161 1576 6207
rect 1622 6161 1690 6207
rect 1736 6161 1804 6207
rect 1850 6161 1918 6207
rect 1964 6161 2032 6207
rect 2078 6161 2146 6207
rect 2192 6161 2260 6207
rect 2306 6161 2374 6207
rect 2420 6161 2488 6207
rect 2534 6161 2602 6207
rect 2648 6161 2716 6207
rect 2762 6161 2830 6207
rect 2876 6161 2944 6207
rect 2990 6161 3058 6207
rect 3104 6161 3172 6207
rect 3218 6161 3286 6207
rect 3332 6161 3400 6207
rect 3446 6161 3514 6207
rect 3560 6161 3628 6207
rect 3674 6161 3742 6207
rect 3788 6161 3856 6207
rect 3902 6161 3970 6207
rect 4016 6161 4084 6207
rect 4130 6161 4198 6207
rect 4244 6161 4312 6207
rect 4358 6161 4426 6207
rect 4472 6161 4540 6207
rect 4586 6161 4654 6207
rect 4700 6161 4768 6207
rect 4814 6161 4882 6207
rect 4928 6161 4996 6207
rect 5042 6161 5110 6207
rect 5156 6161 5224 6207
rect 5270 6161 5338 6207
rect 5384 6161 5452 6207
rect 5498 6161 5566 6207
rect 5612 6161 5680 6207
rect 5726 6161 5794 6207
rect 5840 6161 5908 6207
rect 5954 6161 6022 6207
rect 6068 6161 6136 6207
rect 6182 6161 6250 6207
rect 6296 6161 6364 6207
rect 6410 6161 6478 6207
rect 6524 6161 6592 6207
rect 6638 6161 6706 6207
rect 6752 6161 6820 6207
rect 6866 6161 6934 6207
rect 6980 6161 7048 6207
rect 7094 6161 7162 6207
rect 7208 6161 7276 6207
rect 7322 6161 7390 6207
rect 7436 6161 7504 6207
rect 7550 6161 7618 6207
rect 7664 6161 7732 6207
rect 7778 6161 7846 6207
rect 7892 6161 7960 6207
rect 8006 6161 8074 6207
rect 8120 6161 8188 6207
rect 8234 6161 8302 6207
rect 8348 6161 8416 6207
rect 8462 6161 8530 6207
rect 8576 6161 8644 6207
rect 8690 6161 8758 6207
rect 8804 6161 8872 6207
rect 8918 6161 8986 6207
rect 9032 6161 9100 6207
rect 9146 6161 9214 6207
rect 9260 6161 9328 6207
rect 9374 6161 9442 6207
rect 9488 6161 9556 6207
rect 9602 6161 9670 6207
rect 9716 6161 9784 6207
rect 9830 6161 9898 6207
rect 9944 6161 10012 6207
rect 10058 6161 10126 6207
rect 10172 6161 10240 6207
rect 10286 6161 10565 6207
rect 43 6142 10565 6161
rect 43 6096 10394 6142
rect 10440 6096 10508 6142
rect 10554 6096 10565 6142
rect 43 6093 10565 6096
rect 43 6047 322 6093
rect 368 6047 436 6093
rect 482 6047 550 6093
rect 596 6047 664 6093
rect 710 6047 778 6093
rect 824 6047 892 6093
rect 938 6047 1006 6093
rect 1052 6047 1120 6093
rect 1166 6047 1234 6093
rect 1280 6047 1348 6093
rect 1394 6047 1462 6093
rect 1508 6047 1576 6093
rect 1622 6047 1690 6093
rect 1736 6047 1804 6093
rect 1850 6047 1918 6093
rect 1964 6047 2032 6093
rect 2078 6047 2146 6093
rect 2192 6047 2260 6093
rect 2306 6047 2374 6093
rect 2420 6047 2488 6093
rect 2534 6047 2602 6093
rect 2648 6047 2716 6093
rect 2762 6047 2830 6093
rect 2876 6047 2944 6093
rect 2990 6047 3058 6093
rect 3104 6047 3172 6093
rect 3218 6047 3286 6093
rect 3332 6047 3400 6093
rect 3446 6047 3514 6093
rect 3560 6047 3628 6093
rect 3674 6047 3742 6093
rect 3788 6047 3856 6093
rect 3902 6047 3970 6093
rect 4016 6047 4084 6093
rect 4130 6047 4198 6093
rect 4244 6047 4312 6093
rect 4358 6047 4426 6093
rect 4472 6047 4540 6093
rect 4586 6047 4654 6093
rect 4700 6047 4768 6093
rect 4814 6047 4882 6093
rect 4928 6047 4996 6093
rect 5042 6047 5110 6093
rect 5156 6047 5224 6093
rect 5270 6047 5338 6093
rect 5384 6047 5452 6093
rect 5498 6047 5566 6093
rect 5612 6047 5680 6093
rect 5726 6047 5794 6093
rect 5840 6047 5908 6093
rect 5954 6047 6022 6093
rect 6068 6047 6136 6093
rect 6182 6047 6250 6093
rect 6296 6047 6364 6093
rect 6410 6047 6478 6093
rect 6524 6047 6592 6093
rect 6638 6047 6706 6093
rect 6752 6047 6820 6093
rect 6866 6047 6934 6093
rect 6980 6047 7048 6093
rect 7094 6047 7162 6093
rect 7208 6047 7276 6093
rect 7322 6047 7390 6093
rect 7436 6047 7504 6093
rect 7550 6047 7618 6093
rect 7664 6047 7732 6093
rect 7778 6047 7846 6093
rect 7892 6047 7960 6093
rect 8006 6047 8074 6093
rect 8120 6047 8188 6093
rect 8234 6047 8302 6093
rect 8348 6047 8416 6093
rect 8462 6047 8530 6093
rect 8576 6047 8644 6093
rect 8690 6047 8758 6093
rect 8804 6047 8872 6093
rect 8918 6047 8986 6093
rect 9032 6047 9100 6093
rect 9146 6047 9214 6093
rect 9260 6047 9328 6093
rect 9374 6047 9442 6093
rect 9488 6047 9556 6093
rect 9602 6047 9670 6093
rect 9716 6047 9784 6093
rect 9830 6047 9898 6093
rect 9944 6047 10012 6093
rect 10058 6047 10126 6093
rect 10172 6047 10240 6093
rect 10286 6047 10565 6093
rect 43 6028 10565 6047
rect 43 5982 10394 6028
rect 10440 5982 10508 6028
rect 10554 5982 10565 6028
rect 43 5951 10565 5982
rect 43 5905 5020 5951
rect 5066 5914 10565 5951
rect 5066 5905 10394 5914
rect 43 5868 10394 5905
rect 10440 5868 10508 5914
rect 10554 5868 10565 5914
rect 43 5827 10565 5868
rect 43 5781 5020 5827
rect 5066 5800 10565 5827
rect 5066 5781 10394 5800
rect 43 5771 10394 5781
rect 5009 5703 5501 5771
rect 5009 5657 5020 5703
rect 5066 5657 5501 5703
rect 5009 5584 5501 5657
rect 5561 5700 7477 5711
rect 5561 5654 5572 5700
rect 7466 5654 7477 5700
rect 5561 5643 7477 5654
rect 5009 5579 5444 5584
rect 5009 5533 5020 5579
rect 5066 5533 5444 5579
rect 5009 5455 5444 5533
rect 5009 5409 5020 5455
rect 5066 5409 5444 5455
rect 5009 5331 5444 5409
rect 5009 5285 5020 5331
rect 5066 5285 5444 5331
rect 5009 5207 5444 5285
rect 5009 5161 5020 5207
rect 5066 5161 5444 5207
rect 5009 5083 5444 5161
rect 5009 5037 5020 5083
rect 5066 5037 5444 5083
rect 5009 4959 5444 5037
rect 5009 4913 5020 4959
rect 5066 4913 5444 4959
rect 5009 4835 5444 4913
rect 5009 4789 5020 4835
rect 5066 4789 5444 4835
rect 5009 4711 5444 4789
rect 5009 4665 5020 4711
rect 5066 4665 5444 4711
rect 5009 4587 5444 4665
rect 5009 4541 5020 4587
rect 5066 4541 5444 4587
rect 5009 4463 5444 4541
rect 5009 4417 5020 4463
rect 5066 4417 5444 4463
rect 5009 4339 5444 4417
rect 5009 4293 5020 4339
rect 5066 4293 5444 4339
rect 5009 4215 5444 4293
rect 5009 4169 5020 4215
rect 5066 4169 5444 4215
rect 5009 4091 5444 4169
rect 5009 4045 5020 4091
rect 5066 4045 5444 4091
rect 5009 3967 5444 4045
rect 5009 3921 5020 3967
rect 5066 3921 5444 3967
rect 5009 3843 5444 3921
rect 5009 3797 5020 3843
rect 5066 3797 5444 3843
rect 5009 3719 5444 3797
rect 5009 3673 5020 3719
rect 5066 3673 5444 3719
rect 5009 3595 5444 3673
rect 5009 3549 5020 3595
rect 5066 3549 5444 3595
rect 5009 3471 5444 3549
rect 5009 3425 5020 3471
rect 5066 3425 5444 3471
rect 5009 3347 5444 3425
rect 5009 3301 5020 3347
rect 5066 3301 5444 3347
rect 5009 3223 5444 3301
rect 5009 3177 5020 3223
rect 5066 3177 5444 3223
rect 5009 3099 5444 3177
rect 5009 3053 5020 3099
rect 5066 3053 5444 3099
rect 5009 2975 5444 3053
rect 5009 2929 5020 2975
rect 5066 2929 5444 2975
rect 5009 2851 5444 2929
rect 5009 2805 5020 2851
rect 5066 2805 5444 2851
rect 5009 2727 5444 2805
rect 5009 2681 5020 2727
rect 5066 2681 5444 2727
rect 5009 2603 5444 2681
rect 5009 2557 5020 2603
rect 5066 2557 5444 2603
rect 5009 2479 5444 2557
rect 5009 2433 5020 2479
rect 5066 2433 5444 2479
rect 5009 2355 5444 2433
rect 5009 2309 5020 2355
rect 5066 2309 5444 2355
rect 5009 2231 5444 2309
rect 5009 2185 5020 2231
rect 5066 2185 5444 2231
rect 5009 2107 5444 2185
rect 5009 2061 5020 2107
rect 5066 2061 5444 2107
rect 5009 1983 5444 2061
rect 5009 1937 5020 1983
rect 5066 1937 5444 1983
rect 5009 1859 5444 1937
rect 5009 1813 5020 1859
rect 5066 1813 5444 1859
rect 5009 1735 5444 1813
rect 5009 1689 5020 1735
rect 5066 1689 5444 1735
rect 5009 1611 5444 1689
rect 5009 1565 5020 1611
rect 5066 1565 5444 1611
rect 5009 1487 5444 1565
rect 5009 1441 5020 1487
rect 5066 1441 5444 1487
rect 5009 1363 5444 1441
rect 5009 1317 5020 1363
rect 5066 1317 5444 1363
rect 5009 1239 5444 1317
rect 5009 1193 5020 1239
rect 5066 1193 5444 1239
rect 5009 1115 5444 1193
rect 5009 1069 5020 1115
rect 5066 1069 5444 1115
rect 5009 991 5444 1069
rect 5009 945 5020 991
rect 5066 945 5444 991
rect 5009 867 5444 945
rect 5009 821 5020 867
rect 5066 821 5444 867
rect 5009 743 5444 821
rect 5009 697 5020 743
rect 5066 697 5444 743
rect 5009 658 5444 697
rect 5490 658 5501 5584
rect 5009 621 5501 658
rect 5009 619 5301 621
rect 5009 573 5020 619
rect 5066 573 5301 619
rect 6019 599 7019 5643
rect 7537 5584 7937 5771
rect 9973 5754 10394 5771
rect 10440 5754 10508 5800
rect 10554 5754 10565 5800
rect 7997 5700 9913 5711
rect 7997 5654 8008 5700
rect 9902 5654 9913 5700
rect 7997 5643 9913 5654
rect 9973 5686 10565 5754
rect 7537 658 7548 5584
rect 7594 658 7880 5584
rect 7926 658 7937 5584
rect 7537 621 7937 658
rect 8455 599 9455 5643
rect 9973 5640 10394 5686
rect 10440 5640 10508 5686
rect 10554 5640 10565 5686
rect 9973 5584 10565 5640
rect 9973 658 9984 5584
rect 10030 5572 10565 5584
rect 10030 5526 10394 5572
rect 10440 5526 10508 5572
rect 10554 5526 10565 5572
rect 10030 5458 10565 5526
rect 10030 5412 10394 5458
rect 10440 5412 10508 5458
rect 10554 5412 10565 5458
rect 10030 5344 10565 5412
rect 10030 5298 10394 5344
rect 10440 5298 10508 5344
rect 10554 5298 10565 5344
rect 10030 5230 10565 5298
rect 10030 5184 10394 5230
rect 10440 5184 10508 5230
rect 10554 5184 10565 5230
rect 10030 5116 10565 5184
rect 10030 5070 10394 5116
rect 10440 5070 10508 5116
rect 10554 5070 10565 5116
rect 10030 5002 10565 5070
rect 10030 4956 10394 5002
rect 10440 4956 10508 5002
rect 10554 4956 10565 5002
rect 10030 4888 10565 4956
rect 10030 4842 10394 4888
rect 10440 4842 10508 4888
rect 10554 4842 10565 4888
rect 10030 4774 10565 4842
rect 10030 4728 10394 4774
rect 10440 4728 10508 4774
rect 10554 4728 10565 4774
rect 10030 4660 10565 4728
rect 10030 4614 10394 4660
rect 10440 4614 10508 4660
rect 10554 4614 10565 4660
rect 10030 4546 10565 4614
rect 10030 4500 10394 4546
rect 10440 4500 10508 4546
rect 10554 4500 10565 4546
rect 10030 4432 10565 4500
rect 10030 4386 10394 4432
rect 10440 4386 10508 4432
rect 10554 4386 10565 4432
rect 10030 4318 10565 4386
rect 10030 4272 10394 4318
rect 10440 4272 10508 4318
rect 10554 4272 10565 4318
rect 10030 4204 10565 4272
rect 10030 4158 10394 4204
rect 10440 4158 10508 4204
rect 10554 4158 10565 4204
rect 10030 4090 10565 4158
rect 10030 4044 10394 4090
rect 10440 4044 10508 4090
rect 10554 4044 10565 4090
rect 10030 3976 10565 4044
rect 10030 3930 10394 3976
rect 10440 3930 10508 3976
rect 10554 3930 10565 3976
rect 10030 3862 10565 3930
rect 10030 3816 10394 3862
rect 10440 3816 10508 3862
rect 10554 3816 10565 3862
rect 10030 3748 10565 3816
rect 10030 3702 10394 3748
rect 10440 3702 10508 3748
rect 10554 3702 10565 3748
rect 10030 3634 10565 3702
rect 10030 3588 10394 3634
rect 10440 3588 10508 3634
rect 10554 3588 10565 3634
rect 10030 3520 10565 3588
rect 10030 3474 10394 3520
rect 10440 3474 10508 3520
rect 10554 3474 10565 3520
rect 10030 3406 10565 3474
rect 10030 3360 10394 3406
rect 10440 3360 10508 3406
rect 10554 3360 10565 3406
rect 10030 3292 10565 3360
rect 10030 3246 10394 3292
rect 10440 3246 10508 3292
rect 10554 3246 10565 3292
rect 10030 3178 10565 3246
rect 10030 3132 10394 3178
rect 10440 3132 10508 3178
rect 10554 3132 10565 3178
rect 10030 3064 10565 3132
rect 10030 3018 10394 3064
rect 10440 3018 10508 3064
rect 10554 3018 10565 3064
rect 10030 2950 10565 3018
rect 10030 2904 10394 2950
rect 10440 2904 10508 2950
rect 10554 2904 10565 2950
rect 10030 2836 10565 2904
rect 10030 2790 10394 2836
rect 10440 2790 10508 2836
rect 10554 2790 10565 2836
rect 10030 2722 10565 2790
rect 10030 2676 10394 2722
rect 10440 2676 10508 2722
rect 10554 2676 10565 2722
rect 10030 2608 10565 2676
rect 10030 2562 10394 2608
rect 10440 2562 10508 2608
rect 10554 2562 10565 2608
rect 10030 2494 10565 2562
rect 10030 2448 10394 2494
rect 10440 2448 10508 2494
rect 10554 2448 10565 2494
rect 10030 2380 10565 2448
rect 10030 2334 10394 2380
rect 10440 2334 10508 2380
rect 10554 2334 10565 2380
rect 10030 2266 10565 2334
rect 10030 2220 10394 2266
rect 10440 2220 10508 2266
rect 10554 2220 10565 2266
rect 10030 2152 10565 2220
rect 10030 2106 10394 2152
rect 10440 2106 10508 2152
rect 10554 2106 10565 2152
rect 10030 2038 10565 2106
rect 10030 1992 10394 2038
rect 10440 1992 10508 2038
rect 10554 1992 10565 2038
rect 10030 1924 10565 1992
rect 10030 1878 10394 1924
rect 10440 1878 10508 1924
rect 10554 1878 10565 1924
rect 10030 1810 10565 1878
rect 10030 1764 10394 1810
rect 10440 1764 10508 1810
rect 10554 1764 10565 1810
rect 10030 1696 10565 1764
rect 10030 1650 10394 1696
rect 10440 1650 10508 1696
rect 10554 1650 10565 1696
rect 10030 1582 10565 1650
rect 10030 1536 10394 1582
rect 10440 1536 10508 1582
rect 10554 1536 10565 1582
rect 10030 1468 10565 1536
rect 10030 1422 10394 1468
rect 10440 1422 10508 1468
rect 10554 1422 10565 1468
rect 10030 1354 10565 1422
rect 10030 1308 10394 1354
rect 10440 1308 10508 1354
rect 10554 1308 10565 1354
rect 10030 1240 10565 1308
rect 10030 1194 10394 1240
rect 10440 1194 10508 1240
rect 10554 1194 10565 1240
rect 10030 1126 10565 1194
rect 10030 1080 10394 1126
rect 10440 1080 10508 1126
rect 10554 1080 10565 1126
rect 10030 1012 10565 1080
rect 10030 966 10394 1012
rect 10440 966 10508 1012
rect 10554 966 10565 1012
rect 10030 898 10565 966
rect 10030 852 10394 898
rect 10440 852 10508 898
rect 10554 852 10565 898
rect 10030 784 10565 852
rect 10030 738 10394 784
rect 10440 738 10508 784
rect 10554 738 10565 784
rect 10030 670 10565 738
rect 10030 658 10394 670
rect 9973 624 10394 658
rect 10440 624 10508 670
rect 10554 624 10565 670
rect 9973 621 10565 624
rect 5009 495 5301 573
rect 5009 449 5020 495
rect 5066 449 5301 495
rect 5009 371 5301 449
rect 5561 588 7477 599
rect 5561 542 5572 588
rect 7466 542 7477 588
rect 5561 531 7477 542
rect 7997 588 9913 599
rect 7997 542 8008 588
rect 9902 542 9913 588
rect 7997 531 9913 542
rect 5561 399 9913 531
rect 10383 556 10565 621
rect 10383 510 10394 556
rect 10440 510 10508 556
rect 10554 510 10565 556
rect 10383 442 10565 510
rect 5009 325 5020 371
rect 5066 325 5301 371
rect 5009 247 5301 325
rect 5009 201 5020 247
rect 5066 226 5301 247
rect 10383 396 10394 442
rect 10440 396 10508 442
rect 10554 396 10565 442
rect 10383 328 10565 396
rect 10383 282 10394 328
rect 10440 282 10508 328
rect 10554 282 10565 328
rect 10383 226 10565 282
rect 5066 214 10565 226
rect 5066 201 5354 214
rect 5009 168 5354 201
rect 5400 168 5468 214
rect 5514 168 5582 214
rect 5628 168 5696 214
rect 5742 168 5810 214
rect 5856 168 5924 214
rect 5970 168 6038 214
rect 6084 168 6152 214
rect 6198 168 6266 214
rect 6312 168 6380 214
rect 6426 168 6494 214
rect 6540 168 6608 214
rect 6654 168 6722 214
rect 6768 168 6836 214
rect 6882 168 6950 214
rect 6996 168 7064 214
rect 7110 168 7178 214
rect 7224 168 7292 214
rect 7338 168 7406 214
rect 7452 168 7520 214
rect 7566 168 7634 214
rect 7680 168 7748 214
rect 7794 168 7862 214
rect 7908 168 7976 214
rect 8022 168 8090 214
rect 8136 168 8204 214
rect 8250 168 8318 214
rect 8364 168 8432 214
rect 8478 168 8546 214
rect 8592 168 8660 214
rect 8706 168 8774 214
rect 8820 168 8888 214
rect 8934 168 9002 214
rect 9048 168 9116 214
rect 9162 168 9230 214
rect 9276 168 9344 214
rect 9390 168 9458 214
rect 9504 168 9572 214
rect 9618 168 9686 214
rect 9732 168 9800 214
rect 9846 168 9914 214
rect 9960 168 10028 214
rect 10074 168 10142 214
rect 10188 168 10256 214
rect 10302 168 10394 214
rect 10440 168 10508 214
rect 10554 168 10565 214
rect 5009 123 10565 168
rect 5009 77 5020 123
rect 5066 100 10565 123
rect 5066 77 5354 100
rect 5009 54 5354 77
rect 5400 54 5468 100
rect 5514 54 5582 100
rect 5628 54 5696 100
rect 5742 54 5810 100
rect 5856 54 5924 100
rect 5970 54 6038 100
rect 6084 54 6152 100
rect 6198 54 6266 100
rect 6312 54 6380 100
rect 6426 54 6494 100
rect 6540 54 6608 100
rect 6654 54 6722 100
rect 6768 54 6836 100
rect 6882 54 6950 100
rect 6996 54 7064 100
rect 7110 54 7178 100
rect 7224 54 7292 100
rect 7338 54 7406 100
rect 7452 54 7520 100
rect 7566 54 7634 100
rect 7680 54 7748 100
rect 7794 54 7862 100
rect 7908 54 7976 100
rect 8022 54 8090 100
rect 8136 54 8204 100
rect 8250 54 8318 100
rect 8364 54 8432 100
rect 8478 54 8546 100
rect 8592 54 8660 100
rect 8706 54 8774 100
rect 8820 54 8888 100
rect 8934 54 9002 100
rect 9048 54 9116 100
rect 9162 54 9230 100
rect 9276 54 9344 100
rect 9390 54 9458 100
rect 9504 54 9572 100
rect 9618 54 9686 100
rect 9732 54 9800 100
rect 9846 54 9914 100
rect 9960 54 10028 100
rect 10074 54 10142 100
rect 10188 54 10256 100
rect 10302 54 10394 100
rect 10440 54 10508 100
rect 10554 54 10565 100
rect 5009 42 10565 54
use M1_PSUB_CDNS_40661953145126  M1_PSUB_CDNS_40661953145126_0
timestamp 1749760379
transform 1 0 10474 0 1 6176
box 0 0 1 1
use M1_PSUB_CDNS_40661953145129  M1_PSUB_CDNS_40661953145129_0
timestamp 1749760379
transform 0 -1 5304 1 0 12218
box 0 0 1 1
use M1_PSUB_CDNS_40661953145129  M1_PSUB_CDNS_40661953145129_1
timestamp 1749760379
transform 0 -1 5304 1 0 6127
box 0 0 1 1
use M1_PSUB_CDNS_40661953145679  M1_PSUB_CDNS_40661953145679_0
timestamp 1749760379
transform 0 -1 7828 1 0 134
box 0 0 1 1
use M1_PSUB_CDNS_40661953145680  M1_PSUB_CDNS_40661953145680_0
timestamp 1749760379
transform 1 0 5043 0 1 3014
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_0
timestamp 1749760379
transform 1 0 7955 0 -1 5621
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_1
timestamp 1749760379
transform 1 0 5519 0 -1 5621
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_2
timestamp 1749760379
transform 1 0 7955 0 1 6633
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_3
timestamp 1749760379
transform 1 0 5519 0 1 6633
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_4
timestamp 1749760379
transform 1 0 3083 0 1 6633
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_5
timestamp 1749760379
transform 1 0 647 0 1 6633
box 0 0 1 1
<< labels >>
rlabel metal1 s 5302 6126 5302 6126 4 VMINUS
port 1 nsew
<< properties >>
string GDS_END 5159068
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 5150820
<< end >>
