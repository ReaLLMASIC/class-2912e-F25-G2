magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 352 1878 870
<< pwell >>
rect -86 -86 1878 352
<< mvnmos >>
rect 179 68 299 140
rect 403 68 523 140
rect 571 68 691 140
rect 1027 68 1147 141
rect 1195 68 1315 141
rect 1525 68 1645 232
<< mvpmos >>
rect 179 644 279 716
rect 403 644 503 716
rect 571 644 671 716
rect 1027 622 1127 694
rect 1195 622 1295 694
rect 1525 472 1625 716
<< mvndiff >>
rect 47 180 119 193
rect 47 134 60 180
rect 106 140 119 180
rect 751 200 823 213
rect 751 154 764 200
rect 810 154 823 200
rect 751 140 823 154
rect 106 134 179 140
rect 47 68 179 134
rect 299 127 403 140
rect 299 81 328 127
rect 374 81 403 127
rect 299 68 403 81
rect 523 68 571 140
rect 691 68 823 140
rect 895 200 967 213
rect 895 154 908 200
rect 954 154 967 200
rect 895 141 967 154
rect 1445 141 1525 232
rect 895 68 1027 141
rect 1147 68 1195 141
rect 1315 127 1525 141
rect 1315 81 1344 127
rect 1390 81 1525 127
rect 1315 68 1525 81
rect 1645 192 1733 232
rect 1645 146 1674 192
rect 1720 146 1733 192
rect 1645 68 1733 146
<< mvpdiff >>
rect 47 644 179 716
rect 279 703 403 716
rect 279 657 308 703
rect 354 657 403 703
rect 279 644 403 657
rect 503 644 571 716
rect 671 644 803 716
rect 1445 694 1525 716
rect 47 621 119 644
rect 47 575 60 621
rect 106 575 119 621
rect 47 562 119 575
rect 731 621 803 644
rect 731 575 744 621
rect 790 575 803 621
rect 731 562 803 575
rect 895 622 1027 694
rect 1127 622 1195 694
rect 1295 681 1525 694
rect 1295 635 1324 681
rect 1370 635 1525 681
rect 1295 622 1525 635
rect 895 621 967 622
rect 895 575 908 621
rect 954 575 967 621
rect 895 562 967 575
rect 1445 472 1525 622
rect 1625 639 1713 716
rect 1625 593 1654 639
rect 1700 593 1713 639
rect 1625 531 1713 593
rect 1625 485 1654 531
rect 1700 485 1713 531
rect 1625 472 1713 485
<< mvndiffc >>
rect 60 134 106 180
rect 764 154 810 200
rect 328 81 374 127
rect 908 154 954 200
rect 1344 81 1390 127
rect 1674 146 1720 192
<< mvpdiffc >>
rect 308 657 354 703
rect 60 575 106 621
rect 744 575 790 621
rect 1324 635 1370 681
rect 908 575 954 621
rect 1654 593 1700 639
rect 1654 485 1700 531
<< polysilicon >>
rect 179 716 279 760
rect 403 716 503 760
rect 571 716 671 760
rect 1027 694 1127 738
rect 1195 694 1295 738
rect 1525 716 1625 760
rect 179 303 279 644
rect 179 257 192 303
rect 238 257 279 303
rect 179 184 279 257
rect 403 483 503 644
rect 571 483 671 644
rect 403 470 671 483
rect 403 424 416 470
rect 462 424 596 470
rect 642 424 671 470
rect 403 411 671 424
rect 403 184 503 411
rect 571 184 671 411
rect 1027 399 1127 622
rect 1195 399 1295 622
rect 1027 382 1295 399
rect 1027 336 1040 382
rect 1086 344 1295 382
rect 1086 336 1127 344
rect 1027 251 1127 336
rect 1195 251 1295 344
rect 1525 325 1625 472
rect 1525 279 1538 325
rect 1584 323 1625 325
rect 1584 279 1645 323
rect 179 140 299 184
rect 403 140 523 184
rect 571 140 691 184
rect 1027 141 1147 251
rect 1195 141 1315 251
rect 1525 232 1645 279
rect 179 24 299 68
rect 403 24 523 68
rect 571 24 691 68
rect 1027 24 1147 68
rect 1195 24 1315 68
rect 1525 24 1645 68
<< polycontact >>
rect 192 257 238 303
rect 416 424 462 470
rect 596 424 642 470
rect 1040 336 1086 382
rect 1538 279 1584 325
<< metal1 >>
rect 0 724 1792 844
rect 297 703 365 724
rect 297 657 308 703
rect 354 657 365 703
rect 1313 681 1381 724
rect 1313 635 1324 681
rect 1370 635 1381 681
rect 744 621 790 632
rect 49 575 60 621
rect 106 575 117 621
rect 49 481 117 575
rect 49 470 653 481
rect 49 424 416 470
rect 462 424 596 470
rect 642 424 653 470
rect 49 413 653 424
rect 49 180 95 413
rect 744 382 790 575
rect 908 621 954 632
rect 908 493 954 575
rect 1643 593 1654 639
rect 1700 593 1720 639
rect 1643 542 1720 593
rect 1362 531 1720 542
rect 908 447 1231 493
rect 1362 485 1654 531
rect 1700 485 1720 531
rect 1362 466 1720 485
rect 744 336 1040 382
rect 1086 336 1097 382
rect 186 303 671 320
rect 186 257 192 303
rect 238 257 671 303
rect 186 240 671 257
rect 744 200 821 336
rect 1167 325 1231 447
rect 1167 279 1538 325
rect 1584 279 1595 325
rect 1167 211 1231 279
rect 49 134 60 180
rect 106 134 117 180
rect 744 154 764 200
rect 810 154 821 200
rect 908 200 1231 211
rect 954 154 1231 200
rect 908 143 1231 154
rect 1674 192 1720 466
rect 1344 127 1390 138
rect 1674 135 1720 146
rect 317 81 328 127
rect 374 81 385 127
rect 317 60 385 81
rect 1344 60 1390 81
rect 0 -60 1792 60
<< labels >>
flabel metal1 s 0 724 1792 844 0 FreeSans 400 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 186 240 671 320 0 FreeSans 400 0 0 0 I
port 1 nsew default input
flabel metal1 s 1344 127 1390 138 0 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 1643 542 1720 639 0 FreeSans 400 0 0 0 Z
port 2 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 1362 466 1720 542 1 Z
port 2 nsew default output
rlabel metal1 s 1674 135 1720 466 1 Z
port 2 nsew default output
rlabel metal1 s 1313 657 1381 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 297 657 365 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1313 635 1381 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1344 60 1390 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 317 60 385 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1792 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1792 784
string GDS_END 1094044
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1090088
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
