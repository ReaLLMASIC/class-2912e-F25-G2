magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< metal1 >>
rect 28 945 972 957
rect 28 893 40 945
rect 92 893 164 945
rect 216 893 288 945
rect 340 893 412 945
rect 464 893 536 945
rect 588 893 660 945
rect 712 893 784 945
rect 836 893 908 945
rect 960 893 972 945
rect 28 821 972 893
rect 28 769 40 821
rect 92 769 164 821
rect 216 769 288 821
rect 340 769 412 821
rect 464 769 536 821
rect 588 769 660 821
rect 712 769 784 821
rect 836 769 908 821
rect 960 769 972 821
rect 28 697 972 769
rect 28 645 40 697
rect 92 645 164 697
rect 216 645 288 697
rect 340 645 412 697
rect 464 645 536 697
rect 588 645 660 697
rect 712 645 784 697
rect 836 645 908 697
rect 960 645 972 697
rect 28 573 972 645
rect 28 521 40 573
rect 92 521 164 573
rect 216 521 288 573
rect 340 521 412 573
rect 464 521 536 573
rect 588 521 660 573
rect 712 521 784 573
rect 836 521 908 573
rect 960 521 972 573
rect 28 449 972 521
rect 28 397 40 449
rect 92 397 164 449
rect 216 397 288 449
rect 340 397 412 449
rect 464 397 536 449
rect 588 397 660 449
rect 712 397 784 449
rect 836 397 908 449
rect 960 397 972 449
rect 28 325 972 397
rect 28 273 40 325
rect 92 273 164 325
rect 216 273 288 325
rect 340 273 412 325
rect 464 273 536 325
rect 588 273 660 325
rect 712 273 784 325
rect 836 273 908 325
rect 960 273 972 325
rect 28 201 972 273
rect 28 149 40 201
rect 92 149 164 201
rect 216 149 288 201
rect 340 149 412 201
rect 464 149 536 201
rect 588 149 660 201
rect 712 149 784 201
rect 836 149 908 201
rect 960 149 972 201
rect 28 77 972 149
rect 28 25 40 77
rect 92 25 164 77
rect 216 25 288 77
rect 340 25 412 77
rect 464 25 536 77
rect 588 25 660 77
rect 712 25 784 77
rect 836 25 908 77
rect 960 25 972 77
rect 28 13 972 25
<< via1 >>
rect 40 893 92 945
rect 164 893 216 945
rect 288 893 340 945
rect 412 893 464 945
rect 536 893 588 945
rect 660 893 712 945
rect 784 893 836 945
rect 908 893 960 945
rect 40 769 92 821
rect 164 769 216 821
rect 288 769 340 821
rect 412 769 464 821
rect 536 769 588 821
rect 660 769 712 821
rect 784 769 836 821
rect 908 769 960 821
rect 40 645 92 697
rect 164 645 216 697
rect 288 645 340 697
rect 412 645 464 697
rect 536 645 588 697
rect 660 645 712 697
rect 784 645 836 697
rect 908 645 960 697
rect 40 521 92 573
rect 164 521 216 573
rect 288 521 340 573
rect 412 521 464 573
rect 536 521 588 573
rect 660 521 712 573
rect 784 521 836 573
rect 908 521 960 573
rect 40 397 92 449
rect 164 397 216 449
rect 288 397 340 449
rect 412 397 464 449
rect 536 397 588 449
rect 660 397 712 449
rect 784 397 836 449
rect 908 397 960 449
rect 40 273 92 325
rect 164 273 216 325
rect 288 273 340 325
rect 412 273 464 325
rect 536 273 588 325
rect 660 273 712 325
rect 784 273 836 325
rect 908 273 960 325
rect 40 149 92 201
rect 164 149 216 201
rect 288 149 340 201
rect 412 149 464 201
rect 536 149 588 201
rect 660 149 712 201
rect 784 149 836 201
rect 908 149 960 201
rect 40 25 92 77
rect 164 25 216 77
rect 288 25 340 77
rect 412 25 464 77
rect 536 25 588 77
rect 660 25 712 77
rect 784 25 836 77
rect 908 25 960 77
<< metal2 >>
rect 0 945 1000 1000
rect 0 893 40 945
rect 92 893 164 945
rect 216 893 288 945
rect 340 893 412 945
rect 464 893 536 945
rect 588 893 660 945
rect 712 893 784 945
rect 836 893 908 945
rect 960 893 1000 945
rect 0 821 1000 893
rect 0 769 40 821
rect 92 769 164 821
rect 216 769 288 821
rect 340 769 412 821
rect 464 769 536 821
rect 588 769 660 821
rect 712 769 784 821
rect 836 769 908 821
rect 960 769 1000 821
rect 0 697 1000 769
rect 0 645 40 697
rect 92 645 164 697
rect 216 645 288 697
rect 340 645 412 697
rect 464 645 536 697
rect 588 645 660 697
rect 712 645 784 697
rect 836 645 908 697
rect 960 645 1000 697
rect 0 575 1000 645
rect 0 519 38 575
rect 94 519 162 575
rect 218 519 286 575
rect 342 519 410 575
rect 466 519 534 575
rect 590 519 658 575
rect 714 519 782 575
rect 838 519 906 575
rect 962 519 1000 575
rect 0 451 1000 519
rect 0 395 38 451
rect 94 395 162 451
rect 218 395 286 451
rect 342 395 410 451
rect 466 395 534 451
rect 590 395 658 451
rect 714 395 782 451
rect 838 395 906 451
rect 962 395 1000 451
rect 0 327 1000 395
rect 0 271 38 327
rect 94 271 162 327
rect 218 271 286 327
rect 342 271 410 327
rect 466 271 534 327
rect 590 271 658 327
rect 714 271 782 327
rect 838 271 906 327
rect 962 271 1000 327
rect 0 203 1000 271
rect 0 147 38 203
rect 94 147 162 203
rect 218 147 286 203
rect 342 147 410 203
rect 466 147 534 203
rect 590 147 658 203
rect 714 147 782 203
rect 838 147 906 203
rect 962 147 1000 203
rect 0 79 1000 147
rect 0 23 38 79
rect 94 23 162 79
rect 218 23 286 79
rect 342 23 410 79
rect 466 23 534 79
rect 590 23 658 79
rect 714 23 782 79
rect 838 23 906 79
rect 962 23 1000 79
rect 0 0 1000 23
<< via2 >>
rect 38 573 94 575
rect 38 521 40 573
rect 40 521 92 573
rect 92 521 94 573
rect 38 519 94 521
rect 162 573 218 575
rect 162 521 164 573
rect 164 521 216 573
rect 216 521 218 573
rect 162 519 218 521
rect 286 573 342 575
rect 286 521 288 573
rect 288 521 340 573
rect 340 521 342 573
rect 286 519 342 521
rect 410 573 466 575
rect 410 521 412 573
rect 412 521 464 573
rect 464 521 466 573
rect 410 519 466 521
rect 534 573 590 575
rect 534 521 536 573
rect 536 521 588 573
rect 588 521 590 573
rect 534 519 590 521
rect 658 573 714 575
rect 658 521 660 573
rect 660 521 712 573
rect 712 521 714 573
rect 658 519 714 521
rect 782 573 838 575
rect 782 521 784 573
rect 784 521 836 573
rect 836 521 838 573
rect 782 519 838 521
rect 906 573 962 575
rect 906 521 908 573
rect 908 521 960 573
rect 960 521 962 573
rect 906 519 962 521
rect 38 449 94 451
rect 38 397 40 449
rect 40 397 92 449
rect 92 397 94 449
rect 38 395 94 397
rect 162 449 218 451
rect 162 397 164 449
rect 164 397 216 449
rect 216 397 218 449
rect 162 395 218 397
rect 286 449 342 451
rect 286 397 288 449
rect 288 397 340 449
rect 340 397 342 449
rect 286 395 342 397
rect 410 449 466 451
rect 410 397 412 449
rect 412 397 464 449
rect 464 397 466 449
rect 410 395 466 397
rect 534 449 590 451
rect 534 397 536 449
rect 536 397 588 449
rect 588 397 590 449
rect 534 395 590 397
rect 658 449 714 451
rect 658 397 660 449
rect 660 397 712 449
rect 712 397 714 449
rect 658 395 714 397
rect 782 449 838 451
rect 782 397 784 449
rect 784 397 836 449
rect 836 397 838 449
rect 782 395 838 397
rect 906 449 962 451
rect 906 397 908 449
rect 908 397 960 449
rect 960 397 962 449
rect 906 395 962 397
rect 38 325 94 327
rect 38 273 40 325
rect 40 273 92 325
rect 92 273 94 325
rect 38 271 94 273
rect 162 325 218 327
rect 162 273 164 325
rect 164 273 216 325
rect 216 273 218 325
rect 162 271 218 273
rect 286 325 342 327
rect 286 273 288 325
rect 288 273 340 325
rect 340 273 342 325
rect 286 271 342 273
rect 410 325 466 327
rect 410 273 412 325
rect 412 273 464 325
rect 464 273 466 325
rect 410 271 466 273
rect 534 325 590 327
rect 534 273 536 325
rect 536 273 588 325
rect 588 273 590 325
rect 534 271 590 273
rect 658 325 714 327
rect 658 273 660 325
rect 660 273 712 325
rect 712 273 714 325
rect 658 271 714 273
rect 782 325 838 327
rect 782 273 784 325
rect 784 273 836 325
rect 836 273 838 325
rect 782 271 838 273
rect 906 325 962 327
rect 906 273 908 325
rect 908 273 960 325
rect 960 273 962 325
rect 906 271 962 273
rect 38 201 94 203
rect 38 149 40 201
rect 40 149 92 201
rect 92 149 94 201
rect 38 147 94 149
rect 162 201 218 203
rect 162 149 164 201
rect 164 149 216 201
rect 216 149 218 201
rect 162 147 218 149
rect 286 201 342 203
rect 286 149 288 201
rect 288 149 340 201
rect 340 149 342 201
rect 286 147 342 149
rect 410 201 466 203
rect 410 149 412 201
rect 412 149 464 201
rect 464 149 466 201
rect 410 147 466 149
rect 534 201 590 203
rect 534 149 536 201
rect 536 149 588 201
rect 588 149 590 201
rect 534 147 590 149
rect 658 201 714 203
rect 658 149 660 201
rect 660 149 712 201
rect 712 149 714 201
rect 658 147 714 149
rect 782 201 838 203
rect 782 149 784 201
rect 784 149 836 201
rect 836 149 838 201
rect 782 147 838 149
rect 906 201 962 203
rect 906 149 908 201
rect 908 149 960 201
rect 960 149 962 201
rect 906 147 962 149
rect 38 77 94 79
rect 38 25 40 77
rect 40 25 92 77
rect 92 25 94 77
rect 38 23 94 25
rect 162 77 218 79
rect 162 25 164 77
rect 164 25 216 77
rect 216 25 218 77
rect 162 23 218 25
rect 286 77 342 79
rect 286 25 288 77
rect 288 25 340 77
rect 340 25 342 77
rect 286 23 342 25
rect 410 77 466 79
rect 410 25 412 77
rect 412 25 464 77
rect 464 25 466 77
rect 410 23 466 25
rect 534 77 590 79
rect 534 25 536 77
rect 536 25 588 77
rect 588 25 590 77
rect 534 23 590 25
rect 658 77 714 79
rect 658 25 660 77
rect 660 25 712 77
rect 712 25 714 77
rect 658 23 714 25
rect 782 77 838 79
rect 782 25 784 77
rect 784 25 836 77
rect 836 25 838 77
rect 782 23 838 25
rect 906 77 962 79
rect 906 25 908 77
rect 908 25 960 77
rect 960 25 962 77
rect 906 23 962 25
<< metal3 >>
rect 0 575 1000 650
rect 0 519 38 575
rect 94 519 162 575
rect 218 519 286 575
rect 342 519 410 575
rect 466 519 534 575
rect 590 519 658 575
rect 714 519 782 575
rect 838 519 906 575
rect 962 519 1000 575
rect 0 451 1000 519
rect 0 395 38 451
rect 94 395 162 451
rect 218 395 286 451
rect 342 395 410 451
rect 466 395 534 451
rect 590 395 658 451
rect 714 395 782 451
rect 838 395 906 451
rect 962 395 1000 451
rect 0 327 1000 395
rect 0 271 38 327
rect 94 271 162 327
rect 218 271 286 327
rect 342 271 410 327
rect 466 271 534 327
rect 590 271 658 327
rect 714 271 782 327
rect 838 271 906 327
rect 962 271 1000 327
rect 0 203 1000 271
rect 0 147 38 203
rect 94 147 162 203
rect 218 147 286 203
rect 342 147 410 203
rect 466 147 534 203
rect 590 147 658 203
rect 714 147 782 203
rect 838 147 906 203
rect 962 147 1000 203
rect 0 79 1000 147
rect 0 23 38 79
rect 94 23 162 79
rect 218 23 286 79
rect 342 23 410 79
rect 466 23 534 79
rect 590 23 658 79
rect 714 23 782 79
rect 838 23 906 79
rect 962 23 1000 79
rect 0 -282 1000 23
use M2_M143105905487110_128x8m81  M2_M143105905487110_128x8m81_0
timestamp 1749760379
transform 1 0 500 0 1 485
box 0 0 1 1
use M3_M243105905487111_128x8m81  M3_M243105905487111_128x8m81_0
timestamp 1749760379
transform 1 0 500 0 1 299
box 0 0 1 1
<< properties >>
string GDS_END 2231532
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2231296
<< end >>
