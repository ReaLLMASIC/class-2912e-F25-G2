magic
tech gf180mcuD
magscale 1 5
timestamp 1749760379
use pmos_6p0_esd  pmos_6p0_esd_0
timestamp 1749760379
transform -1 0 1040 0 1 0
box 0 6 598 6126
use pmos_6p0_esd  pmos_6p0_esd_1
timestamp 1749760379
transform 1 0 0 0 1 0
box 0 6 598 6126
<< properties >>
string GDS_END 2653174
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2653080
<< end >>
