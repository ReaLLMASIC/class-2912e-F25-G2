magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
use M1_NACTIVE4310590548729_128x8m81  M1_NACTIVE4310590548729_128x8m81_0
timestamp 1749760379
transform 1 0 1937 0 1 7871
box 0 0 1 1
use M1_NACTIVE4310590548729_128x8m81  M1_NACTIVE4310590548729_128x8m81_1
timestamp 1749760379
transform 1 0 4414 0 1 7871
box 0 0 1 1
use M1_NACTIVE4310590548729_128x8m81  M1_NACTIVE4310590548729_128x8m81_2
timestamp 1749760379
transform 1 0 3175 0 1 7871
box 0 0 1 1
use M1_NACTIVE4310590548729_128x8m81  M1_NACTIVE4310590548729_128x8m81_3
timestamp 1749760379
transform 1 0 698 0 1 7871
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_0
timestamp 1749760379
transform 1 0 1318 0 1 513
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_1
timestamp 1749760379
transform 1 0 2557 0 1 513
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_2
timestamp 1749760379
transform 1 0 5034 0 1 513
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_3
timestamp 1749760379
transform 1 0 3795 0 1 513
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_4
timestamp 1749760379
transform 1 0 -9 0 1 513
box 0 0 1 1
use M1_PSUB$$45111340_128x8m81  M1_PSUB$$45111340_128x8m81_0
timestamp 1749760379
transform 1 0 1937 0 1 5328
box 0 0 1 1
use M1_PSUB$$45111340_128x8m81  M1_PSUB$$45111340_128x8m81_1
timestamp 1749760379
transform 1 0 698 0 1 5328
box 0 0 1 1
use M1_PSUB$$45111340_128x8m81  M1_PSUB$$45111340_128x8m81_2
timestamp 1749760379
transform 1 0 3175 0 1 5328
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_0
timestamp 1749760379
transform 1 0 1937 0 1 7885
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_1
timestamp 1749760379
transform 1 0 3175 0 1 7885
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_2
timestamp 1749760379
transform 1 0 4414 0 1 7885
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_3
timestamp 1749760379
transform 1 0 698 0 1 7885
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_0
timestamp 1749760379
transform 1 0 1463 0 1 1483
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_1
timestamp 1749760379
transform 1 0 2702 0 1 1483
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_2
timestamp 1749760379
transform 1 0 2411 0 1 1483
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_3
timestamp 1749760379
transform 1 0 3940 0 1 1483
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_4
timestamp 1749760379
transform 1 0 3649 0 1 1483
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_5
timestamp 1749760379
transform 1 0 1172 0 1 1483
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_0
timestamp 1749760379
transform 1 0 1463 0 1 1431
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_1
timestamp 1749760379
transform 1 0 2411 0 1 1431
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_2
timestamp 1749760379
transform 1 0 2702 0 1 1431
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_3
timestamp 1749760379
transform 1 0 3649 0 1 1431
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_4
timestamp 1749760379
transform 1 0 3940 0 1 1431
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_5
timestamp 1749760379
transform 1 0 1172 0 1 1431
box 0 0 1 1
use M3_M24310590548730_128x8m81  M3_M24310590548730_128x8m81_0
timestamp 1749760379
transform 1 0 698 0 1 7885
box 0 0 1 1
use M3_M24310590548730_128x8m81  M3_M24310590548730_128x8m81_1
timestamp 1749760379
transform 1 0 3175 0 1 7885
box 0 0 1 1
use M3_M24310590548730_128x8m81  M3_M24310590548730_128x8m81_2
timestamp 1749760379
transform 1 0 4414 0 1 7885
box 0 0 1 1
use M3_M24310590548730_128x8m81  M3_M24310590548730_128x8m81_3
timestamp 1749760379
transform 1 0 1937 0 1 7885
box 0 0 1 1
use ypass_gate_128x8m81  ypass_gate_128x8m81_0
timestamp 1749760379
transform -1 0 3175 0 1 91
box 0 73 527 12143
use ypass_gate_128x8m81  ypass_gate_128x8m81_1
timestamp 1749760379
transform -1 0 4414 0 1 91
box 0 73 527 12143
use ypass_gate_128x8m81  ypass_gate_128x8m81_2
timestamp 1749760379
transform -1 0 1937 0 1 91
box 0 73 527 12143
use ypass_gate_128x8m81  ypass_gate_128x8m81_3
timestamp 1749760379
transform -1 0 698 0 1 91
box 0 73 527 12143
use ypass_gate_128x8m81  ypass_gate_128x8m81_4
timestamp 1749760379
transform 1 0 3175 0 1 91
box 0 73 527 12143
use ypass_gate_128x8m81  ypass_gate_128x8m81_5
timestamp 1749760379
transform 1 0 1937 0 1 91
box 0 73 527 12143
use ypass_gate_128x8m81  ypass_gate_128x8m81_6
timestamp 1749760379
transform 1 0 698 0 1 91
box 0 73 527 12143
use ypass_gate_a_128x8m81  ypass_gate_a_128x8m81_0
timestamp 1749760379
transform 1 0 4414 0 1 91
box 0 73 621 12143
<< properties >>
string GDS_END 431884
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 428428
<< end >>
