magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 352 1430 870
<< pwell >>
rect -86 -86 1430 352
<< metal1 >>
rect 0 724 1344 844
rect 542 558 610 724
rect 176 512 465 546
rect 950 539 1208 585
rect 176 466 899 512
rect 176 338 312 466
rect 851 431 899 466
rect 375 364 803 420
rect 757 314 803 364
rect 851 360 1098 431
rect 757 268 905 314
rect 1144 222 1208 539
rect 38 60 106 152
rect 757 175 1208 222
rect 522 60 590 152
rect 757 106 803 175
rect 1154 60 1222 127
rect 0 -60 1344 60
<< obsm1 >>
rect 58 258 126 670
rect 718 631 1224 678
rect 634 258 702 311
rect 58 198 702 258
rect 262 106 330 198
<< labels >>
rlabel metal1 s 757 268 905 314 6 A1
port 1 nsew default input
rlabel metal1 s 757 314 803 364 6 A1
port 1 nsew default input
rlabel metal1 s 375 364 803 420 6 A1
port 1 nsew default input
rlabel metal1 s 851 360 1098 431 6 A2
port 2 nsew default input
rlabel metal1 s 851 431 899 466 6 A2
port 2 nsew default input
rlabel metal1 s 176 338 312 466 6 A2
port 2 nsew default input
rlabel metal1 s 176 466 899 512 6 A2
port 2 nsew default input
rlabel metal1 s 176 512 465 546 6 A2
port 2 nsew default input
rlabel metal1 s 757 106 803 175 6 Z
port 3 nsew default output
rlabel metal1 s 757 175 1208 222 6 Z
port 3 nsew default output
rlabel metal1 s 1144 222 1208 539 6 Z
port 3 nsew default output
rlabel metal1 s 950 539 1208 585 6 Z
port 3 nsew default output
rlabel metal1 s 542 558 610 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 724 1344 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel nwell s -86 352 1430 870 6 VNW
port 5 nsew power bidirectional
rlabel pwell s -86 -86 1430 352 6 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 0 -60 1344 60 8 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1154 60 1222 127 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 522 60 590 152 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 152 6 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1344 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 360014
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 356412
<< end >>
