magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 352 4790 870
<< pwell >>
rect -86 -86 4790 352
<< mvnmos >>
rect 124 124 244 232
rect 348 124 468 232
rect 720 156 840 232
rect 964 156 1084 232
rect 1188 156 1308 232
rect 1356 156 1476 232
rect 1588 156 1708 232
rect 1816 156 1936 232
rect 2040 156 2160 232
rect 2264 156 2384 232
rect 2888 145 3008 232
rect 3148 170 3268 232
rect 3416 157 3536 232
rect 3784 69 3904 232
rect 4008 69 4128 232
rect 4232 69 4352 232
rect 4456 69 4576 232
<< mvpmos >>
rect 144 472 244 660
rect 348 472 448 660
rect 740 472 840 593
rect 944 472 1044 593
rect 1148 472 1248 593
rect 1296 472 1396 593
rect 1588 472 1688 586
rect 1836 521 1936 647
rect 2264 472 2364 579
rect 2504 472 2604 602
rect 2908 507 3008 648
rect 3168 472 3268 588
rect 3424 472 3524 603
rect 3804 472 3904 715
rect 4008 472 4108 715
rect 4212 472 4312 715
rect 4416 472 4516 715
<< mvndiff >>
rect 36 189 124 232
rect 36 143 49 189
rect 95 143 124 189
rect 36 124 124 143
rect 244 187 348 232
rect 244 141 273 187
rect 319 141 348 187
rect 244 124 348 141
rect 468 189 556 232
rect 468 143 497 189
rect 543 143 556 189
rect 632 218 720 232
rect 632 172 645 218
rect 691 172 720 218
rect 632 156 720 172
rect 840 219 964 232
rect 840 173 869 219
rect 915 173 964 219
rect 840 156 964 173
rect 1084 219 1188 232
rect 1084 173 1113 219
rect 1159 173 1188 219
rect 1084 156 1188 173
rect 1308 156 1356 232
rect 1476 218 1588 232
rect 1476 172 1505 218
rect 1551 172 1588 218
rect 1476 156 1588 172
rect 1708 156 1816 232
rect 1936 219 2040 232
rect 1936 173 1965 219
rect 2011 173 2040 219
rect 1936 156 2040 173
rect 2160 219 2264 232
rect 2160 173 2189 219
rect 2235 173 2264 219
rect 2160 156 2264 173
rect 2384 215 2472 232
rect 2384 169 2413 215
rect 2459 169 2472 215
rect 2384 156 2472 169
rect 468 124 556 143
rect 2800 216 2888 232
rect 2800 170 2813 216
rect 2859 170 2888 216
rect 2800 145 2888 170
rect 3008 170 3148 232
rect 3268 216 3416 232
rect 3268 170 3341 216
rect 3387 170 3416 216
rect 3008 145 3088 170
rect 3328 157 3416 170
rect 3536 216 3624 232
rect 3536 170 3565 216
rect 3611 170 3624 216
rect 3536 157 3624 170
rect 3696 142 3784 232
rect 3696 96 3709 142
rect 3755 96 3784 142
rect 3696 69 3784 96
rect 3904 218 4008 232
rect 3904 172 3933 218
rect 3979 172 4008 218
rect 3904 69 4008 172
rect 4128 142 4232 232
rect 4128 96 4157 142
rect 4203 96 4232 142
rect 4128 69 4232 96
rect 4352 213 4456 232
rect 4352 167 4381 213
rect 4427 167 4456 213
rect 4352 69 4456 167
rect 4576 142 4664 232
rect 4576 96 4605 142
rect 4651 96 4664 142
rect 4576 69 4664 96
<< mvpdiff >>
rect 56 647 144 660
rect 56 507 69 647
rect 115 507 144 647
rect 56 472 144 507
rect 244 647 348 660
rect 244 601 273 647
rect 319 601 348 647
rect 244 472 348 601
rect 448 647 536 660
rect 448 507 477 647
rect 523 507 536 647
rect 448 472 536 507
rect 608 647 680 660
rect 608 601 621 647
rect 667 601 680 647
rect 608 593 680 601
rect 1456 694 1528 707
rect 1456 648 1469 694
rect 1515 648 1528 694
rect 1456 593 1528 648
rect 608 472 740 593
rect 840 550 944 593
rect 840 504 869 550
rect 915 504 944 550
rect 840 472 944 504
rect 1044 531 1148 593
rect 1044 485 1073 531
rect 1119 485 1148 531
rect 1044 472 1148 485
rect 1248 472 1296 593
rect 1396 586 1528 593
rect 1756 586 1836 647
rect 1396 472 1588 586
rect 1688 531 1836 586
rect 1688 485 1717 531
rect 1763 521 1836 531
rect 1936 634 2024 647
rect 1936 588 1965 634
rect 2011 588 2024 634
rect 1936 521 2024 588
rect 3716 665 3804 715
rect 2820 635 2908 648
rect 2424 579 2504 602
rect 2176 531 2264 579
rect 1763 485 1776 521
rect 1688 472 1776 485
rect 2176 485 2189 531
rect 2235 485 2264 531
rect 2176 472 2264 485
rect 2364 531 2504 579
rect 2364 485 2429 531
rect 2475 485 2504 531
rect 2364 472 2504 485
rect 2604 531 2692 602
rect 2604 485 2633 531
rect 2679 485 2692 531
rect 2820 589 2833 635
rect 2879 589 2908 635
rect 2820 507 2908 589
rect 3008 588 3096 648
rect 3336 588 3424 603
rect 3008 531 3168 588
rect 3008 507 3089 531
rect 2604 472 2692 485
rect 3076 485 3089 507
rect 3135 485 3168 531
rect 3076 472 3168 485
rect 3268 577 3424 588
rect 3268 531 3349 577
rect 3395 531 3424 577
rect 3268 472 3424 531
rect 3524 535 3612 603
rect 3524 489 3553 535
rect 3599 489 3612 535
rect 3524 472 3612 489
rect 3716 525 3729 665
rect 3775 525 3804 665
rect 3716 472 3804 525
rect 3904 665 4008 715
rect 3904 525 3933 665
rect 3979 525 4008 665
rect 3904 472 4008 525
rect 4108 665 4212 715
rect 4108 525 4137 665
rect 4183 525 4212 665
rect 4108 472 4212 525
rect 4312 665 4416 715
rect 4312 525 4341 665
rect 4387 525 4416 665
rect 4312 472 4416 525
rect 4516 665 4604 715
rect 4516 525 4545 665
rect 4591 525 4604 665
rect 4516 472 4604 525
<< mvndiffc >>
rect 49 143 95 189
rect 273 141 319 187
rect 497 143 543 189
rect 645 172 691 218
rect 869 173 915 219
rect 1113 173 1159 219
rect 1505 172 1551 218
rect 1965 173 2011 219
rect 2189 173 2235 219
rect 2413 169 2459 215
rect 2813 170 2859 216
rect 3341 170 3387 216
rect 3565 170 3611 216
rect 3709 96 3755 142
rect 3933 172 3979 218
rect 4157 96 4203 142
rect 4381 167 4427 213
rect 4605 96 4651 142
<< mvpdiffc >>
rect 69 507 115 647
rect 273 601 319 647
rect 477 507 523 647
rect 621 601 667 647
rect 1469 648 1515 694
rect 869 504 915 550
rect 1073 485 1119 531
rect 1717 485 1763 531
rect 1965 588 2011 634
rect 2189 485 2235 531
rect 2429 485 2475 531
rect 2633 485 2679 531
rect 2833 589 2879 635
rect 3089 485 3135 531
rect 3349 531 3395 577
rect 3553 489 3599 535
rect 3729 525 3775 665
rect 3933 525 3979 665
rect 4137 525 4183 665
rect 4341 525 4387 665
rect 4545 525 4591 665
<< polysilicon >>
rect 348 720 1044 760
rect 144 660 244 705
rect 348 660 448 720
rect 740 593 840 637
rect 944 593 1044 720
rect 1836 720 3008 760
rect 1148 672 1248 685
rect 1148 626 1189 672
rect 1235 626 1248 672
rect 1148 593 1248 626
rect 1296 593 1396 637
rect 1836 647 1936 720
rect 2264 659 2364 672
rect 1588 586 1688 630
rect 2264 613 2277 659
rect 2323 613 2364 659
rect 2908 648 3008 720
rect 3804 715 3904 760
rect 4008 715 4108 760
rect 4212 715 4312 760
rect 4416 715 4516 760
rect 2264 579 2364 613
rect 2504 602 2604 646
rect 144 410 244 472
rect 144 364 157 410
rect 203 364 244 410
rect 144 288 244 364
rect 124 232 244 288
rect 348 326 448 472
rect 348 280 385 326
rect 431 288 448 326
rect 740 415 840 472
rect 944 428 1044 472
rect 740 369 753 415
rect 799 369 840 415
rect 1148 376 1248 472
rect 431 280 468 288
rect 348 232 468 280
rect 740 276 840 369
rect 720 232 840 276
rect 964 336 1248 376
rect 1296 439 1396 472
rect 1296 393 1337 439
rect 1383 393 1396 439
rect 1296 336 1396 393
rect 964 232 1084 336
rect 1356 314 1396 336
rect 1588 326 1688 472
rect 1188 232 1308 276
rect 1356 232 1476 314
rect 1588 280 1601 326
rect 1647 280 1688 326
rect 1588 276 1688 280
rect 1836 276 1936 521
rect 3168 588 3268 632
rect 3424 603 3524 648
rect 2264 276 2364 472
rect 2504 392 2604 472
rect 2504 304 2632 392
rect 1588 232 1708 276
rect 1816 232 1936 276
rect 2040 232 2160 276
rect 2264 232 2384 276
rect 124 80 244 124
rect 348 64 468 124
rect 720 112 840 156
rect 964 112 1084 156
rect 1188 64 1308 156
rect 1356 112 1476 156
rect 1588 112 1708 156
rect 1816 112 1936 156
rect 2040 64 2160 156
rect 2264 112 2384 156
rect 2532 64 2632 304
rect 2908 323 3008 507
rect 2908 288 2942 323
rect 2888 277 2942 288
rect 2988 277 3008 323
rect 3168 323 3268 472
rect 3168 288 3209 323
rect 2888 232 3008 277
rect 3148 277 3209 288
rect 3255 277 3268 323
rect 3424 439 3524 472
rect 3424 393 3437 439
rect 3483 393 3524 439
rect 3424 288 3524 393
rect 3804 367 3904 472
rect 3804 321 3817 367
rect 3863 344 3904 367
rect 4008 367 4108 472
rect 4008 344 4037 367
rect 3863 321 4037 344
rect 4083 344 4108 367
rect 4212 367 4312 472
rect 4212 344 4239 367
rect 4083 321 4239 344
rect 4285 344 4312 367
rect 4416 344 4516 472
rect 4285 321 4516 344
rect 3804 304 4516 321
rect 3804 288 3904 304
rect 3148 232 3268 277
rect 3416 232 3536 288
rect 3784 232 3904 288
rect 4008 232 4128 304
rect 4232 232 4352 304
rect 4456 288 4516 304
rect 4456 232 4576 288
rect 2888 101 3008 145
rect 3148 126 3268 170
rect 3416 101 3536 157
rect 348 24 2632 64
rect 3784 24 3904 69
rect 4008 24 4128 69
rect 4232 24 4352 69
rect 4456 24 4576 69
<< polycontact >>
rect 1189 626 1235 672
rect 2277 613 2323 659
rect 157 364 203 410
rect 385 280 431 326
rect 753 369 799 415
rect 1337 393 1383 439
rect 1601 280 1647 326
rect 2942 277 2988 323
rect 3209 277 3255 323
rect 3437 393 3483 439
rect 3817 321 3863 367
rect 4037 321 4083 367
rect 4239 321 4285 367
<< metal1 >>
rect 0 724 4704 844
rect 69 647 115 660
rect 262 647 330 724
rect 262 601 273 647
rect 319 601 330 647
rect 477 647 543 660
rect 115 507 431 519
rect 69 472 431 507
rect 56 410 318 426
rect 56 364 157 410
rect 203 364 318 410
rect 56 354 318 364
rect 385 326 431 472
rect 385 279 431 280
rect 49 233 431 279
rect 523 555 543 647
rect 610 647 678 724
rect 1458 694 1526 724
rect 610 601 621 647
rect 667 601 678 647
rect 724 626 1189 672
rect 1235 626 1246 672
rect 1458 648 1469 694
rect 1515 648 1526 694
rect 724 624 1246 626
rect 724 555 770 624
rect 523 509 770 555
rect 1188 576 1246 624
rect 1965 634 2011 724
rect 1595 577 1866 623
rect 1965 577 2011 588
rect 2057 613 2277 659
rect 2323 613 2334 659
rect 2822 635 2890 724
rect 1595 576 1641 577
rect 523 507 543 509
rect 49 189 95 233
rect 477 189 543 507
rect 858 504 869 550
rect 915 504 1018 550
rect 690 415 878 430
rect 690 369 753 415
rect 799 369 878 415
rect 690 354 878 369
rect 49 132 95 143
rect 262 141 273 187
rect 319 141 330 187
rect 262 60 330 141
rect 477 143 497 189
rect 477 132 543 143
rect 645 218 691 229
rect 972 219 1018 504
rect 858 173 869 219
rect 915 173 1018 219
rect 1073 531 1119 542
rect 1188 530 1641 576
rect 1820 531 1866 577
rect 2057 531 2103 613
rect 2429 588 2771 635
rect 2822 589 2833 635
rect 2879 589 2890 635
rect 2429 531 2475 588
rect 2725 543 2771 588
rect 2951 577 3276 624
rect 2951 543 2997 577
rect 1073 326 1119 485
rect 1706 485 1717 531
rect 1763 485 1774 531
rect 1820 485 2103 531
rect 2178 485 2189 531
rect 2235 485 2246 531
rect 1706 439 1774 485
rect 2178 439 2246 485
rect 1326 393 1337 439
rect 1383 393 2246 439
rect 1965 386 2246 393
rect 1073 280 1601 326
rect 1647 280 1658 326
rect 1073 279 1658 280
rect 1073 219 1170 279
rect 1073 173 1113 219
rect 1159 173 1170 219
rect 1965 219 2011 386
rect 2429 317 2475 485
rect 645 60 691 172
rect 1494 172 1505 218
rect 1551 172 1562 218
rect 1494 60 1562 172
rect 1965 162 2011 173
rect 2189 271 2475 317
rect 2633 531 2679 542
rect 2725 496 2997 543
rect 2633 439 2679 485
rect 3076 485 3089 531
rect 3135 485 3146 531
rect 3076 439 3146 485
rect 2633 393 3146 439
rect 3230 439 3276 577
rect 3349 577 3395 724
rect 3729 665 3775 724
rect 3349 520 3395 531
rect 3553 535 3599 575
rect 3729 514 3775 525
rect 3933 665 3979 676
rect 3230 393 3437 439
rect 3483 393 3494 439
rect 2189 219 2235 271
rect 2633 227 2679 393
rect 3230 392 3494 393
rect 3553 368 3599 489
rect 3933 464 3979 525
rect 4137 665 4183 724
rect 4137 514 4183 525
rect 4338 665 4462 676
rect 4338 525 4341 665
rect 4387 525 4462 665
rect 4338 464 4462 525
rect 4545 665 4591 724
rect 4545 514 4591 525
rect 3933 418 4462 464
rect 3553 367 4312 368
rect 2912 323 3118 334
rect 3553 323 3817 367
rect 2912 277 2942 323
rect 2988 277 3118 323
rect 3198 277 3209 323
rect 3255 321 3817 323
rect 3863 321 4037 367
rect 4083 321 4239 367
rect 4285 321 4312 367
rect 3255 277 3611 321
rect 2912 244 3118 277
rect 2633 216 2859 227
rect 3565 216 3611 277
rect 4386 258 4462 418
rect 2633 215 2813 216
rect 2189 162 2235 173
rect 2402 169 2413 215
rect 2459 170 2813 215
rect 2459 169 2859 170
rect 2402 159 2859 169
rect 3330 170 3341 216
rect 3387 170 3398 216
rect 3330 60 3398 170
rect 3565 159 3611 170
rect 3933 218 4462 258
rect 3979 213 4462 218
rect 3979 212 4381 213
rect 3933 161 3979 172
rect 4427 167 4462 213
rect 3709 142 3755 153
rect 3709 60 3755 96
rect 4157 142 4203 153
rect 4381 110 4462 167
rect 4605 142 4651 153
rect 4157 60 4203 96
rect 4605 60 4651 96
rect 0 -60 4704 60
<< labels >>
flabel metal1 s 690 354 878 430 0 FreeSans 600 0 0 0 D
port 1 nsew default input
flabel metal1 s 4338 464 4462 676 0 FreeSans 600 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2912 244 3118 334 0 FreeSans 600 0 0 0 SETN
port 2 nsew default input
flabel metal1 s 0 724 4704 844 0 FreeSans 600 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 645 218 691 229 0 FreeSans 600 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 56 354 318 426 0 FreeSans 600 0 0 0 CLKN
port 3 nsew clock input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 3933 464 3979 676 1 Q
port 4 nsew default output
rlabel metal1 s 3933 418 4462 464 1 Q
port 4 nsew default output
rlabel metal1 s 4386 258 4462 418 1 Q
port 4 nsew default output
rlabel metal1 s 3933 212 4462 258 1 Q
port 4 nsew default output
rlabel metal1 s 4381 161 4462 212 1 Q
port 4 nsew default output
rlabel metal1 s 3933 161 3979 212 1 Q
port 4 nsew default output
rlabel metal1 s 4381 110 4462 161 1 Q
port 4 nsew default output
rlabel metal1 s 4545 648 4591 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4137 648 4183 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3729 648 3775 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 648 3395 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2822 648 2890 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1965 648 2011 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1458 648 1526 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 610 648 678 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 262 648 330 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4545 601 4591 648 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4137 601 4183 648 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3729 601 3775 648 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 601 3395 648 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2822 601 2890 648 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1965 601 2011 648 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 610 601 678 648 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 262 601 330 648 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4545 589 4591 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4137 589 4183 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3729 589 3775 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 589 3395 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2822 589 2890 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1965 589 2011 601 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4545 577 4591 589 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4137 577 4183 589 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3729 577 3775 589 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 577 3395 589 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1965 577 2011 589 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4545 520 4591 577 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4137 520 4183 577 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3729 520 3775 577 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 520 3395 577 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4545 514 4591 520 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4137 514 4183 520 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3729 514 3775 520 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1494 216 1562 218 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 645 216 691 218 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3330 187 3398 216 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1494 187 1562 216 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 645 187 691 216 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3330 153 3398 187 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1494 153 1562 187 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 645 153 691 187 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 153 330 187 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4605 60 4651 153 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4157 60 4203 153 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3709 60 3755 153 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3330 60 3398 153 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1494 60 1562 153 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 645 60 691 153 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 153 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4704 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4704 784
string GDS_END 967302
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 957954
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
