magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< deepnwell >>
rect -680 -680 788 1080
<< pbase >>
rect -180 -180 288 580
<< ndiff >>
rect 0 363 108 400
rect 0 35 31 363
rect 77 35 108 363
rect 0 0 108 35
<< ndiffc >>
rect 31 35 77 363
<< psubdiff >>
rect -1264 1645 1372 1664
rect -1264 1599 -1097 1645
rect 1205 1599 1372 1645
rect -1264 1580 1372 1599
rect -1264 1492 -1180 1580
rect -1264 -1092 -1245 1492
rect -1199 -1092 -1180 1492
rect 1288 1492 1372 1580
rect -148 529 256 548
rect -148 483 -109 529
rect 219 483 256 529
rect -148 464 256 483
rect -148 419 -64 464
rect -148 -97 -129 419
rect -83 -64 -64 419
rect 172 419 256 464
rect 172 -64 191 419
rect -83 -97 191 -64
rect 237 -97 256 419
rect -148 -148 256 -97
rect -1264 -1180 -1180 -1092
rect 1288 -1092 1307 1492
rect 1353 -1092 1372 1492
rect 1288 -1180 1372 -1092
rect -1264 -1199 1372 -1180
rect -1264 -1245 -1097 -1199
rect -769 -1245 877 -1199
rect 1205 -1245 1372 -1199
rect -1264 -1264 1372 -1245
<< nsubdiff >>
rect -296 677 404 696
rect -296 631 -251 677
rect 359 631 404 677
rect -296 612 404 631
rect -296 557 -212 612
rect -296 -241 -277 557
rect -231 -212 -212 557
rect 320 557 404 612
rect 320 -212 339 557
rect -231 -241 339 -212
rect 385 -241 404 557
rect -296 -296 404 -241
<< psubdiffcont >>
rect -1097 1599 1205 1645
rect -1245 -1092 -1199 1492
rect -109 483 219 529
rect -129 -97 -83 419
rect 191 -97 237 419
rect 1307 -1092 1353 1492
rect -1097 -1245 -769 -1199
rect 877 -1245 1205 -1199
<< nsubdiffcont >>
rect -251 631 359 677
rect -277 -241 -231 557
rect 339 -241 385 557
<< metal1 >>
rect -1264 1645 1372 1664
rect -1264 1599 -1097 1645
rect 1205 1599 1372 1645
rect -1264 1580 1372 1599
rect -1264 1492 -1180 1580
rect -1264 -1092 -1245 1492
rect -1199 -1092 -1180 1492
rect 1288 1492 1372 1580
rect -296 677 404 696
rect -296 631 -251 677
rect 359 631 404 677
rect -296 612 404 631
rect -296 557 -212 612
rect -296 -241 -277 557
rect -231 -241 -212 557
rect 320 557 404 612
rect -148 529 256 548
rect -148 483 -109 529
rect 219 483 256 529
rect -148 464 256 483
rect -148 419 -64 464
rect -148 -97 -129 419
rect -83 -97 -64 419
rect 172 419 256 464
rect 0 363 108 400
rect 0 35 31 363
rect 77 35 108 363
rect 0 0 108 35
rect -148 -148 -64 -97
rect 172 -97 191 419
rect 237 -97 256 419
rect 172 -148 256 -97
rect -296 -296 -212 -241
rect 320 -241 339 557
rect 385 -241 404 557
rect 320 -296 404 -241
rect -1264 -1180 -1180 -1092
rect 1288 -1092 1307 1492
rect 1353 -1092 1372 1492
rect 1288 -1180 1372 -1092
rect -1264 -1199 -680 -1180
rect -1264 -1245 -1097 -1199
rect -769 -1245 -680 -1199
rect -1264 -1264 -680 -1245
rect 788 -1199 1372 -1180
rect 788 -1245 877 -1199
rect 1205 -1245 1372 -1199
rect 788 -1264 1372 -1245
<< labels >>
flabel ndiffc 50 199 50 199 0 FreeSans 400 0 0 0 E
flabel psubdiffcont -104 506 -104 506 0 FreeSans 400 0 0 0 B
flabel metal1 211 -106 211 -106 0 FreeSans 400 0 0 0 B
flabel psubdiffcont 212 507 212 507 0 FreeSans 400 0 0 0 B
flabel metal1 -255 654 -255 654 0 FreeSans 400 0 0 0 C
flabel metal1 365 -253 365 -253 0 FreeSans 400 0 0 0 C
flabel metal1 367 652 367 652 0 FreeSans 400 0 0 0 C
flabel metal1 -1218 -1223 -1218 -1223 0 FreeSans 400 0 0 0 S
flabel metal1 -1218 -1223 -1218 -1223 0 FreeSans 400 0 0 0 S
flabel metal1 1327 -1214 1327 -1214 0 FreeSans 400 0 0 0 S
flabel metal1 1327 -1214 1327 -1214 0 FreeSans 400 0 0 0 S
flabel metal1 1331 1627 1331 1627 0 FreeSans 400 0 0 0 S
<< properties >>
string GDS_END 11884
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/npn_00p54x02p00.gds
string GDS_START 112
string gencell npn_00p54x02p00
string library gf180mcu
string parameter m=1
<< end >>
