magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 453 4678 1094
<< pwell >>
rect -86 -86 4678 453
<< mvnmos >>
rect 124 187 244 303
rect 348 187 468 303
rect 516 187 636 303
rect 740 187 860 303
rect 908 187 1028 303
rect 1308 166 1428 324
rect 1532 166 1652 324
rect 1900 185 2020 301
rect 2124 185 2244 301
rect 2292 185 2412 301
rect 2460 185 2580 301
rect 2772 185 2892 301
rect 2996 185 3116 301
rect 3220 185 3340 301
rect 3491 185 3611 301
rect 3715 185 3835 301
rect 3899 185 4019 301
rect 4285 69 4405 333
<< mvpmos >>
rect 134 652 234 852
rect 348 652 448 852
rect 496 652 596 852
rect 740 652 840 852
rect 888 652 988 852
rect 1318 589 1418 865
rect 1532 589 1632 865
rect 1894 652 1994 852
rect 2098 652 2198 852
rect 2302 652 2402 852
rect 2506 652 2606 852
rect 2866 652 2966 852
rect 3070 652 3170 852
rect 3307 652 3407 852
rect 3511 652 3611 852
rect 3715 652 3815 852
rect 3919 652 4019 852
rect 4295 574 4395 940
<< mvndiff >>
rect 36 246 124 303
rect 36 200 49 246
rect 95 200 124 246
rect 36 187 124 200
rect 244 246 348 303
rect 244 200 273 246
rect 319 200 348 246
rect 244 187 348 200
rect 468 187 516 303
rect 636 246 740 303
rect 636 200 665 246
rect 711 200 740 246
rect 636 187 740 200
rect 860 187 908 303
rect 1028 187 1148 303
rect 1088 108 1148 187
rect 1220 299 1308 324
rect 1220 253 1233 299
rect 1279 253 1308 299
rect 1220 166 1308 253
rect 1428 225 1532 324
rect 1428 179 1457 225
rect 1503 179 1532 225
rect 1428 166 1532 179
rect 1652 285 1740 324
rect 4197 320 4285 333
rect 1652 239 1681 285
rect 1727 239 1740 285
rect 1652 166 1740 239
rect 1812 244 1900 301
rect 1812 198 1825 244
rect 1871 198 1900 244
rect 1812 185 1900 198
rect 2020 246 2124 301
rect 2020 200 2049 246
rect 2095 200 2124 246
rect 2020 185 2124 200
rect 2244 185 2292 301
rect 2412 185 2460 301
rect 2580 277 2772 301
rect 2580 231 2653 277
rect 2699 231 2772 277
rect 2580 185 2772 231
rect 2892 288 2996 301
rect 2892 242 2921 288
rect 2967 242 2996 288
rect 2892 185 2996 242
rect 3116 288 3220 301
rect 3116 242 3145 288
rect 3191 242 3220 288
rect 3116 185 3220 242
rect 3340 288 3491 301
rect 3340 242 3416 288
rect 3462 242 3491 288
rect 3340 185 3491 242
rect 3611 244 3715 301
rect 3611 198 3640 244
rect 3686 198 3715 244
rect 3611 185 3715 198
rect 3835 185 3899 301
rect 4019 246 4107 301
rect 4019 200 4048 246
rect 4094 200 4107 246
rect 4019 185 4107 200
rect 1077 100 1148 108
rect 1077 95 1149 100
rect 1077 49 1090 95
rect 1136 49 1149 95
rect 1077 36 1149 49
rect 4197 180 4210 320
rect 4256 180 4285 320
rect 4197 69 4285 180
rect 4405 320 4493 333
rect 4405 180 4434 320
rect 4480 180 4493 320
rect 4405 69 4493 180
<< mvpdiff >>
rect 46 839 134 852
rect 46 699 59 839
rect 105 699 134 839
rect 46 652 134 699
rect 234 839 348 852
rect 234 699 263 839
rect 309 699 348 839
rect 234 652 348 699
rect 448 652 496 852
rect 596 839 740 852
rect 596 699 665 839
rect 711 699 740 839
rect 596 652 740 699
rect 840 652 888 852
rect 988 839 1076 852
rect 988 699 1017 839
rect 1063 699 1076 839
rect 988 652 1076 699
rect 1230 648 1318 865
rect 1230 602 1243 648
rect 1289 602 1318 648
rect 1230 589 1318 602
rect 1418 852 1532 865
rect 1418 806 1447 852
rect 1493 806 1532 852
rect 1418 589 1532 806
rect 1632 648 1720 865
rect 1806 751 1894 852
rect 1806 705 1819 751
rect 1865 705 1894 751
rect 1806 652 1894 705
rect 1994 839 2098 852
rect 1994 699 2023 839
rect 2069 699 2098 839
rect 1994 652 2098 699
rect 2198 839 2302 852
rect 2198 699 2227 839
rect 2273 699 2302 839
rect 2198 652 2302 699
rect 2402 839 2506 852
rect 2402 793 2431 839
rect 2477 793 2506 839
rect 2402 652 2506 793
rect 2606 839 2694 852
rect 2606 699 2635 839
rect 2681 699 2694 839
rect 2606 652 2694 699
rect 2778 839 2866 852
rect 2778 699 2791 839
rect 2837 699 2866 839
rect 2778 652 2866 699
rect 2966 839 3070 852
rect 2966 699 2995 839
rect 3041 699 3070 839
rect 2966 652 3070 699
rect 3170 839 3307 852
rect 3170 699 3199 839
rect 3245 699 3307 839
rect 3170 652 3307 699
rect 3407 745 3511 852
rect 3407 699 3436 745
rect 3482 699 3511 745
rect 3407 652 3511 699
rect 3611 839 3715 852
rect 3611 793 3640 839
rect 3686 793 3715 839
rect 3611 652 3715 793
rect 3815 745 3919 852
rect 3815 699 3844 745
rect 3890 699 3919 745
rect 3815 652 3919 699
rect 4019 839 4107 852
rect 4019 699 4048 839
rect 4094 699 4107 839
rect 4019 652 4107 699
rect 4207 839 4295 940
rect 4207 699 4220 839
rect 4266 699 4295 839
rect 1632 602 1661 648
rect 1707 602 1720 648
rect 1632 589 1720 602
rect 4207 574 4295 699
rect 4395 839 4483 940
rect 4395 699 4424 839
rect 4470 699 4483 839
rect 4395 574 4483 699
<< mvndiffc >>
rect 49 200 95 246
rect 273 200 319 246
rect 665 200 711 246
rect 1233 253 1279 299
rect 1457 179 1503 225
rect 1681 239 1727 285
rect 1825 198 1871 244
rect 2049 200 2095 246
rect 2653 231 2699 277
rect 2921 242 2967 288
rect 3145 242 3191 288
rect 3416 242 3462 288
rect 3640 198 3686 244
rect 4048 200 4094 246
rect 1090 49 1136 95
rect 4210 180 4256 320
rect 4434 180 4480 320
<< mvpdiffc >>
rect 59 699 105 839
rect 263 699 309 839
rect 665 699 711 839
rect 1017 699 1063 839
rect 1243 602 1289 648
rect 1447 806 1493 852
rect 1819 705 1865 751
rect 2023 699 2069 839
rect 2227 699 2273 839
rect 2431 793 2477 839
rect 2635 699 2681 839
rect 2791 699 2837 839
rect 2995 699 3041 839
rect 3199 699 3245 839
rect 3436 699 3482 745
rect 3640 793 3686 839
rect 3844 699 3890 745
rect 4048 699 4094 839
rect 4220 699 4266 839
rect 1661 602 1707 648
rect 4424 699 4470 839
<< polysilicon >>
rect 134 944 988 984
rect 134 852 234 944
rect 348 852 448 896
rect 496 852 596 896
rect 740 852 840 896
rect 888 852 988 944
rect 1532 944 3170 984
rect 1318 865 1418 909
rect 1532 865 1632 944
rect 134 529 234 652
rect 124 516 234 529
rect 124 470 137 516
rect 183 470 234 516
rect 124 347 234 470
rect 348 516 448 652
rect 348 470 361 516
rect 407 470 448 516
rect 348 347 448 470
rect 496 516 596 652
rect 496 470 509 516
rect 555 470 596 516
rect 496 457 596 470
rect 740 516 840 652
rect 888 608 988 652
rect 1894 852 1994 896
rect 2098 852 2198 944
rect 2302 852 2402 896
rect 2506 852 2606 896
rect 2866 852 2966 896
rect 3070 852 3170 944
rect 4295 940 4395 984
rect 3307 852 3407 896
rect 3511 852 3611 896
rect 3715 852 3815 896
rect 3919 852 4019 896
rect 1318 529 1418 589
rect 740 470 753 516
rect 799 470 840 516
rect 740 347 840 470
rect 908 516 1028 529
rect 908 470 921 516
rect 967 470 1028 516
rect 124 303 244 347
rect 348 303 468 347
rect 516 303 636 347
rect 740 303 860 347
rect 908 303 1028 470
rect 1308 516 1418 529
rect 1308 470 1321 516
rect 1367 470 1418 516
rect 1308 368 1418 470
rect 1532 516 1632 589
rect 1532 470 1545 516
rect 1591 470 1632 516
rect 1532 457 1632 470
rect 1894 529 1994 652
rect 2098 608 2198 652
rect 2302 529 2402 652
rect 2506 608 2606 652
rect 1894 516 2244 529
rect 1894 470 1907 516
rect 1953 470 2165 516
rect 2211 470 2244 516
rect 1894 457 2244 470
rect 1532 368 1572 457
rect 1308 324 1428 368
rect 1532 324 1652 368
rect 124 64 244 187
rect 348 143 468 187
rect 516 64 636 187
rect 740 143 860 187
rect 908 143 1028 187
rect 1900 301 2020 345
rect 2124 301 2244 457
rect 2302 516 2412 529
rect 2302 470 2353 516
rect 2399 470 2412 516
rect 2302 345 2412 470
rect 2506 345 2580 608
rect 2866 577 2966 652
rect 2292 301 2412 345
rect 2460 301 2580 345
rect 2772 564 2966 577
rect 2772 518 2805 564
rect 2851 518 2966 564
rect 2772 509 2966 518
rect 3070 550 3170 652
rect 3307 619 3407 652
rect 3307 573 3320 619
rect 3366 573 3407 619
rect 3307 560 3407 573
rect 2772 301 2892 509
rect 3070 478 3260 550
rect 2996 380 3116 393
rect 2996 334 3013 380
rect 3059 334 3116 380
rect 2996 301 3116 334
rect 3220 345 3260 478
rect 3511 516 3611 652
rect 3511 470 3552 516
rect 3598 470 3611 516
rect 3511 345 3611 470
rect 3220 301 3340 345
rect 3491 301 3611 345
rect 3715 516 3815 652
rect 3715 470 3728 516
rect 3774 470 3815 516
rect 3715 345 3815 470
rect 3919 516 4019 652
rect 3919 470 3936 516
rect 3982 470 4019 516
rect 3919 345 4019 470
rect 4067 516 4167 529
rect 4067 470 4080 516
rect 4126 514 4167 516
rect 4295 514 4395 574
rect 4126 470 4395 514
rect 4067 442 4395 470
rect 3715 301 3835 345
rect 3899 301 4019 345
rect 4285 377 4395 442
rect 4285 333 4405 377
rect 1308 122 1428 166
rect 124 24 636 64
rect 1532 96 1652 166
rect 1900 96 2020 185
rect 2124 141 2244 185
rect 2292 141 2412 185
rect 1532 24 2020 96
rect 2460 64 2580 185
rect 2772 141 2892 185
rect 2996 141 3116 185
rect 3220 141 3340 185
rect 3491 141 3611 185
rect 3715 64 3835 185
rect 3899 141 4019 185
rect 2460 24 3835 64
rect 4285 25 4405 69
<< polycontact >>
rect 137 470 183 516
rect 361 470 407 516
rect 509 470 555 516
rect 753 470 799 516
rect 921 470 967 516
rect 1321 470 1367 516
rect 1545 470 1591 516
rect 1907 470 1953 516
rect 2165 470 2211 516
rect 2353 470 2399 516
rect 2805 518 2851 564
rect 3320 573 3366 619
rect 3013 334 3059 380
rect 3552 470 3598 516
rect 3728 470 3774 516
rect 3936 470 3982 516
rect 4080 470 4126 516
<< metal1 >>
rect 0 918 4592 1098
rect 59 839 105 850
rect 59 642 105 699
rect 263 839 309 918
rect 263 688 309 699
rect 665 839 711 850
rect 665 642 711 699
rect 1017 839 1063 918
rect 1436 852 1504 918
rect 1436 806 1447 852
rect 1493 806 1504 852
rect 2023 839 2069 850
rect 1017 688 1063 699
rect 1109 705 1819 751
rect 1865 705 1876 751
rect 1109 642 1155 705
rect 1661 648 1707 659
rect 59 596 555 642
rect 665 596 1155 642
rect 1232 602 1243 648
rect 1289 602 1591 648
rect 30 516 194 542
rect 30 470 137 516
rect 183 470 194 516
rect 30 466 194 470
rect 254 516 418 542
rect 254 470 361 516
rect 407 470 418 516
rect 254 466 418 470
rect 509 516 555 596
rect 509 420 555 470
rect 702 516 866 542
rect 702 470 753 516
rect 799 470 866 516
rect 702 466 866 470
rect 921 516 967 527
rect 921 420 967 470
rect 1262 516 1426 542
rect 1262 470 1321 516
rect 1367 470 1426 516
rect 1262 466 1426 470
rect 1545 516 1591 602
rect 1661 516 1707 602
rect 2023 619 2069 699
rect 2227 839 2273 850
rect 2431 839 2477 918
rect 2431 782 2477 793
rect 2635 839 2681 850
rect 2273 699 2635 734
rect 2227 688 2681 699
rect 2791 839 2837 918
rect 2791 688 2837 699
rect 2995 839 3041 850
rect 2023 573 2862 619
rect 1661 478 1907 516
rect 1545 420 1591 470
rect 49 374 967 420
rect 1233 374 1591 420
rect 1681 470 1907 478
rect 1953 470 1964 516
rect 49 246 95 374
rect 1233 299 1279 374
rect 49 189 95 200
rect 273 246 319 257
rect 273 90 319 200
rect 665 246 711 257
rect 1233 242 1279 253
rect 1325 282 1635 328
rect 665 198 711 200
rect 665 196 1219 198
rect 1325 196 1371 282
rect 665 152 1371 196
rect 1205 150 1371 152
rect 1457 225 1503 236
rect 1090 95 1136 106
rect 0 49 1090 90
rect 1457 90 1503 179
rect 1589 182 1635 282
rect 1681 285 1727 470
rect 1681 228 1727 239
rect 1825 244 1871 255
rect 1825 182 1871 198
rect 2023 246 2095 573
rect 2794 564 2862 573
rect 2165 516 2211 527
rect 2165 380 2211 470
rect 2353 516 2399 527
rect 2794 518 2805 564
rect 2851 518 2862 564
rect 2995 487 3041 699
rect 2933 472 3041 487
rect 2399 470 3041 472
rect 2353 441 3041 470
rect 3199 839 3594 850
rect 3245 804 3594 839
rect 2353 426 2967 441
rect 2165 334 2875 380
rect 2023 200 2049 246
rect 2023 189 2095 200
rect 2653 277 2699 288
rect 1589 136 1871 182
rect 2653 90 2699 231
rect 2829 185 2875 334
rect 2921 288 2967 426
rect 2921 231 2967 242
rect 3013 380 3059 391
rect 3013 185 3059 334
rect 3199 288 3245 699
rect 3416 745 3482 756
rect 3416 699 3436 745
rect 3134 242 3145 288
rect 3191 242 3245 288
rect 3320 619 3366 630
rect 3320 185 3366 573
rect 3416 288 3482 699
rect 3548 736 3594 804
rect 3640 839 3686 918
rect 3640 782 3686 793
rect 3732 802 3982 848
rect 3732 736 3778 802
rect 3548 690 3778 736
rect 3844 745 3890 756
rect 3844 634 3890 699
rect 3552 588 3890 634
rect 3552 516 3598 588
rect 3552 459 3598 470
rect 3726 516 3778 542
rect 3726 470 3728 516
rect 3774 470 3778 516
rect 3726 354 3778 470
rect 3844 413 3890 588
rect 3936 516 3982 802
rect 4048 839 4094 918
rect 4048 688 4094 699
rect 4174 839 4266 850
rect 4174 699 4220 839
rect 3936 459 3982 470
rect 4080 516 4126 527
rect 4080 413 4126 470
rect 3844 367 4126 413
rect 3462 242 3482 288
rect 3416 231 3482 242
rect 3640 244 3686 255
rect 2829 139 3366 185
rect 3640 90 3686 198
rect 4048 246 4126 367
rect 4094 200 4126 246
rect 4048 189 4126 200
rect 4174 320 4266 699
rect 4424 839 4470 918
rect 4424 688 4470 699
rect 4174 180 4210 320
rect 4256 180 4266 320
rect 4174 169 4266 180
rect 4434 320 4480 331
rect 4434 90 4480 180
rect 1136 49 4592 90
rect 0 -90 4592 49
<< labels >>
flabel metal1 s 1262 466 1426 542 0 FreeSans 200 0 0 0 CLK
port 5 nsew clock input
flabel metal1 s 702 466 866 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4174 169 4266 850 0 FreeSans 200 0 0 0 Q
port 6 nsew default output
flabel metal1 s 3726 354 3778 542 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 30 466 194 542 0 FreeSans 200 0 0 0 SE
port 3 nsew default input
flabel metal1 s 254 466 418 542 0 FreeSans 200 0 0 0 SI
port 4 nsew default input
flabel metal1 s 0 918 4592 1098 0 FreeSans 200 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 4434 288 4480 331 0 FreeSans 200 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 8 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 9 nsew ground bidirectional
rlabel metal1 s 4424 806 4470 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4048 806 4094 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3640 806 3686 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2791 806 2837 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2431 806 2477 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1436 806 1504 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1017 806 1063 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 263 806 309 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4424 782 4470 806 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4048 782 4094 806 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3640 782 3686 806 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2791 782 2837 806 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2431 782 2477 806 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1017 782 1063 806 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 263 782 309 806 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4424 688 4470 782 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4048 688 4094 782 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2791 688 2837 782 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1017 688 1063 782 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 263 688 309 782 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4434 257 4480 288 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2653 257 2699 288 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4434 255 4480 257 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2653 255 2699 257 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 255 319 257 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4434 236 4480 255 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 3640 236 3686 255 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2653 236 2699 255 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 236 319 255 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4434 106 4480 236 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 3640 106 3686 236 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2653 106 2699 236 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1457 106 1503 236 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 106 319 236 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4434 90 4480 106 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 3640 90 3686 106 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2653 90 2699 106 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1457 90 1503 106 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1090 90 1136 106 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 106 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4592 90 1 VSS
port 10 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4592 1008
string GDS_END 344184
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 333480
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
