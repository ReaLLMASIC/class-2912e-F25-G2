magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 453 1654 1094
<< pwell >>
rect -86 -86 1654 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
rect 1244 69 1364 333
<< mvpmos >>
rect 144 573 244 939
rect 358 573 458 939
rect 582 573 682 939
rect 806 573 906 939
rect 1030 573 1130 939
rect 1244 573 1344 939
<< mvndiff >>
rect 36 294 124 333
rect 36 154 49 294
rect 95 154 124 294
rect 36 69 124 154
rect 244 294 348 333
rect 244 154 273 294
rect 319 154 348 294
rect 244 69 348 154
rect 468 294 572 333
rect 468 154 497 294
rect 543 154 572 294
rect 468 69 572 154
rect 692 294 796 333
rect 692 154 721 294
rect 767 154 796 294
rect 692 69 796 154
rect 916 285 1020 333
rect 916 239 945 285
rect 991 239 1020 285
rect 916 69 1020 239
rect 1140 294 1244 333
rect 1140 154 1169 294
rect 1215 154 1244 294
rect 1140 69 1244 154
rect 1364 294 1452 333
rect 1364 154 1393 294
rect 1439 154 1452 294
rect 1364 69 1452 154
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 573 358 939
rect 458 573 582 939
rect 682 861 806 939
rect 682 721 731 861
rect 777 721 806 861
rect 682 573 806 721
rect 906 573 1030 939
rect 1130 573 1244 939
rect 1344 861 1432 939
rect 1344 721 1373 861
rect 1419 721 1432 861
rect 1344 573 1432 721
<< mvndiffc >>
rect 49 154 95 294
rect 273 154 319 294
rect 497 154 543 294
rect 721 154 767 294
rect 945 239 991 285
rect 1169 154 1215 294
rect 1393 154 1439 294
<< mvpdiffc >>
rect 69 721 115 861
rect 731 721 777 861
rect 1373 721 1419 861
<< polysilicon >>
rect 144 939 244 983
rect 358 939 458 983
rect 582 939 682 983
rect 806 939 906 983
rect 1030 939 1130 983
rect 1244 939 1344 983
rect 144 500 244 573
rect 144 454 157 500
rect 203 454 244 500
rect 144 377 244 454
rect 358 500 458 573
rect 358 454 371 500
rect 417 454 458 500
rect 358 377 458 454
rect 582 500 682 573
rect 582 454 595 500
rect 641 454 682 500
rect 582 377 682 454
rect 806 500 906 573
rect 806 454 819 500
rect 865 454 906 500
rect 806 377 906 454
rect 1030 500 1130 573
rect 1030 454 1043 500
rect 1089 454 1130 500
rect 1030 377 1130 454
rect 1244 500 1344 573
rect 1244 454 1257 500
rect 1303 454 1344 500
rect 1244 377 1344 454
rect 124 333 244 377
rect 348 333 468 377
rect 572 333 692 377
rect 796 333 916 377
rect 1020 333 1140 377
rect 1244 333 1364 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
<< polycontact >>
rect 157 454 203 500
rect 371 454 417 500
rect 595 454 641 500
rect 819 454 865 500
rect 1043 454 1089 500
rect 1257 454 1303 500
<< metal1 >>
rect 0 918 1568 1098
rect 69 861 115 918
rect 69 710 115 721
rect 731 861 777 872
rect 731 603 777 721
rect 1373 861 1419 918
rect 1373 710 1419 721
rect 731 557 980 603
rect 142 500 203 542
rect 142 454 157 500
rect 360 500 428 542
rect 360 454 371 500
rect 417 454 428 500
rect 584 500 652 542
rect 584 454 595 500
rect 641 454 652 500
rect 814 500 866 511
rect 814 454 819 500
rect 865 454 866 500
rect 142 443 203 454
rect 273 351 635 397
rect 814 354 866 454
rect 934 397 980 557
rect 1038 500 1090 654
rect 1038 454 1043 500
rect 1089 454 1090 500
rect 1246 500 1314 542
rect 1246 454 1257 500
rect 1303 454 1314 500
rect 1038 443 1090 454
rect 49 294 95 305
rect 49 90 95 154
rect 273 294 319 351
rect 273 143 319 154
rect 497 294 543 305
rect 497 90 543 154
rect 589 182 635 351
rect 934 351 1308 397
rect 721 294 767 305
rect 589 154 721 182
rect 934 285 991 351
rect 1262 318 1308 351
rect 934 239 945 285
rect 934 228 991 239
rect 1169 294 1215 305
rect 767 154 1169 182
rect 1262 294 1439 318
rect 1262 242 1393 294
rect 589 136 1215 154
rect 1393 143 1439 154
rect 0 -90 1568 90
<< labels >>
flabel metal1 s 814 354 866 511 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1038 443 1090 654 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 1246 454 1314 542 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 584 454 652 542 0 FreeSans 200 0 0 0 B1
port 4 nsew default input
flabel metal1 s 360 454 428 542 0 FreeSans 200 0 0 0 B2
port 5 nsew default input
flabel metal1 s 142 443 203 542 0 FreeSans 200 0 0 0 B3
port 6 nsew default input
flabel metal1 s 0 918 1568 1098 0 FreeSans 200 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 497 90 543 305 0 FreeSans 200 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 731 603 777 872 0 FreeSans 200 0 0 0 ZN
port 7 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 9 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 10 nsew ground bidirectional
rlabel metal1 s 731 557 980 603 1 ZN
port 7 nsew default output
rlabel metal1 s 934 397 980 557 1 ZN
port 7 nsew default output
rlabel metal1 s 934 351 1308 397 1 ZN
port 7 nsew default output
rlabel metal1 s 1262 318 1308 351 1 ZN
port 7 nsew default output
rlabel metal1 s 934 318 991 351 1 ZN
port 7 nsew default output
rlabel metal1 s 1262 242 1439 318 1 ZN
port 7 nsew default output
rlabel metal1 s 934 242 991 318 1 ZN
port 7 nsew default output
rlabel metal1 s 1393 228 1439 242 1 ZN
port 7 nsew default output
rlabel metal1 s 934 228 991 242 1 ZN
port 7 nsew default output
rlabel metal1 s 1393 143 1439 228 1 ZN
port 7 nsew default output
rlabel metal1 s 1373 710 1419 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 69 710 115 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 90 95 305 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1568 90 1 VSS
port 11 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1568 1008
string GDS_END 186680
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 181964
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
