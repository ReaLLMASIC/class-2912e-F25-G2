magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -51 24849 13013 25405
rect -51 505 505 24849
rect 12457 505 13013 24849
rect -51 -51 13013 505
<< mvnmos >>
rect 1481 23733 11481 23873
rect 1481 23489 11481 23629
rect 1481 23245 11481 23385
rect 1481 23001 11481 23141
rect 1481 22757 11481 22897
rect 1481 22513 11481 22653
rect 1481 22269 11481 22409
rect 1481 22025 11481 22165
rect 1481 21781 11481 21921
rect 1481 21537 11481 21677
rect 1481 21293 11481 21433
rect 1481 21049 11481 21189
rect 1481 20805 11481 20945
rect 1481 20561 11481 20701
rect 1481 20317 11481 20457
rect 1481 20073 11481 20213
rect 1481 19829 11481 19969
rect 1481 19585 11481 19725
rect 1481 19341 11481 19481
rect 1481 19097 11481 19237
rect 1481 17861 11481 18001
rect 1481 17617 11481 17757
rect 1481 17373 11481 17513
rect 1481 17129 11481 17269
rect 1481 16885 11481 17025
rect 1481 16641 11481 16781
rect 1481 16397 11481 16537
rect 1481 16153 11481 16293
rect 1481 15909 11481 16049
rect 1481 15665 11481 15805
rect 1481 15421 11481 15561
rect 1481 15177 11481 15317
rect 1481 14933 11481 15073
rect 1481 14689 11481 14829
rect 1481 14445 11481 14585
rect 1481 14201 11481 14341
rect 1481 13957 11481 14097
rect 1481 13713 11481 13853
rect 1481 13469 11481 13609
rect 1481 13225 11481 13365
rect 1481 11989 11481 12129
rect 1481 11745 11481 11885
rect 1481 11501 11481 11641
rect 1481 11257 11481 11397
rect 1481 11013 11481 11153
rect 1481 10769 11481 10909
rect 1481 10525 11481 10665
rect 1481 10281 11481 10421
rect 1481 10037 11481 10177
rect 1481 9793 11481 9933
rect 1481 9549 11481 9689
rect 1481 9305 11481 9445
rect 1481 9061 11481 9201
rect 1481 8817 11481 8957
rect 1481 8573 11481 8713
rect 1481 8329 11481 8469
rect 1481 8085 11481 8225
rect 1481 7841 11481 7981
rect 1481 7597 11481 7737
rect 1481 7353 11481 7493
rect 1481 6117 11481 6257
rect 1481 5873 11481 6013
rect 1481 5629 11481 5769
rect 1481 5385 11481 5525
rect 1481 5141 11481 5281
rect 1481 4897 11481 5037
rect 1481 4653 11481 4793
rect 1481 4409 11481 4549
rect 1481 4165 11481 4305
rect 1481 3921 11481 4061
rect 1481 3677 11481 3817
rect 1481 3433 11481 3573
rect 1481 3189 11481 3329
rect 1481 2945 11481 3085
rect 1481 2701 11481 2841
rect 1481 2457 11481 2597
rect 1481 2213 11481 2353
rect 1481 1969 11481 2109
rect 1481 1725 11481 1865
rect 1481 1481 11481 1621
<< mvndiff >>
rect 1481 23948 11481 23961
rect 1481 23902 1494 23948
rect 11468 23902 11481 23948
rect 1481 23873 11481 23902
rect 1481 23704 11481 23733
rect 1481 23658 1494 23704
rect 11468 23658 11481 23704
rect 1481 23629 11481 23658
rect 1481 23460 11481 23489
rect 1481 23414 1494 23460
rect 11468 23414 11481 23460
rect 1481 23385 11481 23414
rect 1481 23216 11481 23245
rect 1481 23170 1494 23216
rect 11468 23170 11481 23216
rect 1481 23141 11481 23170
rect 1481 22972 11481 23001
rect 1481 22926 1494 22972
rect 11468 22926 11481 22972
rect 1481 22897 11481 22926
rect 1481 22728 11481 22757
rect 1481 22682 1494 22728
rect 11468 22682 11481 22728
rect 1481 22653 11481 22682
rect 1481 22484 11481 22513
rect 1481 22438 1494 22484
rect 11468 22438 11481 22484
rect 1481 22409 11481 22438
rect 1481 22240 11481 22269
rect 1481 22194 1494 22240
rect 11468 22194 11481 22240
rect 1481 22165 11481 22194
rect 1481 21996 11481 22025
rect 1481 21950 1494 21996
rect 11468 21950 11481 21996
rect 1481 21921 11481 21950
rect 1481 21752 11481 21781
rect 1481 21706 1494 21752
rect 11468 21706 11481 21752
rect 1481 21677 11481 21706
rect 1481 21508 11481 21537
rect 1481 21462 1494 21508
rect 11468 21462 11481 21508
rect 1481 21433 11481 21462
rect 1481 21264 11481 21293
rect 1481 21218 1494 21264
rect 11468 21218 11481 21264
rect 1481 21189 11481 21218
rect 1481 21020 11481 21049
rect 1481 20974 1494 21020
rect 11468 20974 11481 21020
rect 1481 20945 11481 20974
rect 1481 20776 11481 20805
rect 1481 20730 1494 20776
rect 11468 20730 11481 20776
rect 1481 20701 11481 20730
rect 1481 20532 11481 20561
rect 1481 20486 1494 20532
rect 11468 20486 11481 20532
rect 1481 20457 11481 20486
rect 1481 20288 11481 20317
rect 1481 20242 1494 20288
rect 11468 20242 11481 20288
rect 1481 20213 11481 20242
rect 1481 20044 11481 20073
rect 1481 19998 1494 20044
rect 11468 19998 11481 20044
rect 1481 19969 11481 19998
rect 1481 19800 11481 19829
rect 1481 19754 1494 19800
rect 11468 19754 11481 19800
rect 1481 19725 11481 19754
rect 1481 19556 11481 19585
rect 1481 19510 1494 19556
rect 11468 19510 11481 19556
rect 1481 19481 11481 19510
rect 1481 19312 11481 19341
rect 1481 19266 1494 19312
rect 11468 19266 11481 19312
rect 1481 19237 11481 19266
rect 1481 19068 11481 19097
rect 1481 19022 1494 19068
rect 11468 19022 11481 19068
rect 1481 19009 11481 19022
rect 1481 18076 11481 18089
rect 1481 18030 1494 18076
rect 11468 18030 11481 18076
rect 1481 18001 11481 18030
rect 1481 17832 11481 17861
rect 1481 17786 1494 17832
rect 11468 17786 11481 17832
rect 1481 17757 11481 17786
rect 1481 17588 11481 17617
rect 1481 17542 1494 17588
rect 11468 17542 11481 17588
rect 1481 17513 11481 17542
rect 1481 17344 11481 17373
rect 1481 17298 1494 17344
rect 11468 17298 11481 17344
rect 1481 17269 11481 17298
rect 1481 17100 11481 17129
rect 1481 17054 1494 17100
rect 11468 17054 11481 17100
rect 1481 17025 11481 17054
rect 1481 16856 11481 16885
rect 1481 16810 1494 16856
rect 11468 16810 11481 16856
rect 1481 16781 11481 16810
rect 1481 16612 11481 16641
rect 1481 16566 1494 16612
rect 11468 16566 11481 16612
rect 1481 16537 11481 16566
rect 1481 16368 11481 16397
rect 1481 16322 1494 16368
rect 11468 16322 11481 16368
rect 1481 16293 11481 16322
rect 1481 16124 11481 16153
rect 1481 16078 1494 16124
rect 11468 16078 11481 16124
rect 1481 16049 11481 16078
rect 1481 15880 11481 15909
rect 1481 15834 1494 15880
rect 11468 15834 11481 15880
rect 1481 15805 11481 15834
rect 1481 15636 11481 15665
rect 1481 15590 1494 15636
rect 11468 15590 11481 15636
rect 1481 15561 11481 15590
rect 1481 15392 11481 15421
rect 1481 15346 1494 15392
rect 11468 15346 11481 15392
rect 1481 15317 11481 15346
rect 1481 15148 11481 15177
rect 1481 15102 1494 15148
rect 11468 15102 11481 15148
rect 1481 15073 11481 15102
rect 1481 14904 11481 14933
rect 1481 14858 1494 14904
rect 11468 14858 11481 14904
rect 1481 14829 11481 14858
rect 1481 14660 11481 14689
rect 1481 14614 1494 14660
rect 11468 14614 11481 14660
rect 1481 14585 11481 14614
rect 1481 14416 11481 14445
rect 1481 14370 1494 14416
rect 11468 14370 11481 14416
rect 1481 14341 11481 14370
rect 1481 14172 11481 14201
rect 1481 14126 1494 14172
rect 11468 14126 11481 14172
rect 1481 14097 11481 14126
rect 1481 13928 11481 13957
rect 1481 13882 1494 13928
rect 11468 13882 11481 13928
rect 1481 13853 11481 13882
rect 1481 13684 11481 13713
rect 1481 13638 1494 13684
rect 11468 13638 11481 13684
rect 1481 13609 11481 13638
rect 1481 13440 11481 13469
rect 1481 13394 1494 13440
rect 11468 13394 11481 13440
rect 1481 13365 11481 13394
rect 1481 13196 11481 13225
rect 1481 13150 1494 13196
rect 11468 13150 11481 13196
rect 1481 13137 11481 13150
rect 1481 12204 11481 12217
rect 1481 12158 1494 12204
rect 11468 12158 11481 12204
rect 1481 12129 11481 12158
rect 1481 11960 11481 11989
rect 1481 11914 1494 11960
rect 11468 11914 11481 11960
rect 1481 11885 11481 11914
rect 1481 11716 11481 11745
rect 1481 11670 1494 11716
rect 11468 11670 11481 11716
rect 1481 11641 11481 11670
rect 1481 11472 11481 11501
rect 1481 11426 1494 11472
rect 11468 11426 11481 11472
rect 1481 11397 11481 11426
rect 1481 11228 11481 11257
rect 1481 11182 1494 11228
rect 11468 11182 11481 11228
rect 1481 11153 11481 11182
rect 1481 10984 11481 11013
rect 1481 10938 1494 10984
rect 11468 10938 11481 10984
rect 1481 10909 11481 10938
rect 1481 10740 11481 10769
rect 1481 10694 1494 10740
rect 11468 10694 11481 10740
rect 1481 10665 11481 10694
rect 1481 10496 11481 10525
rect 1481 10450 1494 10496
rect 11468 10450 11481 10496
rect 1481 10421 11481 10450
rect 1481 10252 11481 10281
rect 1481 10206 1494 10252
rect 11468 10206 11481 10252
rect 1481 10177 11481 10206
rect 1481 10008 11481 10037
rect 1481 9962 1494 10008
rect 11468 9962 11481 10008
rect 1481 9933 11481 9962
rect 1481 9764 11481 9793
rect 1481 9718 1494 9764
rect 11468 9718 11481 9764
rect 1481 9689 11481 9718
rect 1481 9520 11481 9549
rect 1481 9474 1494 9520
rect 11468 9474 11481 9520
rect 1481 9445 11481 9474
rect 1481 9276 11481 9305
rect 1481 9230 1494 9276
rect 11468 9230 11481 9276
rect 1481 9201 11481 9230
rect 1481 9032 11481 9061
rect 1481 8986 1494 9032
rect 11468 8986 11481 9032
rect 1481 8957 11481 8986
rect 1481 8788 11481 8817
rect 1481 8742 1494 8788
rect 11468 8742 11481 8788
rect 1481 8713 11481 8742
rect 1481 8544 11481 8573
rect 1481 8498 1494 8544
rect 11468 8498 11481 8544
rect 1481 8469 11481 8498
rect 1481 8300 11481 8329
rect 1481 8254 1494 8300
rect 11468 8254 11481 8300
rect 1481 8225 11481 8254
rect 1481 8056 11481 8085
rect 1481 8010 1494 8056
rect 11468 8010 11481 8056
rect 1481 7981 11481 8010
rect 1481 7812 11481 7841
rect 1481 7766 1494 7812
rect 11468 7766 11481 7812
rect 1481 7737 11481 7766
rect 1481 7568 11481 7597
rect 1481 7522 1494 7568
rect 11468 7522 11481 7568
rect 1481 7493 11481 7522
rect 1481 7324 11481 7353
rect 1481 7278 1494 7324
rect 11468 7278 11481 7324
rect 1481 7265 11481 7278
rect 1481 6332 11481 6345
rect 1481 6286 1494 6332
rect 11468 6286 11481 6332
rect 1481 6257 11481 6286
rect 1481 6088 11481 6117
rect 1481 6042 1494 6088
rect 11468 6042 11481 6088
rect 1481 6013 11481 6042
rect 1481 5844 11481 5873
rect 1481 5798 1494 5844
rect 11468 5798 11481 5844
rect 1481 5769 11481 5798
rect 1481 5600 11481 5629
rect 1481 5554 1494 5600
rect 11468 5554 11481 5600
rect 1481 5525 11481 5554
rect 1481 5356 11481 5385
rect 1481 5310 1494 5356
rect 11468 5310 11481 5356
rect 1481 5281 11481 5310
rect 1481 5112 11481 5141
rect 1481 5066 1494 5112
rect 11468 5066 11481 5112
rect 1481 5037 11481 5066
rect 1481 4868 11481 4897
rect 1481 4822 1494 4868
rect 11468 4822 11481 4868
rect 1481 4793 11481 4822
rect 1481 4624 11481 4653
rect 1481 4578 1494 4624
rect 11468 4578 11481 4624
rect 1481 4549 11481 4578
rect 1481 4380 11481 4409
rect 1481 4334 1494 4380
rect 11468 4334 11481 4380
rect 1481 4305 11481 4334
rect 1481 4136 11481 4165
rect 1481 4090 1494 4136
rect 11468 4090 11481 4136
rect 1481 4061 11481 4090
rect 1481 3892 11481 3921
rect 1481 3846 1494 3892
rect 11468 3846 11481 3892
rect 1481 3817 11481 3846
rect 1481 3648 11481 3677
rect 1481 3602 1494 3648
rect 11468 3602 11481 3648
rect 1481 3573 11481 3602
rect 1481 3404 11481 3433
rect 1481 3358 1494 3404
rect 11468 3358 11481 3404
rect 1481 3329 11481 3358
rect 1481 3160 11481 3189
rect 1481 3114 1494 3160
rect 11468 3114 11481 3160
rect 1481 3085 11481 3114
rect 1481 2916 11481 2945
rect 1481 2870 1494 2916
rect 11468 2870 11481 2916
rect 1481 2841 11481 2870
rect 1481 2672 11481 2701
rect 1481 2626 1494 2672
rect 11468 2626 11481 2672
rect 1481 2597 11481 2626
rect 1481 2428 11481 2457
rect 1481 2382 1494 2428
rect 11468 2382 11481 2428
rect 1481 2353 11481 2382
rect 1481 2184 11481 2213
rect 1481 2138 1494 2184
rect 11468 2138 11481 2184
rect 1481 2109 11481 2138
rect 1481 1940 11481 1969
rect 1481 1894 1494 1940
rect 11468 1894 11481 1940
rect 1481 1865 11481 1894
rect 1481 1696 11481 1725
rect 1481 1650 1494 1696
rect 11468 1650 11481 1696
rect 1481 1621 11481 1650
rect 1481 1452 11481 1481
rect 1481 1406 1494 1452
rect 11468 1406 11481 1452
rect 1481 1393 11481 1406
<< mvndiffc >>
rect 1494 23902 11468 23948
rect 1494 23658 11468 23704
rect 1494 23414 11468 23460
rect 1494 23170 11468 23216
rect 1494 22926 11468 22972
rect 1494 22682 11468 22728
rect 1494 22438 11468 22484
rect 1494 22194 11468 22240
rect 1494 21950 11468 21996
rect 1494 21706 11468 21752
rect 1494 21462 11468 21508
rect 1494 21218 11468 21264
rect 1494 20974 11468 21020
rect 1494 20730 11468 20776
rect 1494 20486 11468 20532
rect 1494 20242 11468 20288
rect 1494 19998 11468 20044
rect 1494 19754 11468 19800
rect 1494 19510 11468 19556
rect 1494 19266 11468 19312
rect 1494 19022 11468 19068
rect 1494 18030 11468 18076
rect 1494 17786 11468 17832
rect 1494 17542 11468 17588
rect 1494 17298 11468 17344
rect 1494 17054 11468 17100
rect 1494 16810 11468 16856
rect 1494 16566 11468 16612
rect 1494 16322 11468 16368
rect 1494 16078 11468 16124
rect 1494 15834 11468 15880
rect 1494 15590 11468 15636
rect 1494 15346 11468 15392
rect 1494 15102 11468 15148
rect 1494 14858 11468 14904
rect 1494 14614 11468 14660
rect 1494 14370 11468 14416
rect 1494 14126 11468 14172
rect 1494 13882 11468 13928
rect 1494 13638 11468 13684
rect 1494 13394 11468 13440
rect 1494 13150 11468 13196
rect 1494 12158 11468 12204
rect 1494 11914 11468 11960
rect 1494 11670 11468 11716
rect 1494 11426 11468 11472
rect 1494 11182 11468 11228
rect 1494 10938 11468 10984
rect 1494 10694 11468 10740
rect 1494 10450 11468 10496
rect 1494 10206 11468 10252
rect 1494 9962 11468 10008
rect 1494 9718 11468 9764
rect 1494 9474 11468 9520
rect 1494 9230 11468 9276
rect 1494 8986 11468 9032
rect 1494 8742 11468 8788
rect 1494 8498 11468 8544
rect 1494 8254 11468 8300
rect 1494 8010 11468 8056
rect 1494 7766 11468 7812
rect 1494 7522 11468 7568
rect 1494 7278 11468 7324
rect 1494 6286 11468 6332
rect 1494 6042 11468 6088
rect 1494 5798 11468 5844
rect 1494 5554 11468 5600
rect 1494 5310 11468 5356
rect 1494 5066 11468 5112
rect 1494 4822 11468 4868
rect 1494 4578 11468 4624
rect 1494 4334 11468 4380
rect 1494 4090 11468 4136
rect 1494 3846 11468 3892
rect 1494 3602 11468 3648
rect 1494 3358 11468 3404
rect 1494 3114 11468 3160
rect 1494 2870 11468 2916
rect 1494 2626 11468 2672
rect 1494 2382 11468 2428
rect 1494 2138 11468 2184
rect 1494 1894 11468 1940
rect 1494 1650 11468 1696
rect 1494 1406 11468 1452
<< psubdiff >>
rect 582 24700 12380 24722
rect 582 654 604 24700
rect 950 24354 1058 24700
rect 11904 24354 12012 24700
rect 950 24332 12012 24354
rect 950 18644 972 24332
rect 11990 18644 12012 24332
rect 950 18622 12012 18644
rect 950 18476 1058 18622
rect 11904 18476 12012 18622
rect 950 18454 12012 18476
rect 950 12772 972 18454
rect 11990 12772 12012 18454
rect 950 12750 12012 12772
rect 950 12604 1058 12750
rect 11904 12604 12012 12750
rect 950 12582 12012 12604
rect 950 6900 972 12582
rect 11990 6900 12012 12582
rect 950 6878 12012 6900
rect 950 6732 1058 6878
rect 11904 6732 12012 6878
rect 950 6710 12012 6732
rect 950 1022 972 6710
rect 11990 1022 12012 6710
rect 950 1000 12012 1022
rect 950 654 1058 1000
rect 11904 654 12012 1000
rect 12358 654 12380 24700
rect 582 632 12380 654
<< nsubdiff >>
rect 32 25300 12930 25322
rect 32 54 54 25300
rect 400 24954 508 25300
rect 12454 24954 12562 25300
rect 400 24932 12562 24954
rect 400 422 422 24932
rect 12540 422 12562 24932
rect 400 400 12562 422
rect 400 54 508 400
rect 12454 54 12562 400
rect 12908 54 12930 25300
rect 32 32 12930 54
<< psubdiffcont >>
rect 604 654 950 24700
rect 1058 24354 11904 24700
rect 1058 18476 11904 18622
rect 1058 12604 11904 12750
rect 1058 6732 11904 6878
rect 1058 654 11904 1000
rect 12012 654 12358 24700
<< nsubdiffcont >>
rect 54 54 400 25300
rect 508 24954 12454 25300
rect 508 54 12454 400
rect 12562 54 12908 25300
<< polysilicon >>
rect 1237 23808 1481 23873
rect 1237 19162 1256 23808
rect 1402 23733 1481 23808
rect 11481 23808 11725 23873
rect 11481 23733 11560 23808
rect 1402 23629 1421 23733
rect 11541 23629 11560 23733
rect 1402 23489 1481 23629
rect 11481 23489 11560 23629
rect 1402 23385 1421 23489
rect 11541 23385 11560 23489
rect 1402 23245 1481 23385
rect 11481 23245 11560 23385
rect 1402 23141 1421 23245
rect 11541 23141 11560 23245
rect 1402 23001 1481 23141
rect 11481 23001 11560 23141
rect 1402 22897 1421 23001
rect 11541 22897 11560 23001
rect 1402 22757 1481 22897
rect 11481 22757 11560 22897
rect 1402 22653 1421 22757
rect 11541 22653 11560 22757
rect 1402 22513 1481 22653
rect 11481 22513 11560 22653
rect 1402 22409 1421 22513
rect 11541 22409 11560 22513
rect 1402 22269 1481 22409
rect 11481 22269 11560 22409
rect 1402 22165 1421 22269
rect 11541 22165 11560 22269
rect 1402 22025 1481 22165
rect 11481 22025 11560 22165
rect 1402 21921 1421 22025
rect 11541 21921 11560 22025
rect 1402 21781 1481 21921
rect 11481 21781 11560 21921
rect 1402 21677 1421 21781
rect 11541 21677 11560 21781
rect 1402 21537 1481 21677
rect 11481 21537 11560 21677
rect 1402 21433 1421 21537
rect 11541 21433 11560 21537
rect 1402 21293 1481 21433
rect 11481 21293 11560 21433
rect 1402 21189 1421 21293
rect 11541 21189 11560 21293
rect 1402 21049 1481 21189
rect 11481 21049 11560 21189
rect 1402 20945 1421 21049
rect 11541 20945 11560 21049
rect 1402 20805 1481 20945
rect 11481 20805 11560 20945
rect 1402 20701 1421 20805
rect 11541 20701 11560 20805
rect 1402 20561 1481 20701
rect 11481 20561 11560 20701
rect 1402 20457 1421 20561
rect 11541 20457 11560 20561
rect 1402 20317 1481 20457
rect 11481 20317 11560 20457
rect 1402 20213 1421 20317
rect 11541 20213 11560 20317
rect 1402 20073 1481 20213
rect 11481 20073 11560 20213
rect 1402 19969 1421 20073
rect 11541 19969 11560 20073
rect 1402 19829 1481 19969
rect 11481 19829 11560 19969
rect 1402 19725 1421 19829
rect 11541 19725 11560 19829
rect 1402 19585 1481 19725
rect 11481 19585 11560 19725
rect 1402 19481 1421 19585
rect 11541 19481 11560 19585
rect 1402 19341 1481 19481
rect 11481 19341 11560 19481
rect 1402 19237 1421 19341
rect 11541 19237 11560 19341
rect 1402 19162 1481 19237
rect 1237 19097 1481 19162
rect 11481 19162 11560 19237
rect 11706 19162 11725 23808
rect 11481 19097 11725 19162
rect 1237 17936 1481 18001
rect 1237 13290 1256 17936
rect 1402 17861 1481 17936
rect 11481 17936 11725 18001
rect 11481 17861 11560 17936
rect 1402 17757 1421 17861
rect 11541 17757 11560 17861
rect 1402 17617 1481 17757
rect 11481 17617 11560 17757
rect 1402 17513 1421 17617
rect 11541 17513 11560 17617
rect 1402 17373 1481 17513
rect 11481 17373 11560 17513
rect 1402 17269 1421 17373
rect 11541 17269 11560 17373
rect 1402 17129 1481 17269
rect 11481 17129 11560 17269
rect 1402 17025 1421 17129
rect 11541 17025 11560 17129
rect 1402 16885 1481 17025
rect 11481 16885 11560 17025
rect 1402 16781 1421 16885
rect 11541 16781 11560 16885
rect 1402 16641 1481 16781
rect 11481 16641 11560 16781
rect 1402 16537 1421 16641
rect 11541 16537 11560 16641
rect 1402 16397 1481 16537
rect 11481 16397 11560 16537
rect 1402 16293 1421 16397
rect 11541 16293 11560 16397
rect 1402 16153 1481 16293
rect 11481 16153 11560 16293
rect 1402 16049 1421 16153
rect 11541 16049 11560 16153
rect 1402 15909 1481 16049
rect 11481 15909 11560 16049
rect 1402 15805 1421 15909
rect 11541 15805 11560 15909
rect 1402 15665 1481 15805
rect 11481 15665 11560 15805
rect 1402 15561 1421 15665
rect 11541 15561 11560 15665
rect 1402 15421 1481 15561
rect 11481 15421 11560 15561
rect 1402 15317 1421 15421
rect 11541 15317 11560 15421
rect 1402 15177 1481 15317
rect 11481 15177 11560 15317
rect 1402 15073 1421 15177
rect 11541 15073 11560 15177
rect 1402 14933 1481 15073
rect 11481 14933 11560 15073
rect 1402 14829 1421 14933
rect 11541 14829 11560 14933
rect 1402 14689 1481 14829
rect 11481 14689 11560 14829
rect 1402 14585 1421 14689
rect 11541 14585 11560 14689
rect 1402 14445 1481 14585
rect 11481 14445 11560 14585
rect 1402 14341 1421 14445
rect 11541 14341 11560 14445
rect 1402 14201 1481 14341
rect 11481 14201 11560 14341
rect 1402 14097 1421 14201
rect 11541 14097 11560 14201
rect 1402 13957 1481 14097
rect 11481 13957 11560 14097
rect 1402 13853 1421 13957
rect 11541 13853 11560 13957
rect 1402 13713 1481 13853
rect 11481 13713 11560 13853
rect 1402 13609 1421 13713
rect 11541 13609 11560 13713
rect 1402 13469 1481 13609
rect 11481 13469 11560 13609
rect 1402 13365 1421 13469
rect 11541 13365 11560 13469
rect 1402 13290 1481 13365
rect 1237 13225 1481 13290
rect 11481 13290 11560 13365
rect 11706 13290 11725 17936
rect 11481 13225 11725 13290
rect 1237 12064 1481 12129
rect 1237 7418 1256 12064
rect 1402 11989 1481 12064
rect 11481 12064 11725 12129
rect 11481 11989 11560 12064
rect 1402 11885 1421 11989
rect 11541 11885 11560 11989
rect 1402 11745 1481 11885
rect 11481 11745 11560 11885
rect 1402 11641 1421 11745
rect 11541 11641 11560 11745
rect 1402 11501 1481 11641
rect 11481 11501 11560 11641
rect 1402 11397 1421 11501
rect 11541 11397 11560 11501
rect 1402 11257 1481 11397
rect 11481 11257 11560 11397
rect 1402 11153 1421 11257
rect 11541 11153 11560 11257
rect 1402 11013 1481 11153
rect 11481 11013 11560 11153
rect 1402 10909 1421 11013
rect 11541 10909 11560 11013
rect 1402 10769 1481 10909
rect 11481 10769 11560 10909
rect 1402 10665 1421 10769
rect 11541 10665 11560 10769
rect 1402 10525 1481 10665
rect 11481 10525 11560 10665
rect 1402 10421 1421 10525
rect 11541 10421 11560 10525
rect 1402 10281 1481 10421
rect 11481 10281 11560 10421
rect 1402 10177 1421 10281
rect 11541 10177 11560 10281
rect 1402 10037 1481 10177
rect 11481 10037 11560 10177
rect 1402 9933 1421 10037
rect 11541 9933 11560 10037
rect 1402 9793 1481 9933
rect 11481 9793 11560 9933
rect 1402 9689 1421 9793
rect 11541 9689 11560 9793
rect 1402 9549 1481 9689
rect 11481 9549 11560 9689
rect 1402 9445 1421 9549
rect 11541 9445 11560 9549
rect 1402 9305 1481 9445
rect 11481 9305 11560 9445
rect 1402 9201 1421 9305
rect 11541 9201 11560 9305
rect 1402 9061 1481 9201
rect 11481 9061 11560 9201
rect 1402 8957 1421 9061
rect 11541 8957 11560 9061
rect 1402 8817 1481 8957
rect 11481 8817 11560 8957
rect 1402 8713 1421 8817
rect 11541 8713 11560 8817
rect 1402 8573 1481 8713
rect 11481 8573 11560 8713
rect 1402 8469 1421 8573
rect 11541 8469 11560 8573
rect 1402 8329 1481 8469
rect 11481 8329 11560 8469
rect 1402 8225 1421 8329
rect 11541 8225 11560 8329
rect 1402 8085 1481 8225
rect 11481 8085 11560 8225
rect 1402 7981 1421 8085
rect 11541 7981 11560 8085
rect 1402 7841 1481 7981
rect 11481 7841 11560 7981
rect 1402 7737 1421 7841
rect 11541 7737 11560 7841
rect 1402 7597 1481 7737
rect 11481 7597 11560 7737
rect 1402 7493 1421 7597
rect 11541 7493 11560 7597
rect 1402 7418 1481 7493
rect 1237 7353 1481 7418
rect 11481 7418 11560 7493
rect 11706 7418 11725 12064
rect 11481 7353 11725 7418
rect 1237 6192 1481 6257
rect 1237 1546 1256 6192
rect 1402 6117 1481 6192
rect 11481 6192 11725 6257
rect 11481 6117 11560 6192
rect 1402 6013 1421 6117
rect 11541 6013 11560 6117
rect 1402 5873 1481 6013
rect 11481 5873 11560 6013
rect 1402 5769 1421 5873
rect 11541 5769 11560 5873
rect 1402 5629 1481 5769
rect 11481 5629 11560 5769
rect 1402 5525 1421 5629
rect 11541 5525 11560 5629
rect 1402 5385 1481 5525
rect 11481 5385 11560 5525
rect 1402 5281 1421 5385
rect 11541 5281 11560 5385
rect 1402 5141 1481 5281
rect 11481 5141 11560 5281
rect 1402 5037 1421 5141
rect 11541 5037 11560 5141
rect 1402 4897 1481 5037
rect 11481 4897 11560 5037
rect 1402 4793 1421 4897
rect 11541 4793 11560 4897
rect 1402 4653 1481 4793
rect 11481 4653 11560 4793
rect 1402 4549 1421 4653
rect 11541 4549 11560 4653
rect 1402 4409 1481 4549
rect 11481 4409 11560 4549
rect 1402 4305 1421 4409
rect 11541 4305 11560 4409
rect 1402 4165 1481 4305
rect 11481 4165 11560 4305
rect 1402 4061 1421 4165
rect 11541 4061 11560 4165
rect 1402 3921 1481 4061
rect 11481 3921 11560 4061
rect 1402 3817 1421 3921
rect 11541 3817 11560 3921
rect 1402 3677 1481 3817
rect 11481 3677 11560 3817
rect 1402 3573 1421 3677
rect 11541 3573 11560 3677
rect 1402 3433 1481 3573
rect 11481 3433 11560 3573
rect 1402 3329 1421 3433
rect 11541 3329 11560 3433
rect 1402 3189 1481 3329
rect 11481 3189 11560 3329
rect 1402 3085 1421 3189
rect 11541 3085 11560 3189
rect 1402 2945 1481 3085
rect 11481 2945 11560 3085
rect 1402 2841 1421 2945
rect 11541 2841 11560 2945
rect 1402 2701 1481 2841
rect 11481 2701 11560 2841
rect 1402 2597 1421 2701
rect 11541 2597 11560 2701
rect 1402 2457 1481 2597
rect 11481 2457 11560 2597
rect 1402 2353 1421 2457
rect 11541 2353 11560 2457
rect 1402 2213 1481 2353
rect 11481 2213 11560 2353
rect 1402 2109 1421 2213
rect 11541 2109 11560 2213
rect 1402 1969 1481 2109
rect 11481 1969 11560 2109
rect 1402 1865 1421 1969
rect 11541 1865 11560 1969
rect 1402 1725 1481 1865
rect 11481 1725 11560 1865
rect 1402 1621 1421 1725
rect 11541 1621 11560 1725
rect 1402 1546 1481 1621
rect 1237 1481 1481 1546
rect 11481 1546 11560 1621
rect 11706 1546 11725 6192
rect 11481 1481 11725 1546
<< polycontact >>
rect 1256 19162 1402 23808
rect 11560 19162 11706 23808
rect 1256 13290 1402 17936
rect 11560 13290 11706 17936
rect 1256 7418 1402 12064
rect 11560 7418 11706 12064
rect 1256 1546 1402 6192
rect 11560 1546 11706 6192
<< metal1 >>
rect 43 25300 12919 25311
rect 43 54 54 25300
rect 400 24954 508 25300
rect 12454 24954 12562 25300
rect 400 24943 12562 24954
rect 400 411 411 24943
rect 593 24700 12369 24711
rect 593 654 604 24700
rect 950 24354 1058 24700
rect 11904 24354 12012 24700
rect 950 24343 12012 24354
rect 950 18641 961 24343
rect 1213 24053 11749 24253
rect 1213 23887 1413 24053
rect 1481 23951 11481 23963
rect 1481 23948 1760 23951
rect 1812 23948 1868 23951
rect 1920 23948 1976 23951
rect 2028 23948 2084 23951
rect 2136 23948 2192 23951
rect 2244 23948 2300 23951
rect 2352 23948 2408 23951
rect 2460 23948 2516 23951
rect 2568 23948 2624 23951
rect 2676 23948 2732 23951
rect 2784 23948 2840 23951
rect 2892 23948 2948 23951
rect 3000 23948 3056 23951
rect 3108 23948 3164 23951
rect 3216 23948 3272 23951
rect 3324 23948 3380 23951
rect 3432 23948 3488 23951
rect 3540 23948 3596 23951
rect 3648 23948 3704 23951
rect 3756 23948 4130 23951
rect 4182 23948 4238 23951
rect 4290 23948 4346 23951
rect 4398 23948 4454 23951
rect 4506 23948 4562 23951
rect 4614 23948 4670 23951
rect 4722 23948 4778 23951
rect 4830 23948 4886 23951
rect 4938 23948 4994 23951
rect 5046 23948 5102 23951
rect 5154 23948 5210 23951
rect 5262 23948 5318 23951
rect 5370 23948 5426 23951
rect 5478 23948 5534 23951
rect 5586 23948 5642 23951
rect 5694 23948 5750 23951
rect 5802 23948 5858 23951
rect 5910 23948 5966 23951
rect 6018 23948 6074 23951
rect 6126 23948 6836 23951
rect 6888 23948 6944 23951
rect 6996 23948 7052 23951
rect 7104 23948 7160 23951
rect 7212 23948 7268 23951
rect 7320 23948 7376 23951
rect 7428 23948 7484 23951
rect 7536 23948 7592 23951
rect 7644 23948 7700 23951
rect 7752 23948 7808 23951
rect 7860 23948 7916 23951
rect 7968 23948 8024 23951
rect 8076 23948 8132 23951
rect 8184 23948 8240 23951
rect 8292 23948 8348 23951
rect 8400 23948 8456 23951
rect 8508 23948 8564 23951
rect 8616 23948 8672 23951
rect 8724 23948 8780 23951
rect 8832 23948 9206 23951
rect 9258 23948 9314 23951
rect 9366 23948 9422 23951
rect 9474 23948 9530 23951
rect 9582 23948 9638 23951
rect 9690 23948 9746 23951
rect 9798 23948 9854 23951
rect 9906 23948 9962 23951
rect 10014 23948 10070 23951
rect 10122 23948 10178 23951
rect 10230 23948 10286 23951
rect 10338 23948 10394 23951
rect 10446 23948 10502 23951
rect 10554 23948 10610 23951
rect 10662 23948 10718 23951
rect 10770 23948 10826 23951
rect 10878 23948 10934 23951
rect 10986 23948 11042 23951
rect 11094 23948 11150 23951
rect 11202 23948 11481 23951
rect 1481 23902 1494 23948
rect 11468 23902 11481 23948
rect 1481 23899 1760 23902
rect 1812 23899 1868 23902
rect 1920 23899 1976 23902
rect 2028 23899 2084 23902
rect 2136 23899 2192 23902
rect 2244 23899 2300 23902
rect 2352 23899 2408 23902
rect 2460 23899 2516 23902
rect 2568 23899 2624 23902
rect 2676 23899 2732 23902
rect 2784 23899 2840 23902
rect 2892 23899 2948 23902
rect 3000 23899 3056 23902
rect 3108 23899 3164 23902
rect 3216 23899 3272 23902
rect 3324 23899 3380 23902
rect 3432 23899 3488 23902
rect 3540 23899 3596 23902
rect 3648 23899 3704 23902
rect 3756 23899 4130 23902
rect 4182 23899 4238 23902
rect 4290 23899 4346 23902
rect 4398 23899 4454 23902
rect 4506 23899 4562 23902
rect 4614 23899 4670 23902
rect 4722 23899 4778 23902
rect 4830 23899 4886 23902
rect 4938 23899 4994 23902
rect 5046 23899 5102 23902
rect 5154 23899 5210 23902
rect 5262 23899 5318 23902
rect 5370 23899 5426 23902
rect 5478 23899 5534 23902
rect 5586 23899 5642 23902
rect 5694 23899 5750 23902
rect 5802 23899 5858 23902
rect 5910 23899 5966 23902
rect 6018 23899 6074 23902
rect 6126 23899 6836 23902
rect 6888 23899 6944 23902
rect 6996 23899 7052 23902
rect 7104 23899 7160 23902
rect 7212 23899 7268 23902
rect 7320 23899 7376 23902
rect 7428 23899 7484 23902
rect 7536 23899 7592 23902
rect 7644 23899 7700 23902
rect 7752 23899 7808 23902
rect 7860 23899 7916 23902
rect 7968 23899 8024 23902
rect 8076 23899 8132 23902
rect 8184 23899 8240 23902
rect 8292 23899 8348 23902
rect 8400 23899 8456 23902
rect 8508 23899 8564 23902
rect 8616 23899 8672 23902
rect 8724 23899 8780 23902
rect 8832 23899 9206 23902
rect 9258 23899 9314 23902
rect 9366 23899 9422 23902
rect 9474 23899 9530 23902
rect 9582 23899 9638 23902
rect 9690 23899 9746 23902
rect 9798 23899 9854 23902
rect 9906 23899 9962 23902
rect 10014 23899 10070 23902
rect 10122 23899 10178 23902
rect 10230 23899 10286 23902
rect 10338 23899 10394 23902
rect 10446 23899 10502 23902
rect 10554 23899 10610 23902
rect 10662 23899 10718 23902
rect 10770 23899 10826 23902
rect 10878 23899 10934 23902
rect 10986 23899 11042 23902
rect 11094 23899 11150 23902
rect 11202 23899 11481 23902
rect 1481 23887 11481 23899
rect 11549 23887 11749 24053
rect 1213 23835 1233 23887
rect 1285 23835 1341 23887
rect 1393 23835 1413 23887
rect 1213 23808 1413 23835
rect 1213 23779 1256 23808
rect 1213 23727 1233 23779
rect 1213 23671 1256 23727
rect 1213 23619 1233 23671
rect 1213 23563 1256 23619
rect 1213 23511 1233 23563
rect 1213 23455 1256 23511
rect 1213 23403 1233 23455
rect 1213 23347 1256 23403
rect 1213 23295 1233 23347
rect 1213 23239 1256 23295
rect 1213 23187 1233 23239
rect 1213 23131 1256 23187
rect 1213 23079 1233 23131
rect 1213 23023 1256 23079
rect 1213 22971 1233 23023
rect 1213 22915 1256 22971
rect 1213 22863 1233 22915
rect 1213 22807 1256 22863
rect 1213 22755 1233 22807
rect 1213 22699 1256 22755
rect 1213 22647 1233 22699
rect 1213 22591 1256 22647
rect 1213 22539 1233 22591
rect 1213 22483 1256 22539
rect 1213 22431 1233 22483
rect 1213 22375 1256 22431
rect 1213 22323 1233 22375
rect 1213 22267 1256 22323
rect 1213 22215 1233 22267
rect 1213 22159 1256 22215
rect 1213 22107 1233 22159
rect 1213 22051 1256 22107
rect 1213 21999 1233 22051
rect 1213 21943 1256 21999
rect 1213 21891 1233 21943
rect 1213 21835 1256 21891
rect 1213 21783 1233 21835
rect 1213 21727 1256 21783
rect 1213 21675 1233 21727
rect 1213 21619 1256 21675
rect 1213 21567 1233 21619
rect 1213 21511 1256 21567
rect 1213 21459 1233 21511
rect 1213 21403 1256 21459
rect 1213 21351 1233 21403
rect 1213 21295 1256 21351
rect 1213 21243 1233 21295
rect 1213 21187 1256 21243
rect 1213 21135 1233 21187
rect 1213 21079 1256 21135
rect 1213 21027 1233 21079
rect 1213 20971 1256 21027
rect 1213 20919 1233 20971
rect 1213 20863 1256 20919
rect 1213 20811 1233 20863
rect 1213 20755 1256 20811
rect 1213 20703 1233 20755
rect 1213 20647 1256 20703
rect 1213 20595 1233 20647
rect 1213 20539 1256 20595
rect 1213 20487 1233 20539
rect 1213 20431 1256 20487
rect 1213 20379 1233 20431
rect 1213 20323 1256 20379
rect 1213 20271 1233 20323
rect 1213 20215 1256 20271
rect 1213 20163 1233 20215
rect 1213 20107 1256 20163
rect 1213 20055 1233 20107
rect 1213 19999 1256 20055
rect 1213 19947 1233 19999
rect 1213 19891 1256 19947
rect 1213 19839 1233 19891
rect 1213 19783 1256 19839
rect 1213 19731 1233 19783
rect 1213 19675 1256 19731
rect 1213 19623 1233 19675
rect 1213 19567 1256 19623
rect 1213 19515 1233 19567
rect 1213 19459 1256 19515
rect 1213 19407 1233 19459
rect 1213 19351 1256 19407
rect 1213 19299 1233 19351
rect 1213 19243 1256 19299
rect 1213 19191 1233 19243
rect 1213 19162 1256 19191
rect 1402 19162 1413 23808
rect 11549 23835 11569 23887
rect 11621 23835 11677 23887
rect 11729 23835 11749 23887
rect 11549 23808 11749 23835
rect 1481 23707 11481 23719
rect 1481 23655 1493 23707
rect 1545 23704 1601 23707
rect 1653 23704 3863 23707
rect 3915 23704 3971 23707
rect 4023 23704 6239 23707
rect 6291 23704 6347 23707
rect 6399 23704 6455 23707
rect 6507 23704 6563 23707
rect 6615 23704 6671 23707
rect 6723 23704 8939 23707
rect 8991 23704 9047 23707
rect 9099 23704 11309 23707
rect 11361 23704 11417 23707
rect 1545 23655 1601 23658
rect 1653 23655 3863 23658
rect 3915 23655 3971 23658
rect 4023 23655 6239 23658
rect 6291 23655 6347 23658
rect 6399 23655 6455 23658
rect 6507 23655 6563 23658
rect 6615 23655 6671 23658
rect 6723 23655 8939 23658
rect 8991 23655 9047 23658
rect 9099 23655 11309 23658
rect 11361 23655 11417 23658
rect 11469 23655 11481 23707
rect 1481 23643 11481 23655
rect 1481 23463 11481 23475
rect 1481 23460 1760 23463
rect 1812 23460 1868 23463
rect 1920 23460 1976 23463
rect 2028 23460 2084 23463
rect 2136 23460 2192 23463
rect 2244 23460 2300 23463
rect 2352 23460 2408 23463
rect 2460 23460 2516 23463
rect 2568 23460 2624 23463
rect 2676 23460 2732 23463
rect 2784 23460 2840 23463
rect 2892 23460 2948 23463
rect 3000 23460 3056 23463
rect 3108 23460 3164 23463
rect 3216 23460 3272 23463
rect 3324 23460 3380 23463
rect 3432 23460 3488 23463
rect 3540 23460 3596 23463
rect 3648 23460 3704 23463
rect 3756 23460 4130 23463
rect 4182 23460 4238 23463
rect 4290 23460 4346 23463
rect 4398 23460 4454 23463
rect 4506 23460 4562 23463
rect 4614 23460 4670 23463
rect 4722 23460 4778 23463
rect 4830 23460 4886 23463
rect 4938 23460 4994 23463
rect 5046 23460 5102 23463
rect 5154 23460 5210 23463
rect 5262 23460 5318 23463
rect 5370 23460 5426 23463
rect 5478 23460 5534 23463
rect 5586 23460 5642 23463
rect 5694 23460 5750 23463
rect 5802 23460 5858 23463
rect 5910 23460 5966 23463
rect 6018 23460 6074 23463
rect 6126 23460 6836 23463
rect 6888 23460 6944 23463
rect 6996 23460 7052 23463
rect 7104 23460 7160 23463
rect 7212 23460 7268 23463
rect 7320 23460 7376 23463
rect 7428 23460 7484 23463
rect 7536 23460 7592 23463
rect 7644 23460 7700 23463
rect 7752 23460 7808 23463
rect 7860 23460 7916 23463
rect 7968 23460 8024 23463
rect 8076 23460 8132 23463
rect 8184 23460 8240 23463
rect 8292 23460 8348 23463
rect 8400 23460 8456 23463
rect 8508 23460 8564 23463
rect 8616 23460 8672 23463
rect 8724 23460 8780 23463
rect 8832 23460 9206 23463
rect 9258 23460 9314 23463
rect 9366 23460 9422 23463
rect 9474 23460 9530 23463
rect 9582 23460 9638 23463
rect 9690 23460 9746 23463
rect 9798 23460 9854 23463
rect 9906 23460 9962 23463
rect 10014 23460 10070 23463
rect 10122 23460 10178 23463
rect 10230 23460 10286 23463
rect 10338 23460 10394 23463
rect 10446 23460 10502 23463
rect 10554 23460 10610 23463
rect 10662 23460 10718 23463
rect 10770 23460 10826 23463
rect 10878 23460 10934 23463
rect 10986 23460 11042 23463
rect 11094 23460 11150 23463
rect 11202 23460 11481 23463
rect 1481 23414 1494 23460
rect 11468 23414 11481 23460
rect 1481 23411 1760 23414
rect 1812 23411 1868 23414
rect 1920 23411 1976 23414
rect 2028 23411 2084 23414
rect 2136 23411 2192 23414
rect 2244 23411 2300 23414
rect 2352 23411 2408 23414
rect 2460 23411 2516 23414
rect 2568 23411 2624 23414
rect 2676 23411 2732 23414
rect 2784 23411 2840 23414
rect 2892 23411 2948 23414
rect 3000 23411 3056 23414
rect 3108 23411 3164 23414
rect 3216 23411 3272 23414
rect 3324 23411 3380 23414
rect 3432 23411 3488 23414
rect 3540 23411 3596 23414
rect 3648 23411 3704 23414
rect 3756 23411 4130 23414
rect 4182 23411 4238 23414
rect 4290 23411 4346 23414
rect 4398 23411 4454 23414
rect 4506 23411 4562 23414
rect 4614 23411 4670 23414
rect 4722 23411 4778 23414
rect 4830 23411 4886 23414
rect 4938 23411 4994 23414
rect 5046 23411 5102 23414
rect 5154 23411 5210 23414
rect 5262 23411 5318 23414
rect 5370 23411 5426 23414
rect 5478 23411 5534 23414
rect 5586 23411 5642 23414
rect 5694 23411 5750 23414
rect 5802 23411 5858 23414
rect 5910 23411 5966 23414
rect 6018 23411 6074 23414
rect 6126 23411 6836 23414
rect 6888 23411 6944 23414
rect 6996 23411 7052 23414
rect 7104 23411 7160 23414
rect 7212 23411 7268 23414
rect 7320 23411 7376 23414
rect 7428 23411 7484 23414
rect 7536 23411 7592 23414
rect 7644 23411 7700 23414
rect 7752 23411 7808 23414
rect 7860 23411 7916 23414
rect 7968 23411 8024 23414
rect 8076 23411 8132 23414
rect 8184 23411 8240 23414
rect 8292 23411 8348 23414
rect 8400 23411 8456 23414
rect 8508 23411 8564 23414
rect 8616 23411 8672 23414
rect 8724 23411 8780 23414
rect 8832 23411 9206 23414
rect 9258 23411 9314 23414
rect 9366 23411 9422 23414
rect 9474 23411 9530 23414
rect 9582 23411 9638 23414
rect 9690 23411 9746 23414
rect 9798 23411 9854 23414
rect 9906 23411 9962 23414
rect 10014 23411 10070 23414
rect 10122 23411 10178 23414
rect 10230 23411 10286 23414
rect 10338 23411 10394 23414
rect 10446 23411 10502 23414
rect 10554 23411 10610 23414
rect 10662 23411 10718 23414
rect 10770 23411 10826 23414
rect 10878 23411 10934 23414
rect 10986 23411 11042 23414
rect 11094 23411 11150 23414
rect 11202 23411 11481 23414
rect 1481 23399 11481 23411
rect 1481 23219 11481 23231
rect 1481 23167 1493 23219
rect 1545 23216 1601 23219
rect 1653 23216 3863 23219
rect 3915 23216 3971 23219
rect 4023 23216 6239 23219
rect 6291 23216 6347 23219
rect 6399 23216 6455 23219
rect 6507 23216 6563 23219
rect 6615 23216 6671 23219
rect 6723 23216 8939 23219
rect 8991 23216 9047 23219
rect 9099 23216 11309 23219
rect 11361 23216 11417 23219
rect 1545 23167 1601 23170
rect 1653 23167 3863 23170
rect 3915 23167 3971 23170
rect 4023 23167 6239 23170
rect 6291 23167 6347 23170
rect 6399 23167 6455 23170
rect 6507 23167 6563 23170
rect 6615 23167 6671 23170
rect 6723 23167 8939 23170
rect 8991 23167 9047 23170
rect 9099 23167 11309 23170
rect 11361 23167 11417 23170
rect 11469 23167 11481 23219
rect 1481 23155 11481 23167
rect 1481 22975 11481 22987
rect 1481 22972 1760 22975
rect 1812 22972 1868 22975
rect 1920 22972 1976 22975
rect 2028 22972 2084 22975
rect 2136 22972 2192 22975
rect 2244 22972 2300 22975
rect 2352 22972 2408 22975
rect 2460 22972 2516 22975
rect 2568 22972 2624 22975
rect 2676 22972 2732 22975
rect 2784 22972 2840 22975
rect 2892 22972 2948 22975
rect 3000 22972 3056 22975
rect 3108 22972 3164 22975
rect 3216 22972 3272 22975
rect 3324 22972 3380 22975
rect 3432 22972 3488 22975
rect 3540 22972 3596 22975
rect 3648 22972 3704 22975
rect 3756 22972 4130 22975
rect 4182 22972 4238 22975
rect 4290 22972 4346 22975
rect 4398 22972 4454 22975
rect 4506 22972 4562 22975
rect 4614 22972 4670 22975
rect 4722 22972 4778 22975
rect 4830 22972 4886 22975
rect 4938 22972 4994 22975
rect 5046 22972 5102 22975
rect 5154 22972 5210 22975
rect 5262 22972 5318 22975
rect 5370 22972 5426 22975
rect 5478 22972 5534 22975
rect 5586 22972 5642 22975
rect 5694 22972 5750 22975
rect 5802 22972 5858 22975
rect 5910 22972 5966 22975
rect 6018 22972 6074 22975
rect 6126 22972 6836 22975
rect 6888 22972 6944 22975
rect 6996 22972 7052 22975
rect 7104 22972 7160 22975
rect 7212 22972 7268 22975
rect 7320 22972 7376 22975
rect 7428 22972 7484 22975
rect 7536 22972 7592 22975
rect 7644 22972 7700 22975
rect 7752 22972 7808 22975
rect 7860 22972 7916 22975
rect 7968 22972 8024 22975
rect 8076 22972 8132 22975
rect 8184 22972 8240 22975
rect 8292 22972 8348 22975
rect 8400 22972 8456 22975
rect 8508 22972 8564 22975
rect 8616 22972 8672 22975
rect 8724 22972 8780 22975
rect 8832 22972 9206 22975
rect 9258 22972 9314 22975
rect 9366 22972 9422 22975
rect 9474 22972 9530 22975
rect 9582 22972 9638 22975
rect 9690 22972 9746 22975
rect 9798 22972 9854 22975
rect 9906 22972 9962 22975
rect 10014 22972 10070 22975
rect 10122 22972 10178 22975
rect 10230 22972 10286 22975
rect 10338 22972 10394 22975
rect 10446 22972 10502 22975
rect 10554 22972 10610 22975
rect 10662 22972 10718 22975
rect 10770 22972 10826 22975
rect 10878 22972 10934 22975
rect 10986 22972 11042 22975
rect 11094 22972 11150 22975
rect 11202 22972 11481 22975
rect 1481 22926 1494 22972
rect 11468 22926 11481 22972
rect 1481 22923 1760 22926
rect 1812 22923 1868 22926
rect 1920 22923 1976 22926
rect 2028 22923 2084 22926
rect 2136 22923 2192 22926
rect 2244 22923 2300 22926
rect 2352 22923 2408 22926
rect 2460 22923 2516 22926
rect 2568 22923 2624 22926
rect 2676 22923 2732 22926
rect 2784 22923 2840 22926
rect 2892 22923 2948 22926
rect 3000 22923 3056 22926
rect 3108 22923 3164 22926
rect 3216 22923 3272 22926
rect 3324 22923 3380 22926
rect 3432 22923 3488 22926
rect 3540 22923 3596 22926
rect 3648 22923 3704 22926
rect 3756 22923 4130 22926
rect 4182 22923 4238 22926
rect 4290 22923 4346 22926
rect 4398 22923 4454 22926
rect 4506 22923 4562 22926
rect 4614 22923 4670 22926
rect 4722 22923 4778 22926
rect 4830 22923 4886 22926
rect 4938 22923 4994 22926
rect 5046 22923 5102 22926
rect 5154 22923 5210 22926
rect 5262 22923 5318 22926
rect 5370 22923 5426 22926
rect 5478 22923 5534 22926
rect 5586 22923 5642 22926
rect 5694 22923 5750 22926
rect 5802 22923 5858 22926
rect 5910 22923 5966 22926
rect 6018 22923 6074 22926
rect 6126 22923 6836 22926
rect 6888 22923 6944 22926
rect 6996 22923 7052 22926
rect 7104 22923 7160 22926
rect 7212 22923 7268 22926
rect 7320 22923 7376 22926
rect 7428 22923 7484 22926
rect 7536 22923 7592 22926
rect 7644 22923 7700 22926
rect 7752 22923 7808 22926
rect 7860 22923 7916 22926
rect 7968 22923 8024 22926
rect 8076 22923 8132 22926
rect 8184 22923 8240 22926
rect 8292 22923 8348 22926
rect 8400 22923 8456 22926
rect 8508 22923 8564 22926
rect 8616 22923 8672 22926
rect 8724 22923 8780 22926
rect 8832 22923 9206 22926
rect 9258 22923 9314 22926
rect 9366 22923 9422 22926
rect 9474 22923 9530 22926
rect 9582 22923 9638 22926
rect 9690 22923 9746 22926
rect 9798 22923 9854 22926
rect 9906 22923 9962 22926
rect 10014 22923 10070 22926
rect 10122 22923 10178 22926
rect 10230 22923 10286 22926
rect 10338 22923 10394 22926
rect 10446 22923 10502 22926
rect 10554 22923 10610 22926
rect 10662 22923 10718 22926
rect 10770 22923 10826 22926
rect 10878 22923 10934 22926
rect 10986 22923 11042 22926
rect 11094 22923 11150 22926
rect 11202 22923 11481 22926
rect 1481 22911 11481 22923
rect 1481 22731 11481 22743
rect 1481 22679 1493 22731
rect 1545 22728 1601 22731
rect 1653 22728 3863 22731
rect 3915 22728 3971 22731
rect 4023 22728 6239 22731
rect 6291 22728 6347 22731
rect 6399 22728 6455 22731
rect 6507 22728 6563 22731
rect 6615 22728 6671 22731
rect 6723 22728 8939 22731
rect 8991 22728 9047 22731
rect 9099 22728 11309 22731
rect 11361 22728 11417 22731
rect 1545 22679 1601 22682
rect 1653 22679 3863 22682
rect 3915 22679 3971 22682
rect 4023 22679 6239 22682
rect 6291 22679 6347 22682
rect 6399 22679 6455 22682
rect 6507 22679 6563 22682
rect 6615 22679 6671 22682
rect 6723 22679 8939 22682
rect 8991 22679 9047 22682
rect 9099 22679 11309 22682
rect 11361 22679 11417 22682
rect 11469 22679 11481 22731
rect 1481 22667 11481 22679
rect 1481 22487 11481 22499
rect 1481 22484 1760 22487
rect 1812 22484 1868 22487
rect 1920 22484 1976 22487
rect 2028 22484 2084 22487
rect 2136 22484 2192 22487
rect 2244 22484 2300 22487
rect 2352 22484 2408 22487
rect 2460 22484 2516 22487
rect 2568 22484 2624 22487
rect 2676 22484 2732 22487
rect 2784 22484 2840 22487
rect 2892 22484 2948 22487
rect 3000 22484 3056 22487
rect 3108 22484 3164 22487
rect 3216 22484 3272 22487
rect 3324 22484 3380 22487
rect 3432 22484 3488 22487
rect 3540 22484 3596 22487
rect 3648 22484 3704 22487
rect 3756 22484 4130 22487
rect 4182 22484 4238 22487
rect 4290 22484 4346 22487
rect 4398 22484 4454 22487
rect 4506 22484 4562 22487
rect 4614 22484 4670 22487
rect 4722 22484 4778 22487
rect 4830 22484 4886 22487
rect 4938 22484 4994 22487
rect 5046 22484 5102 22487
rect 5154 22484 5210 22487
rect 5262 22484 5318 22487
rect 5370 22484 5426 22487
rect 5478 22484 5534 22487
rect 5586 22484 5642 22487
rect 5694 22484 5750 22487
rect 5802 22484 5858 22487
rect 5910 22484 5966 22487
rect 6018 22484 6074 22487
rect 6126 22484 6836 22487
rect 6888 22484 6944 22487
rect 6996 22484 7052 22487
rect 7104 22484 7160 22487
rect 7212 22484 7268 22487
rect 7320 22484 7376 22487
rect 7428 22484 7484 22487
rect 7536 22484 7592 22487
rect 7644 22484 7700 22487
rect 7752 22484 7808 22487
rect 7860 22484 7916 22487
rect 7968 22484 8024 22487
rect 8076 22484 8132 22487
rect 8184 22484 8240 22487
rect 8292 22484 8348 22487
rect 8400 22484 8456 22487
rect 8508 22484 8564 22487
rect 8616 22484 8672 22487
rect 8724 22484 8780 22487
rect 8832 22484 9206 22487
rect 9258 22484 9314 22487
rect 9366 22484 9422 22487
rect 9474 22484 9530 22487
rect 9582 22484 9638 22487
rect 9690 22484 9746 22487
rect 9798 22484 9854 22487
rect 9906 22484 9962 22487
rect 10014 22484 10070 22487
rect 10122 22484 10178 22487
rect 10230 22484 10286 22487
rect 10338 22484 10394 22487
rect 10446 22484 10502 22487
rect 10554 22484 10610 22487
rect 10662 22484 10718 22487
rect 10770 22484 10826 22487
rect 10878 22484 10934 22487
rect 10986 22484 11042 22487
rect 11094 22484 11150 22487
rect 11202 22484 11481 22487
rect 1481 22438 1494 22484
rect 11468 22438 11481 22484
rect 1481 22435 1760 22438
rect 1812 22435 1868 22438
rect 1920 22435 1976 22438
rect 2028 22435 2084 22438
rect 2136 22435 2192 22438
rect 2244 22435 2300 22438
rect 2352 22435 2408 22438
rect 2460 22435 2516 22438
rect 2568 22435 2624 22438
rect 2676 22435 2732 22438
rect 2784 22435 2840 22438
rect 2892 22435 2948 22438
rect 3000 22435 3056 22438
rect 3108 22435 3164 22438
rect 3216 22435 3272 22438
rect 3324 22435 3380 22438
rect 3432 22435 3488 22438
rect 3540 22435 3596 22438
rect 3648 22435 3704 22438
rect 3756 22435 4130 22438
rect 4182 22435 4238 22438
rect 4290 22435 4346 22438
rect 4398 22435 4454 22438
rect 4506 22435 4562 22438
rect 4614 22435 4670 22438
rect 4722 22435 4778 22438
rect 4830 22435 4886 22438
rect 4938 22435 4994 22438
rect 5046 22435 5102 22438
rect 5154 22435 5210 22438
rect 5262 22435 5318 22438
rect 5370 22435 5426 22438
rect 5478 22435 5534 22438
rect 5586 22435 5642 22438
rect 5694 22435 5750 22438
rect 5802 22435 5858 22438
rect 5910 22435 5966 22438
rect 6018 22435 6074 22438
rect 6126 22435 6836 22438
rect 6888 22435 6944 22438
rect 6996 22435 7052 22438
rect 7104 22435 7160 22438
rect 7212 22435 7268 22438
rect 7320 22435 7376 22438
rect 7428 22435 7484 22438
rect 7536 22435 7592 22438
rect 7644 22435 7700 22438
rect 7752 22435 7808 22438
rect 7860 22435 7916 22438
rect 7968 22435 8024 22438
rect 8076 22435 8132 22438
rect 8184 22435 8240 22438
rect 8292 22435 8348 22438
rect 8400 22435 8456 22438
rect 8508 22435 8564 22438
rect 8616 22435 8672 22438
rect 8724 22435 8780 22438
rect 8832 22435 9206 22438
rect 9258 22435 9314 22438
rect 9366 22435 9422 22438
rect 9474 22435 9530 22438
rect 9582 22435 9638 22438
rect 9690 22435 9746 22438
rect 9798 22435 9854 22438
rect 9906 22435 9962 22438
rect 10014 22435 10070 22438
rect 10122 22435 10178 22438
rect 10230 22435 10286 22438
rect 10338 22435 10394 22438
rect 10446 22435 10502 22438
rect 10554 22435 10610 22438
rect 10662 22435 10718 22438
rect 10770 22435 10826 22438
rect 10878 22435 10934 22438
rect 10986 22435 11042 22438
rect 11094 22435 11150 22438
rect 11202 22435 11481 22438
rect 1481 22423 11481 22435
rect 1481 22243 11481 22255
rect 1481 22191 1493 22243
rect 1545 22240 1601 22243
rect 1653 22240 3863 22243
rect 3915 22240 3971 22243
rect 4023 22240 6239 22243
rect 6291 22240 6347 22243
rect 6399 22240 6455 22243
rect 6507 22240 6563 22243
rect 6615 22240 6671 22243
rect 6723 22240 8939 22243
rect 8991 22240 9047 22243
rect 9099 22240 11309 22243
rect 11361 22240 11417 22243
rect 1545 22191 1601 22194
rect 1653 22191 3863 22194
rect 3915 22191 3971 22194
rect 4023 22191 6239 22194
rect 6291 22191 6347 22194
rect 6399 22191 6455 22194
rect 6507 22191 6563 22194
rect 6615 22191 6671 22194
rect 6723 22191 8939 22194
rect 8991 22191 9047 22194
rect 9099 22191 11309 22194
rect 11361 22191 11417 22194
rect 11469 22191 11481 22243
rect 1481 22179 11481 22191
rect 1481 21999 11481 22011
rect 1481 21996 1760 21999
rect 1812 21996 1868 21999
rect 1920 21996 1976 21999
rect 2028 21996 2084 21999
rect 2136 21996 2192 21999
rect 2244 21996 2300 21999
rect 2352 21996 2408 21999
rect 2460 21996 2516 21999
rect 2568 21996 2624 21999
rect 2676 21996 2732 21999
rect 2784 21996 2840 21999
rect 2892 21996 2948 21999
rect 3000 21996 3056 21999
rect 3108 21996 3164 21999
rect 3216 21996 3272 21999
rect 3324 21996 3380 21999
rect 3432 21996 3488 21999
rect 3540 21996 3596 21999
rect 3648 21996 3704 21999
rect 3756 21996 4130 21999
rect 4182 21996 4238 21999
rect 4290 21996 4346 21999
rect 4398 21996 4454 21999
rect 4506 21996 4562 21999
rect 4614 21996 4670 21999
rect 4722 21996 4778 21999
rect 4830 21996 4886 21999
rect 4938 21996 4994 21999
rect 5046 21996 5102 21999
rect 5154 21996 5210 21999
rect 5262 21996 5318 21999
rect 5370 21996 5426 21999
rect 5478 21996 5534 21999
rect 5586 21996 5642 21999
rect 5694 21996 5750 21999
rect 5802 21996 5858 21999
rect 5910 21996 5966 21999
rect 6018 21996 6074 21999
rect 6126 21996 6836 21999
rect 6888 21996 6944 21999
rect 6996 21996 7052 21999
rect 7104 21996 7160 21999
rect 7212 21996 7268 21999
rect 7320 21996 7376 21999
rect 7428 21996 7484 21999
rect 7536 21996 7592 21999
rect 7644 21996 7700 21999
rect 7752 21996 7808 21999
rect 7860 21996 7916 21999
rect 7968 21996 8024 21999
rect 8076 21996 8132 21999
rect 8184 21996 8240 21999
rect 8292 21996 8348 21999
rect 8400 21996 8456 21999
rect 8508 21996 8564 21999
rect 8616 21996 8672 21999
rect 8724 21996 8780 21999
rect 8832 21996 9206 21999
rect 9258 21996 9314 21999
rect 9366 21996 9422 21999
rect 9474 21996 9530 21999
rect 9582 21996 9638 21999
rect 9690 21996 9746 21999
rect 9798 21996 9854 21999
rect 9906 21996 9962 21999
rect 10014 21996 10070 21999
rect 10122 21996 10178 21999
rect 10230 21996 10286 21999
rect 10338 21996 10394 21999
rect 10446 21996 10502 21999
rect 10554 21996 10610 21999
rect 10662 21996 10718 21999
rect 10770 21996 10826 21999
rect 10878 21996 10934 21999
rect 10986 21996 11042 21999
rect 11094 21996 11150 21999
rect 11202 21996 11481 21999
rect 1481 21950 1494 21996
rect 11468 21950 11481 21996
rect 1481 21947 1760 21950
rect 1812 21947 1868 21950
rect 1920 21947 1976 21950
rect 2028 21947 2084 21950
rect 2136 21947 2192 21950
rect 2244 21947 2300 21950
rect 2352 21947 2408 21950
rect 2460 21947 2516 21950
rect 2568 21947 2624 21950
rect 2676 21947 2732 21950
rect 2784 21947 2840 21950
rect 2892 21947 2948 21950
rect 3000 21947 3056 21950
rect 3108 21947 3164 21950
rect 3216 21947 3272 21950
rect 3324 21947 3380 21950
rect 3432 21947 3488 21950
rect 3540 21947 3596 21950
rect 3648 21947 3704 21950
rect 3756 21947 4130 21950
rect 4182 21947 4238 21950
rect 4290 21947 4346 21950
rect 4398 21947 4454 21950
rect 4506 21947 4562 21950
rect 4614 21947 4670 21950
rect 4722 21947 4778 21950
rect 4830 21947 4886 21950
rect 4938 21947 4994 21950
rect 5046 21947 5102 21950
rect 5154 21947 5210 21950
rect 5262 21947 5318 21950
rect 5370 21947 5426 21950
rect 5478 21947 5534 21950
rect 5586 21947 5642 21950
rect 5694 21947 5750 21950
rect 5802 21947 5858 21950
rect 5910 21947 5966 21950
rect 6018 21947 6074 21950
rect 6126 21947 6836 21950
rect 6888 21947 6944 21950
rect 6996 21947 7052 21950
rect 7104 21947 7160 21950
rect 7212 21947 7268 21950
rect 7320 21947 7376 21950
rect 7428 21947 7484 21950
rect 7536 21947 7592 21950
rect 7644 21947 7700 21950
rect 7752 21947 7808 21950
rect 7860 21947 7916 21950
rect 7968 21947 8024 21950
rect 8076 21947 8132 21950
rect 8184 21947 8240 21950
rect 8292 21947 8348 21950
rect 8400 21947 8456 21950
rect 8508 21947 8564 21950
rect 8616 21947 8672 21950
rect 8724 21947 8780 21950
rect 8832 21947 9206 21950
rect 9258 21947 9314 21950
rect 9366 21947 9422 21950
rect 9474 21947 9530 21950
rect 9582 21947 9638 21950
rect 9690 21947 9746 21950
rect 9798 21947 9854 21950
rect 9906 21947 9962 21950
rect 10014 21947 10070 21950
rect 10122 21947 10178 21950
rect 10230 21947 10286 21950
rect 10338 21947 10394 21950
rect 10446 21947 10502 21950
rect 10554 21947 10610 21950
rect 10662 21947 10718 21950
rect 10770 21947 10826 21950
rect 10878 21947 10934 21950
rect 10986 21947 11042 21950
rect 11094 21947 11150 21950
rect 11202 21947 11481 21950
rect 1481 21935 11481 21947
rect 1481 21755 11481 21767
rect 1481 21703 1493 21755
rect 1545 21752 1601 21755
rect 1653 21752 3863 21755
rect 3915 21752 3971 21755
rect 4023 21752 6239 21755
rect 6291 21752 6347 21755
rect 6399 21752 6455 21755
rect 6507 21752 6563 21755
rect 6615 21752 6671 21755
rect 6723 21752 8939 21755
rect 8991 21752 9047 21755
rect 9099 21752 11309 21755
rect 11361 21752 11417 21755
rect 1545 21703 1601 21706
rect 1653 21703 3863 21706
rect 3915 21703 3971 21706
rect 4023 21703 6239 21706
rect 6291 21703 6347 21706
rect 6399 21703 6455 21706
rect 6507 21703 6563 21706
rect 6615 21703 6671 21706
rect 6723 21703 8939 21706
rect 8991 21703 9047 21706
rect 9099 21703 11309 21706
rect 11361 21703 11417 21706
rect 11469 21703 11481 21755
rect 1481 21691 11481 21703
rect 1481 21511 11481 21523
rect 1481 21508 1760 21511
rect 1812 21508 1868 21511
rect 1920 21508 1976 21511
rect 2028 21508 2084 21511
rect 2136 21508 2192 21511
rect 2244 21508 2300 21511
rect 2352 21508 2408 21511
rect 2460 21508 2516 21511
rect 2568 21508 2624 21511
rect 2676 21508 2732 21511
rect 2784 21508 2840 21511
rect 2892 21508 2948 21511
rect 3000 21508 3056 21511
rect 3108 21508 3164 21511
rect 3216 21508 3272 21511
rect 3324 21508 3380 21511
rect 3432 21508 3488 21511
rect 3540 21508 3596 21511
rect 3648 21508 3704 21511
rect 3756 21508 4130 21511
rect 4182 21508 4238 21511
rect 4290 21508 4346 21511
rect 4398 21508 4454 21511
rect 4506 21508 4562 21511
rect 4614 21508 4670 21511
rect 4722 21508 4778 21511
rect 4830 21508 4886 21511
rect 4938 21508 4994 21511
rect 5046 21508 5102 21511
rect 5154 21508 5210 21511
rect 5262 21508 5318 21511
rect 5370 21508 5426 21511
rect 5478 21508 5534 21511
rect 5586 21508 5642 21511
rect 5694 21508 5750 21511
rect 5802 21508 5858 21511
rect 5910 21508 5966 21511
rect 6018 21508 6074 21511
rect 6126 21508 6836 21511
rect 6888 21508 6944 21511
rect 6996 21508 7052 21511
rect 7104 21508 7160 21511
rect 7212 21508 7268 21511
rect 7320 21508 7376 21511
rect 7428 21508 7484 21511
rect 7536 21508 7592 21511
rect 7644 21508 7700 21511
rect 7752 21508 7808 21511
rect 7860 21508 7916 21511
rect 7968 21508 8024 21511
rect 8076 21508 8132 21511
rect 8184 21508 8240 21511
rect 8292 21508 8348 21511
rect 8400 21508 8456 21511
rect 8508 21508 8564 21511
rect 8616 21508 8672 21511
rect 8724 21508 8780 21511
rect 8832 21508 9206 21511
rect 9258 21508 9314 21511
rect 9366 21508 9422 21511
rect 9474 21508 9530 21511
rect 9582 21508 9638 21511
rect 9690 21508 9746 21511
rect 9798 21508 9854 21511
rect 9906 21508 9962 21511
rect 10014 21508 10070 21511
rect 10122 21508 10178 21511
rect 10230 21508 10286 21511
rect 10338 21508 10394 21511
rect 10446 21508 10502 21511
rect 10554 21508 10610 21511
rect 10662 21508 10718 21511
rect 10770 21508 10826 21511
rect 10878 21508 10934 21511
rect 10986 21508 11042 21511
rect 11094 21508 11150 21511
rect 11202 21508 11481 21511
rect 1481 21462 1494 21508
rect 11468 21462 11481 21508
rect 1481 21459 1760 21462
rect 1812 21459 1868 21462
rect 1920 21459 1976 21462
rect 2028 21459 2084 21462
rect 2136 21459 2192 21462
rect 2244 21459 2300 21462
rect 2352 21459 2408 21462
rect 2460 21459 2516 21462
rect 2568 21459 2624 21462
rect 2676 21459 2732 21462
rect 2784 21459 2840 21462
rect 2892 21459 2948 21462
rect 3000 21459 3056 21462
rect 3108 21459 3164 21462
rect 3216 21459 3272 21462
rect 3324 21459 3380 21462
rect 3432 21459 3488 21462
rect 3540 21459 3596 21462
rect 3648 21459 3704 21462
rect 3756 21459 4130 21462
rect 4182 21459 4238 21462
rect 4290 21459 4346 21462
rect 4398 21459 4454 21462
rect 4506 21459 4562 21462
rect 4614 21459 4670 21462
rect 4722 21459 4778 21462
rect 4830 21459 4886 21462
rect 4938 21459 4994 21462
rect 5046 21459 5102 21462
rect 5154 21459 5210 21462
rect 5262 21459 5318 21462
rect 5370 21459 5426 21462
rect 5478 21459 5534 21462
rect 5586 21459 5642 21462
rect 5694 21459 5750 21462
rect 5802 21459 5858 21462
rect 5910 21459 5966 21462
rect 6018 21459 6074 21462
rect 6126 21459 6836 21462
rect 6888 21459 6944 21462
rect 6996 21459 7052 21462
rect 7104 21459 7160 21462
rect 7212 21459 7268 21462
rect 7320 21459 7376 21462
rect 7428 21459 7484 21462
rect 7536 21459 7592 21462
rect 7644 21459 7700 21462
rect 7752 21459 7808 21462
rect 7860 21459 7916 21462
rect 7968 21459 8024 21462
rect 8076 21459 8132 21462
rect 8184 21459 8240 21462
rect 8292 21459 8348 21462
rect 8400 21459 8456 21462
rect 8508 21459 8564 21462
rect 8616 21459 8672 21462
rect 8724 21459 8780 21462
rect 8832 21459 9206 21462
rect 9258 21459 9314 21462
rect 9366 21459 9422 21462
rect 9474 21459 9530 21462
rect 9582 21459 9638 21462
rect 9690 21459 9746 21462
rect 9798 21459 9854 21462
rect 9906 21459 9962 21462
rect 10014 21459 10070 21462
rect 10122 21459 10178 21462
rect 10230 21459 10286 21462
rect 10338 21459 10394 21462
rect 10446 21459 10502 21462
rect 10554 21459 10610 21462
rect 10662 21459 10718 21462
rect 10770 21459 10826 21462
rect 10878 21459 10934 21462
rect 10986 21459 11042 21462
rect 11094 21459 11150 21462
rect 11202 21459 11481 21462
rect 1481 21447 11481 21459
rect 1481 21267 11481 21279
rect 1481 21215 1493 21267
rect 1545 21264 1601 21267
rect 1653 21264 3863 21267
rect 3915 21264 3971 21267
rect 4023 21264 6239 21267
rect 6291 21264 6347 21267
rect 6399 21264 6455 21267
rect 6507 21264 6563 21267
rect 6615 21264 6671 21267
rect 6723 21264 8939 21267
rect 8991 21264 9047 21267
rect 9099 21264 11309 21267
rect 11361 21264 11417 21267
rect 1545 21215 1601 21218
rect 1653 21215 3863 21218
rect 3915 21215 3971 21218
rect 4023 21215 6239 21218
rect 6291 21215 6347 21218
rect 6399 21215 6455 21218
rect 6507 21215 6563 21218
rect 6615 21215 6671 21218
rect 6723 21215 8939 21218
rect 8991 21215 9047 21218
rect 9099 21215 11309 21218
rect 11361 21215 11417 21218
rect 11469 21215 11481 21267
rect 1481 21203 11481 21215
rect 1481 21023 11481 21035
rect 1481 21020 1760 21023
rect 1812 21020 1868 21023
rect 1920 21020 1976 21023
rect 2028 21020 2084 21023
rect 2136 21020 2192 21023
rect 2244 21020 2300 21023
rect 2352 21020 2408 21023
rect 2460 21020 2516 21023
rect 2568 21020 2624 21023
rect 2676 21020 2732 21023
rect 2784 21020 2840 21023
rect 2892 21020 2948 21023
rect 3000 21020 3056 21023
rect 3108 21020 3164 21023
rect 3216 21020 3272 21023
rect 3324 21020 3380 21023
rect 3432 21020 3488 21023
rect 3540 21020 3596 21023
rect 3648 21020 3704 21023
rect 3756 21020 4130 21023
rect 4182 21020 4238 21023
rect 4290 21020 4346 21023
rect 4398 21020 4454 21023
rect 4506 21020 4562 21023
rect 4614 21020 4670 21023
rect 4722 21020 4778 21023
rect 4830 21020 4886 21023
rect 4938 21020 4994 21023
rect 5046 21020 5102 21023
rect 5154 21020 5210 21023
rect 5262 21020 5318 21023
rect 5370 21020 5426 21023
rect 5478 21020 5534 21023
rect 5586 21020 5642 21023
rect 5694 21020 5750 21023
rect 5802 21020 5858 21023
rect 5910 21020 5966 21023
rect 6018 21020 6074 21023
rect 6126 21020 6836 21023
rect 6888 21020 6944 21023
rect 6996 21020 7052 21023
rect 7104 21020 7160 21023
rect 7212 21020 7268 21023
rect 7320 21020 7376 21023
rect 7428 21020 7484 21023
rect 7536 21020 7592 21023
rect 7644 21020 7700 21023
rect 7752 21020 7808 21023
rect 7860 21020 7916 21023
rect 7968 21020 8024 21023
rect 8076 21020 8132 21023
rect 8184 21020 8240 21023
rect 8292 21020 8348 21023
rect 8400 21020 8456 21023
rect 8508 21020 8564 21023
rect 8616 21020 8672 21023
rect 8724 21020 8780 21023
rect 8832 21020 9206 21023
rect 9258 21020 9314 21023
rect 9366 21020 9422 21023
rect 9474 21020 9530 21023
rect 9582 21020 9638 21023
rect 9690 21020 9746 21023
rect 9798 21020 9854 21023
rect 9906 21020 9962 21023
rect 10014 21020 10070 21023
rect 10122 21020 10178 21023
rect 10230 21020 10286 21023
rect 10338 21020 10394 21023
rect 10446 21020 10502 21023
rect 10554 21020 10610 21023
rect 10662 21020 10718 21023
rect 10770 21020 10826 21023
rect 10878 21020 10934 21023
rect 10986 21020 11042 21023
rect 11094 21020 11150 21023
rect 11202 21020 11481 21023
rect 1481 20974 1494 21020
rect 11468 20974 11481 21020
rect 1481 20971 1760 20974
rect 1812 20971 1868 20974
rect 1920 20971 1976 20974
rect 2028 20971 2084 20974
rect 2136 20971 2192 20974
rect 2244 20971 2300 20974
rect 2352 20971 2408 20974
rect 2460 20971 2516 20974
rect 2568 20971 2624 20974
rect 2676 20971 2732 20974
rect 2784 20971 2840 20974
rect 2892 20971 2948 20974
rect 3000 20971 3056 20974
rect 3108 20971 3164 20974
rect 3216 20971 3272 20974
rect 3324 20971 3380 20974
rect 3432 20971 3488 20974
rect 3540 20971 3596 20974
rect 3648 20971 3704 20974
rect 3756 20971 4130 20974
rect 4182 20971 4238 20974
rect 4290 20971 4346 20974
rect 4398 20971 4454 20974
rect 4506 20971 4562 20974
rect 4614 20971 4670 20974
rect 4722 20971 4778 20974
rect 4830 20971 4886 20974
rect 4938 20971 4994 20974
rect 5046 20971 5102 20974
rect 5154 20971 5210 20974
rect 5262 20971 5318 20974
rect 5370 20971 5426 20974
rect 5478 20971 5534 20974
rect 5586 20971 5642 20974
rect 5694 20971 5750 20974
rect 5802 20971 5858 20974
rect 5910 20971 5966 20974
rect 6018 20971 6074 20974
rect 6126 20971 6836 20974
rect 6888 20971 6944 20974
rect 6996 20971 7052 20974
rect 7104 20971 7160 20974
rect 7212 20971 7268 20974
rect 7320 20971 7376 20974
rect 7428 20971 7484 20974
rect 7536 20971 7592 20974
rect 7644 20971 7700 20974
rect 7752 20971 7808 20974
rect 7860 20971 7916 20974
rect 7968 20971 8024 20974
rect 8076 20971 8132 20974
rect 8184 20971 8240 20974
rect 8292 20971 8348 20974
rect 8400 20971 8456 20974
rect 8508 20971 8564 20974
rect 8616 20971 8672 20974
rect 8724 20971 8780 20974
rect 8832 20971 9206 20974
rect 9258 20971 9314 20974
rect 9366 20971 9422 20974
rect 9474 20971 9530 20974
rect 9582 20971 9638 20974
rect 9690 20971 9746 20974
rect 9798 20971 9854 20974
rect 9906 20971 9962 20974
rect 10014 20971 10070 20974
rect 10122 20971 10178 20974
rect 10230 20971 10286 20974
rect 10338 20971 10394 20974
rect 10446 20971 10502 20974
rect 10554 20971 10610 20974
rect 10662 20971 10718 20974
rect 10770 20971 10826 20974
rect 10878 20971 10934 20974
rect 10986 20971 11042 20974
rect 11094 20971 11150 20974
rect 11202 20971 11481 20974
rect 1481 20959 11481 20971
rect 1481 20779 11481 20791
rect 1481 20727 1493 20779
rect 1545 20776 1601 20779
rect 1653 20776 3863 20779
rect 3915 20776 3971 20779
rect 4023 20776 6239 20779
rect 6291 20776 6347 20779
rect 6399 20776 6455 20779
rect 6507 20776 6563 20779
rect 6615 20776 6671 20779
rect 6723 20776 8939 20779
rect 8991 20776 9047 20779
rect 9099 20776 11309 20779
rect 11361 20776 11417 20779
rect 1545 20727 1601 20730
rect 1653 20727 3863 20730
rect 3915 20727 3971 20730
rect 4023 20727 6239 20730
rect 6291 20727 6347 20730
rect 6399 20727 6455 20730
rect 6507 20727 6563 20730
rect 6615 20727 6671 20730
rect 6723 20727 8939 20730
rect 8991 20727 9047 20730
rect 9099 20727 11309 20730
rect 11361 20727 11417 20730
rect 11469 20727 11481 20779
rect 1481 20715 11481 20727
rect 1481 20535 11481 20547
rect 1481 20532 1760 20535
rect 1812 20532 1868 20535
rect 1920 20532 1976 20535
rect 2028 20532 2084 20535
rect 2136 20532 2192 20535
rect 2244 20532 2300 20535
rect 2352 20532 2408 20535
rect 2460 20532 2516 20535
rect 2568 20532 2624 20535
rect 2676 20532 2732 20535
rect 2784 20532 2840 20535
rect 2892 20532 2948 20535
rect 3000 20532 3056 20535
rect 3108 20532 3164 20535
rect 3216 20532 3272 20535
rect 3324 20532 3380 20535
rect 3432 20532 3488 20535
rect 3540 20532 3596 20535
rect 3648 20532 3704 20535
rect 3756 20532 4130 20535
rect 4182 20532 4238 20535
rect 4290 20532 4346 20535
rect 4398 20532 4454 20535
rect 4506 20532 4562 20535
rect 4614 20532 4670 20535
rect 4722 20532 4778 20535
rect 4830 20532 4886 20535
rect 4938 20532 4994 20535
rect 5046 20532 5102 20535
rect 5154 20532 5210 20535
rect 5262 20532 5318 20535
rect 5370 20532 5426 20535
rect 5478 20532 5534 20535
rect 5586 20532 5642 20535
rect 5694 20532 5750 20535
rect 5802 20532 5858 20535
rect 5910 20532 5966 20535
rect 6018 20532 6074 20535
rect 6126 20532 6836 20535
rect 6888 20532 6944 20535
rect 6996 20532 7052 20535
rect 7104 20532 7160 20535
rect 7212 20532 7268 20535
rect 7320 20532 7376 20535
rect 7428 20532 7484 20535
rect 7536 20532 7592 20535
rect 7644 20532 7700 20535
rect 7752 20532 7808 20535
rect 7860 20532 7916 20535
rect 7968 20532 8024 20535
rect 8076 20532 8132 20535
rect 8184 20532 8240 20535
rect 8292 20532 8348 20535
rect 8400 20532 8456 20535
rect 8508 20532 8564 20535
rect 8616 20532 8672 20535
rect 8724 20532 8780 20535
rect 8832 20532 9206 20535
rect 9258 20532 9314 20535
rect 9366 20532 9422 20535
rect 9474 20532 9530 20535
rect 9582 20532 9638 20535
rect 9690 20532 9746 20535
rect 9798 20532 9854 20535
rect 9906 20532 9962 20535
rect 10014 20532 10070 20535
rect 10122 20532 10178 20535
rect 10230 20532 10286 20535
rect 10338 20532 10394 20535
rect 10446 20532 10502 20535
rect 10554 20532 10610 20535
rect 10662 20532 10718 20535
rect 10770 20532 10826 20535
rect 10878 20532 10934 20535
rect 10986 20532 11042 20535
rect 11094 20532 11150 20535
rect 11202 20532 11481 20535
rect 1481 20486 1494 20532
rect 11468 20486 11481 20532
rect 1481 20483 1760 20486
rect 1812 20483 1868 20486
rect 1920 20483 1976 20486
rect 2028 20483 2084 20486
rect 2136 20483 2192 20486
rect 2244 20483 2300 20486
rect 2352 20483 2408 20486
rect 2460 20483 2516 20486
rect 2568 20483 2624 20486
rect 2676 20483 2732 20486
rect 2784 20483 2840 20486
rect 2892 20483 2948 20486
rect 3000 20483 3056 20486
rect 3108 20483 3164 20486
rect 3216 20483 3272 20486
rect 3324 20483 3380 20486
rect 3432 20483 3488 20486
rect 3540 20483 3596 20486
rect 3648 20483 3704 20486
rect 3756 20483 4130 20486
rect 4182 20483 4238 20486
rect 4290 20483 4346 20486
rect 4398 20483 4454 20486
rect 4506 20483 4562 20486
rect 4614 20483 4670 20486
rect 4722 20483 4778 20486
rect 4830 20483 4886 20486
rect 4938 20483 4994 20486
rect 5046 20483 5102 20486
rect 5154 20483 5210 20486
rect 5262 20483 5318 20486
rect 5370 20483 5426 20486
rect 5478 20483 5534 20486
rect 5586 20483 5642 20486
rect 5694 20483 5750 20486
rect 5802 20483 5858 20486
rect 5910 20483 5966 20486
rect 6018 20483 6074 20486
rect 6126 20483 6836 20486
rect 6888 20483 6944 20486
rect 6996 20483 7052 20486
rect 7104 20483 7160 20486
rect 7212 20483 7268 20486
rect 7320 20483 7376 20486
rect 7428 20483 7484 20486
rect 7536 20483 7592 20486
rect 7644 20483 7700 20486
rect 7752 20483 7808 20486
rect 7860 20483 7916 20486
rect 7968 20483 8024 20486
rect 8076 20483 8132 20486
rect 8184 20483 8240 20486
rect 8292 20483 8348 20486
rect 8400 20483 8456 20486
rect 8508 20483 8564 20486
rect 8616 20483 8672 20486
rect 8724 20483 8780 20486
rect 8832 20483 9206 20486
rect 9258 20483 9314 20486
rect 9366 20483 9422 20486
rect 9474 20483 9530 20486
rect 9582 20483 9638 20486
rect 9690 20483 9746 20486
rect 9798 20483 9854 20486
rect 9906 20483 9962 20486
rect 10014 20483 10070 20486
rect 10122 20483 10178 20486
rect 10230 20483 10286 20486
rect 10338 20483 10394 20486
rect 10446 20483 10502 20486
rect 10554 20483 10610 20486
rect 10662 20483 10718 20486
rect 10770 20483 10826 20486
rect 10878 20483 10934 20486
rect 10986 20483 11042 20486
rect 11094 20483 11150 20486
rect 11202 20483 11481 20486
rect 1481 20471 11481 20483
rect 1481 20291 11481 20303
rect 1481 20239 1493 20291
rect 1545 20288 1601 20291
rect 1653 20288 3863 20291
rect 3915 20288 3971 20291
rect 4023 20288 6239 20291
rect 6291 20288 6347 20291
rect 6399 20288 6455 20291
rect 6507 20288 6563 20291
rect 6615 20288 6671 20291
rect 6723 20288 8939 20291
rect 8991 20288 9047 20291
rect 9099 20288 11309 20291
rect 11361 20288 11417 20291
rect 1545 20239 1601 20242
rect 1653 20239 3863 20242
rect 3915 20239 3971 20242
rect 4023 20239 6239 20242
rect 6291 20239 6347 20242
rect 6399 20239 6455 20242
rect 6507 20239 6563 20242
rect 6615 20239 6671 20242
rect 6723 20239 8939 20242
rect 8991 20239 9047 20242
rect 9099 20239 11309 20242
rect 11361 20239 11417 20242
rect 11469 20239 11481 20291
rect 1481 20227 11481 20239
rect 1481 20047 11481 20059
rect 1481 20044 1760 20047
rect 1812 20044 1868 20047
rect 1920 20044 1976 20047
rect 2028 20044 2084 20047
rect 2136 20044 2192 20047
rect 2244 20044 2300 20047
rect 2352 20044 2408 20047
rect 2460 20044 2516 20047
rect 2568 20044 2624 20047
rect 2676 20044 2732 20047
rect 2784 20044 2840 20047
rect 2892 20044 2948 20047
rect 3000 20044 3056 20047
rect 3108 20044 3164 20047
rect 3216 20044 3272 20047
rect 3324 20044 3380 20047
rect 3432 20044 3488 20047
rect 3540 20044 3596 20047
rect 3648 20044 3704 20047
rect 3756 20044 4130 20047
rect 4182 20044 4238 20047
rect 4290 20044 4346 20047
rect 4398 20044 4454 20047
rect 4506 20044 4562 20047
rect 4614 20044 4670 20047
rect 4722 20044 4778 20047
rect 4830 20044 4886 20047
rect 4938 20044 4994 20047
rect 5046 20044 5102 20047
rect 5154 20044 5210 20047
rect 5262 20044 5318 20047
rect 5370 20044 5426 20047
rect 5478 20044 5534 20047
rect 5586 20044 5642 20047
rect 5694 20044 5750 20047
rect 5802 20044 5858 20047
rect 5910 20044 5966 20047
rect 6018 20044 6074 20047
rect 6126 20044 6836 20047
rect 6888 20044 6944 20047
rect 6996 20044 7052 20047
rect 7104 20044 7160 20047
rect 7212 20044 7268 20047
rect 7320 20044 7376 20047
rect 7428 20044 7484 20047
rect 7536 20044 7592 20047
rect 7644 20044 7700 20047
rect 7752 20044 7808 20047
rect 7860 20044 7916 20047
rect 7968 20044 8024 20047
rect 8076 20044 8132 20047
rect 8184 20044 8240 20047
rect 8292 20044 8348 20047
rect 8400 20044 8456 20047
rect 8508 20044 8564 20047
rect 8616 20044 8672 20047
rect 8724 20044 8780 20047
rect 8832 20044 9206 20047
rect 9258 20044 9314 20047
rect 9366 20044 9422 20047
rect 9474 20044 9530 20047
rect 9582 20044 9638 20047
rect 9690 20044 9746 20047
rect 9798 20044 9854 20047
rect 9906 20044 9962 20047
rect 10014 20044 10070 20047
rect 10122 20044 10178 20047
rect 10230 20044 10286 20047
rect 10338 20044 10394 20047
rect 10446 20044 10502 20047
rect 10554 20044 10610 20047
rect 10662 20044 10718 20047
rect 10770 20044 10826 20047
rect 10878 20044 10934 20047
rect 10986 20044 11042 20047
rect 11094 20044 11150 20047
rect 11202 20044 11481 20047
rect 1481 19998 1494 20044
rect 11468 19998 11481 20044
rect 1481 19995 1760 19998
rect 1812 19995 1868 19998
rect 1920 19995 1976 19998
rect 2028 19995 2084 19998
rect 2136 19995 2192 19998
rect 2244 19995 2300 19998
rect 2352 19995 2408 19998
rect 2460 19995 2516 19998
rect 2568 19995 2624 19998
rect 2676 19995 2732 19998
rect 2784 19995 2840 19998
rect 2892 19995 2948 19998
rect 3000 19995 3056 19998
rect 3108 19995 3164 19998
rect 3216 19995 3272 19998
rect 3324 19995 3380 19998
rect 3432 19995 3488 19998
rect 3540 19995 3596 19998
rect 3648 19995 3704 19998
rect 3756 19995 4130 19998
rect 4182 19995 4238 19998
rect 4290 19995 4346 19998
rect 4398 19995 4454 19998
rect 4506 19995 4562 19998
rect 4614 19995 4670 19998
rect 4722 19995 4778 19998
rect 4830 19995 4886 19998
rect 4938 19995 4994 19998
rect 5046 19995 5102 19998
rect 5154 19995 5210 19998
rect 5262 19995 5318 19998
rect 5370 19995 5426 19998
rect 5478 19995 5534 19998
rect 5586 19995 5642 19998
rect 5694 19995 5750 19998
rect 5802 19995 5858 19998
rect 5910 19995 5966 19998
rect 6018 19995 6074 19998
rect 6126 19995 6836 19998
rect 6888 19995 6944 19998
rect 6996 19995 7052 19998
rect 7104 19995 7160 19998
rect 7212 19995 7268 19998
rect 7320 19995 7376 19998
rect 7428 19995 7484 19998
rect 7536 19995 7592 19998
rect 7644 19995 7700 19998
rect 7752 19995 7808 19998
rect 7860 19995 7916 19998
rect 7968 19995 8024 19998
rect 8076 19995 8132 19998
rect 8184 19995 8240 19998
rect 8292 19995 8348 19998
rect 8400 19995 8456 19998
rect 8508 19995 8564 19998
rect 8616 19995 8672 19998
rect 8724 19995 8780 19998
rect 8832 19995 9206 19998
rect 9258 19995 9314 19998
rect 9366 19995 9422 19998
rect 9474 19995 9530 19998
rect 9582 19995 9638 19998
rect 9690 19995 9746 19998
rect 9798 19995 9854 19998
rect 9906 19995 9962 19998
rect 10014 19995 10070 19998
rect 10122 19995 10178 19998
rect 10230 19995 10286 19998
rect 10338 19995 10394 19998
rect 10446 19995 10502 19998
rect 10554 19995 10610 19998
rect 10662 19995 10718 19998
rect 10770 19995 10826 19998
rect 10878 19995 10934 19998
rect 10986 19995 11042 19998
rect 11094 19995 11150 19998
rect 11202 19995 11481 19998
rect 1481 19983 11481 19995
rect 1481 19803 11481 19815
rect 1481 19751 1493 19803
rect 1545 19800 1601 19803
rect 1653 19800 3863 19803
rect 3915 19800 3971 19803
rect 4023 19800 6239 19803
rect 6291 19800 6347 19803
rect 6399 19800 6455 19803
rect 6507 19800 6563 19803
rect 6615 19800 6671 19803
rect 6723 19800 8939 19803
rect 8991 19800 9047 19803
rect 9099 19800 11309 19803
rect 11361 19800 11417 19803
rect 1545 19751 1601 19754
rect 1653 19751 3863 19754
rect 3915 19751 3971 19754
rect 4023 19751 6239 19754
rect 6291 19751 6347 19754
rect 6399 19751 6455 19754
rect 6507 19751 6563 19754
rect 6615 19751 6671 19754
rect 6723 19751 8939 19754
rect 8991 19751 9047 19754
rect 9099 19751 11309 19754
rect 11361 19751 11417 19754
rect 11469 19751 11481 19803
rect 1481 19739 11481 19751
rect 1481 19559 11481 19571
rect 1481 19556 1760 19559
rect 1812 19556 1868 19559
rect 1920 19556 1976 19559
rect 2028 19556 2084 19559
rect 2136 19556 2192 19559
rect 2244 19556 2300 19559
rect 2352 19556 2408 19559
rect 2460 19556 2516 19559
rect 2568 19556 2624 19559
rect 2676 19556 2732 19559
rect 2784 19556 2840 19559
rect 2892 19556 2948 19559
rect 3000 19556 3056 19559
rect 3108 19556 3164 19559
rect 3216 19556 3272 19559
rect 3324 19556 3380 19559
rect 3432 19556 3488 19559
rect 3540 19556 3596 19559
rect 3648 19556 3704 19559
rect 3756 19556 4130 19559
rect 4182 19556 4238 19559
rect 4290 19556 4346 19559
rect 4398 19556 4454 19559
rect 4506 19556 4562 19559
rect 4614 19556 4670 19559
rect 4722 19556 4778 19559
rect 4830 19556 4886 19559
rect 4938 19556 4994 19559
rect 5046 19556 5102 19559
rect 5154 19556 5210 19559
rect 5262 19556 5318 19559
rect 5370 19556 5426 19559
rect 5478 19556 5534 19559
rect 5586 19556 5642 19559
rect 5694 19556 5750 19559
rect 5802 19556 5858 19559
rect 5910 19556 5966 19559
rect 6018 19556 6074 19559
rect 6126 19556 6836 19559
rect 6888 19556 6944 19559
rect 6996 19556 7052 19559
rect 7104 19556 7160 19559
rect 7212 19556 7268 19559
rect 7320 19556 7376 19559
rect 7428 19556 7484 19559
rect 7536 19556 7592 19559
rect 7644 19556 7700 19559
rect 7752 19556 7808 19559
rect 7860 19556 7916 19559
rect 7968 19556 8024 19559
rect 8076 19556 8132 19559
rect 8184 19556 8240 19559
rect 8292 19556 8348 19559
rect 8400 19556 8456 19559
rect 8508 19556 8564 19559
rect 8616 19556 8672 19559
rect 8724 19556 8780 19559
rect 8832 19556 9206 19559
rect 9258 19556 9314 19559
rect 9366 19556 9422 19559
rect 9474 19556 9530 19559
rect 9582 19556 9638 19559
rect 9690 19556 9746 19559
rect 9798 19556 9854 19559
rect 9906 19556 9962 19559
rect 10014 19556 10070 19559
rect 10122 19556 10178 19559
rect 10230 19556 10286 19559
rect 10338 19556 10394 19559
rect 10446 19556 10502 19559
rect 10554 19556 10610 19559
rect 10662 19556 10718 19559
rect 10770 19556 10826 19559
rect 10878 19556 10934 19559
rect 10986 19556 11042 19559
rect 11094 19556 11150 19559
rect 11202 19556 11481 19559
rect 1481 19510 1494 19556
rect 11468 19510 11481 19556
rect 1481 19507 1760 19510
rect 1812 19507 1868 19510
rect 1920 19507 1976 19510
rect 2028 19507 2084 19510
rect 2136 19507 2192 19510
rect 2244 19507 2300 19510
rect 2352 19507 2408 19510
rect 2460 19507 2516 19510
rect 2568 19507 2624 19510
rect 2676 19507 2732 19510
rect 2784 19507 2840 19510
rect 2892 19507 2948 19510
rect 3000 19507 3056 19510
rect 3108 19507 3164 19510
rect 3216 19507 3272 19510
rect 3324 19507 3380 19510
rect 3432 19507 3488 19510
rect 3540 19507 3596 19510
rect 3648 19507 3704 19510
rect 3756 19507 4130 19510
rect 4182 19507 4238 19510
rect 4290 19507 4346 19510
rect 4398 19507 4454 19510
rect 4506 19507 4562 19510
rect 4614 19507 4670 19510
rect 4722 19507 4778 19510
rect 4830 19507 4886 19510
rect 4938 19507 4994 19510
rect 5046 19507 5102 19510
rect 5154 19507 5210 19510
rect 5262 19507 5318 19510
rect 5370 19507 5426 19510
rect 5478 19507 5534 19510
rect 5586 19507 5642 19510
rect 5694 19507 5750 19510
rect 5802 19507 5858 19510
rect 5910 19507 5966 19510
rect 6018 19507 6074 19510
rect 6126 19507 6836 19510
rect 6888 19507 6944 19510
rect 6996 19507 7052 19510
rect 7104 19507 7160 19510
rect 7212 19507 7268 19510
rect 7320 19507 7376 19510
rect 7428 19507 7484 19510
rect 7536 19507 7592 19510
rect 7644 19507 7700 19510
rect 7752 19507 7808 19510
rect 7860 19507 7916 19510
rect 7968 19507 8024 19510
rect 8076 19507 8132 19510
rect 8184 19507 8240 19510
rect 8292 19507 8348 19510
rect 8400 19507 8456 19510
rect 8508 19507 8564 19510
rect 8616 19507 8672 19510
rect 8724 19507 8780 19510
rect 8832 19507 9206 19510
rect 9258 19507 9314 19510
rect 9366 19507 9422 19510
rect 9474 19507 9530 19510
rect 9582 19507 9638 19510
rect 9690 19507 9746 19510
rect 9798 19507 9854 19510
rect 9906 19507 9962 19510
rect 10014 19507 10070 19510
rect 10122 19507 10178 19510
rect 10230 19507 10286 19510
rect 10338 19507 10394 19510
rect 10446 19507 10502 19510
rect 10554 19507 10610 19510
rect 10662 19507 10718 19510
rect 10770 19507 10826 19510
rect 10878 19507 10934 19510
rect 10986 19507 11042 19510
rect 11094 19507 11150 19510
rect 11202 19507 11481 19510
rect 1481 19495 11481 19507
rect 1481 19315 11481 19327
rect 1481 19263 1493 19315
rect 1545 19312 1601 19315
rect 1653 19312 3863 19315
rect 3915 19312 3971 19315
rect 4023 19312 6239 19315
rect 6291 19312 6347 19315
rect 6399 19312 6455 19315
rect 6507 19312 6563 19315
rect 6615 19312 6671 19315
rect 6723 19312 8939 19315
rect 8991 19312 9047 19315
rect 9099 19312 11309 19315
rect 11361 19312 11417 19315
rect 1545 19263 1601 19266
rect 1653 19263 3863 19266
rect 3915 19263 3971 19266
rect 4023 19263 6239 19266
rect 6291 19263 6347 19266
rect 6399 19263 6455 19266
rect 6507 19263 6563 19266
rect 6615 19263 6671 19266
rect 6723 19263 8939 19266
rect 8991 19263 9047 19266
rect 9099 19263 11309 19266
rect 11361 19263 11417 19266
rect 11469 19263 11481 19315
rect 1481 19251 11481 19263
rect 1213 19135 1413 19162
rect 1213 19083 1233 19135
rect 1285 19083 1341 19135
rect 1393 19083 1413 19135
rect 11549 19162 11560 23808
rect 11706 23779 11749 23808
rect 11729 23727 11749 23779
rect 11706 23671 11749 23727
rect 11729 23619 11749 23671
rect 11706 23563 11749 23619
rect 11729 23511 11749 23563
rect 11706 23455 11749 23511
rect 11729 23403 11749 23455
rect 11706 23347 11749 23403
rect 11729 23295 11749 23347
rect 11706 23239 11749 23295
rect 11729 23187 11749 23239
rect 11706 23131 11749 23187
rect 11729 23079 11749 23131
rect 11706 23023 11749 23079
rect 11729 22971 11749 23023
rect 11706 22915 11749 22971
rect 11729 22863 11749 22915
rect 11706 22807 11749 22863
rect 11729 22755 11749 22807
rect 11706 22699 11749 22755
rect 11729 22647 11749 22699
rect 11706 22591 11749 22647
rect 11729 22539 11749 22591
rect 11706 22483 11749 22539
rect 11729 22431 11749 22483
rect 11706 22375 11749 22431
rect 11729 22323 11749 22375
rect 11706 22267 11749 22323
rect 11729 22215 11749 22267
rect 11706 22159 11749 22215
rect 11729 22107 11749 22159
rect 11706 22051 11749 22107
rect 11729 21999 11749 22051
rect 11706 21943 11749 21999
rect 11729 21891 11749 21943
rect 11706 21835 11749 21891
rect 11729 21783 11749 21835
rect 11706 21727 11749 21783
rect 11729 21675 11749 21727
rect 11706 21619 11749 21675
rect 11729 21567 11749 21619
rect 11706 21511 11749 21567
rect 11729 21459 11749 21511
rect 11706 21403 11749 21459
rect 11729 21351 11749 21403
rect 11706 21295 11749 21351
rect 11729 21243 11749 21295
rect 11706 21187 11749 21243
rect 11729 21135 11749 21187
rect 11706 21079 11749 21135
rect 11729 21027 11749 21079
rect 11706 20971 11749 21027
rect 11729 20919 11749 20971
rect 11706 20863 11749 20919
rect 11729 20811 11749 20863
rect 11706 20755 11749 20811
rect 11729 20703 11749 20755
rect 11706 20647 11749 20703
rect 11729 20595 11749 20647
rect 11706 20539 11749 20595
rect 11729 20487 11749 20539
rect 11706 20431 11749 20487
rect 11729 20379 11749 20431
rect 11706 20323 11749 20379
rect 11729 20271 11749 20323
rect 11706 20215 11749 20271
rect 11729 20163 11749 20215
rect 11706 20107 11749 20163
rect 11729 20055 11749 20107
rect 11706 19999 11749 20055
rect 11729 19947 11749 19999
rect 11706 19891 11749 19947
rect 11729 19839 11749 19891
rect 11706 19783 11749 19839
rect 11729 19731 11749 19783
rect 11706 19675 11749 19731
rect 11729 19623 11749 19675
rect 11706 19567 11749 19623
rect 11729 19515 11749 19567
rect 11706 19459 11749 19515
rect 11729 19407 11749 19459
rect 11706 19351 11749 19407
rect 11729 19299 11749 19351
rect 11706 19243 11749 19299
rect 11729 19191 11749 19243
rect 11706 19162 11749 19191
rect 11549 19135 11749 19162
rect 11549 19083 11569 19135
rect 11621 19083 11677 19135
rect 11729 19083 11749 19135
rect 1213 18920 1413 19083
rect 1481 19071 11481 19083
rect 1481 19068 1760 19071
rect 1812 19068 1868 19071
rect 1920 19068 1976 19071
rect 2028 19068 2084 19071
rect 2136 19068 2192 19071
rect 2244 19068 2300 19071
rect 2352 19068 2408 19071
rect 2460 19068 2516 19071
rect 2568 19068 2624 19071
rect 2676 19068 2732 19071
rect 2784 19068 2840 19071
rect 2892 19068 2948 19071
rect 3000 19068 3056 19071
rect 3108 19068 3164 19071
rect 3216 19068 3272 19071
rect 3324 19068 3380 19071
rect 3432 19068 3488 19071
rect 3540 19068 3596 19071
rect 3648 19068 3704 19071
rect 3756 19068 4130 19071
rect 4182 19068 4238 19071
rect 4290 19068 4346 19071
rect 4398 19068 4454 19071
rect 4506 19068 4562 19071
rect 4614 19068 4670 19071
rect 4722 19068 4778 19071
rect 4830 19068 4886 19071
rect 4938 19068 4994 19071
rect 5046 19068 5102 19071
rect 5154 19068 5210 19071
rect 5262 19068 5318 19071
rect 5370 19068 5426 19071
rect 5478 19068 5534 19071
rect 5586 19068 5642 19071
rect 5694 19068 5750 19071
rect 5802 19068 5858 19071
rect 5910 19068 5966 19071
rect 6018 19068 6074 19071
rect 6126 19068 6836 19071
rect 6888 19068 6944 19071
rect 6996 19068 7052 19071
rect 7104 19068 7160 19071
rect 7212 19068 7268 19071
rect 7320 19068 7376 19071
rect 7428 19068 7484 19071
rect 7536 19068 7592 19071
rect 7644 19068 7700 19071
rect 7752 19068 7808 19071
rect 7860 19068 7916 19071
rect 7968 19068 8024 19071
rect 8076 19068 8132 19071
rect 8184 19068 8240 19071
rect 8292 19068 8348 19071
rect 8400 19068 8456 19071
rect 8508 19068 8564 19071
rect 8616 19068 8672 19071
rect 8724 19068 8780 19071
rect 8832 19068 9206 19071
rect 9258 19068 9314 19071
rect 9366 19068 9422 19071
rect 9474 19068 9530 19071
rect 9582 19068 9638 19071
rect 9690 19068 9746 19071
rect 9798 19068 9854 19071
rect 9906 19068 9962 19071
rect 10014 19068 10070 19071
rect 10122 19068 10178 19071
rect 10230 19068 10286 19071
rect 10338 19068 10394 19071
rect 10446 19068 10502 19071
rect 10554 19068 10610 19071
rect 10662 19068 10718 19071
rect 10770 19068 10826 19071
rect 10878 19068 10934 19071
rect 10986 19068 11042 19071
rect 11094 19068 11150 19071
rect 11202 19068 11481 19071
rect 1481 19022 1494 19068
rect 11468 19022 11481 19068
rect 1481 19019 1760 19022
rect 1812 19019 1868 19022
rect 1920 19019 1976 19022
rect 2028 19019 2084 19022
rect 2136 19019 2192 19022
rect 2244 19019 2300 19022
rect 2352 19019 2408 19022
rect 2460 19019 2516 19022
rect 2568 19019 2624 19022
rect 2676 19019 2732 19022
rect 2784 19019 2840 19022
rect 2892 19019 2948 19022
rect 3000 19019 3056 19022
rect 3108 19019 3164 19022
rect 3216 19019 3272 19022
rect 3324 19019 3380 19022
rect 3432 19019 3488 19022
rect 3540 19019 3596 19022
rect 3648 19019 3704 19022
rect 3756 19019 4130 19022
rect 4182 19019 4238 19022
rect 4290 19019 4346 19022
rect 4398 19019 4454 19022
rect 4506 19019 4562 19022
rect 4614 19019 4670 19022
rect 4722 19019 4778 19022
rect 4830 19019 4886 19022
rect 4938 19019 4994 19022
rect 5046 19019 5102 19022
rect 5154 19019 5210 19022
rect 5262 19019 5318 19022
rect 5370 19019 5426 19022
rect 5478 19019 5534 19022
rect 5586 19019 5642 19022
rect 5694 19019 5750 19022
rect 5802 19019 5858 19022
rect 5910 19019 5966 19022
rect 6018 19019 6074 19022
rect 6126 19019 6836 19022
rect 6888 19019 6944 19022
rect 6996 19019 7052 19022
rect 7104 19019 7160 19022
rect 7212 19019 7268 19022
rect 7320 19019 7376 19022
rect 7428 19019 7484 19022
rect 7536 19019 7592 19022
rect 7644 19019 7700 19022
rect 7752 19019 7808 19022
rect 7860 19019 7916 19022
rect 7968 19019 8024 19022
rect 8076 19019 8132 19022
rect 8184 19019 8240 19022
rect 8292 19019 8348 19022
rect 8400 19019 8456 19022
rect 8508 19019 8564 19022
rect 8616 19019 8672 19022
rect 8724 19019 8780 19022
rect 8832 19019 9206 19022
rect 9258 19019 9314 19022
rect 9366 19019 9422 19022
rect 9474 19019 9530 19022
rect 9582 19019 9638 19022
rect 9690 19019 9746 19022
rect 9798 19019 9854 19022
rect 9906 19019 9962 19022
rect 10014 19019 10070 19022
rect 10122 19019 10178 19022
rect 10230 19019 10286 19022
rect 10338 19019 10394 19022
rect 10446 19019 10502 19022
rect 10554 19019 10610 19022
rect 10662 19019 10718 19022
rect 10770 19019 10826 19022
rect 10878 19019 10934 19022
rect 10986 19019 11042 19022
rect 11094 19019 11150 19022
rect 11202 19019 11481 19022
rect 1481 19007 11481 19019
rect 11549 18920 11749 19083
rect 1213 18720 11749 18920
rect 12001 18641 12012 24343
rect 950 18629 12012 18641
rect 950 18622 1760 18629
rect 1812 18622 1868 18629
rect 1920 18622 1976 18629
rect 2028 18622 2084 18629
rect 2136 18622 2192 18629
rect 2244 18622 2300 18629
rect 2352 18622 2408 18629
rect 2460 18622 2516 18629
rect 2568 18622 2624 18629
rect 2676 18622 2732 18629
rect 2784 18622 2840 18629
rect 2892 18622 2948 18629
rect 3000 18622 3056 18629
rect 3108 18622 3164 18629
rect 3216 18622 3272 18629
rect 3324 18622 3380 18629
rect 3432 18622 3488 18629
rect 3540 18622 3596 18629
rect 3648 18622 3704 18629
rect 3756 18622 4130 18629
rect 4182 18622 4238 18629
rect 4290 18622 4346 18629
rect 4398 18622 4454 18629
rect 4506 18622 4562 18629
rect 4614 18622 4670 18629
rect 4722 18622 4778 18629
rect 4830 18622 4886 18629
rect 4938 18622 4994 18629
rect 5046 18622 5102 18629
rect 5154 18622 5210 18629
rect 5262 18622 5318 18629
rect 5370 18622 5426 18629
rect 5478 18622 5534 18629
rect 5586 18622 5642 18629
rect 5694 18622 5750 18629
rect 5802 18622 5858 18629
rect 5910 18622 5966 18629
rect 6018 18622 6074 18629
rect 6126 18622 6836 18629
rect 6888 18622 6944 18629
rect 6996 18622 7052 18629
rect 7104 18622 7160 18629
rect 7212 18622 7268 18629
rect 7320 18622 7376 18629
rect 7428 18622 7484 18629
rect 7536 18622 7592 18629
rect 7644 18622 7700 18629
rect 7752 18622 7808 18629
rect 7860 18622 7916 18629
rect 7968 18622 8024 18629
rect 8076 18622 8132 18629
rect 8184 18622 8240 18629
rect 8292 18622 8348 18629
rect 8400 18622 8456 18629
rect 8508 18622 8564 18629
rect 8616 18622 8672 18629
rect 8724 18622 8780 18629
rect 8832 18622 9206 18629
rect 9258 18622 9314 18629
rect 9366 18622 9422 18629
rect 9474 18622 9530 18629
rect 9582 18622 9638 18629
rect 9690 18622 9746 18629
rect 9798 18622 9854 18629
rect 9906 18622 9962 18629
rect 10014 18622 10070 18629
rect 10122 18622 10178 18629
rect 10230 18622 10286 18629
rect 10338 18622 10394 18629
rect 10446 18622 10502 18629
rect 10554 18622 10610 18629
rect 10662 18622 10718 18629
rect 10770 18622 10826 18629
rect 10878 18622 10934 18629
rect 10986 18622 11042 18629
rect 11094 18622 11150 18629
rect 11202 18622 12012 18629
rect 950 18476 1058 18622
rect 11904 18476 12012 18622
rect 950 18469 1760 18476
rect 1812 18469 1868 18476
rect 1920 18469 1976 18476
rect 2028 18469 2084 18476
rect 2136 18469 2192 18476
rect 2244 18469 2300 18476
rect 2352 18469 2408 18476
rect 2460 18469 2516 18476
rect 2568 18469 2624 18476
rect 2676 18469 2732 18476
rect 2784 18469 2840 18476
rect 2892 18469 2948 18476
rect 3000 18469 3056 18476
rect 3108 18469 3164 18476
rect 3216 18469 3272 18476
rect 3324 18469 3380 18476
rect 3432 18469 3488 18476
rect 3540 18469 3596 18476
rect 3648 18469 3704 18476
rect 3756 18469 4130 18476
rect 4182 18469 4238 18476
rect 4290 18469 4346 18476
rect 4398 18469 4454 18476
rect 4506 18469 4562 18476
rect 4614 18469 4670 18476
rect 4722 18469 4778 18476
rect 4830 18469 4886 18476
rect 4938 18469 4994 18476
rect 5046 18469 5102 18476
rect 5154 18469 5210 18476
rect 5262 18469 5318 18476
rect 5370 18469 5426 18476
rect 5478 18469 5534 18476
rect 5586 18469 5642 18476
rect 5694 18469 5750 18476
rect 5802 18469 5858 18476
rect 5910 18469 5966 18476
rect 6018 18469 6074 18476
rect 6126 18469 6836 18476
rect 6888 18469 6944 18476
rect 6996 18469 7052 18476
rect 7104 18469 7160 18476
rect 7212 18469 7268 18476
rect 7320 18469 7376 18476
rect 7428 18469 7484 18476
rect 7536 18469 7592 18476
rect 7644 18469 7700 18476
rect 7752 18469 7808 18476
rect 7860 18469 7916 18476
rect 7968 18469 8024 18476
rect 8076 18469 8132 18476
rect 8184 18469 8240 18476
rect 8292 18469 8348 18476
rect 8400 18469 8456 18476
rect 8508 18469 8564 18476
rect 8616 18469 8672 18476
rect 8724 18469 8780 18476
rect 8832 18469 9206 18476
rect 9258 18469 9314 18476
rect 9366 18469 9422 18476
rect 9474 18469 9530 18476
rect 9582 18469 9638 18476
rect 9690 18469 9746 18476
rect 9798 18469 9854 18476
rect 9906 18469 9962 18476
rect 10014 18469 10070 18476
rect 10122 18469 10178 18476
rect 10230 18469 10286 18476
rect 10338 18469 10394 18476
rect 10446 18469 10502 18476
rect 10554 18469 10610 18476
rect 10662 18469 10718 18476
rect 10770 18469 10826 18476
rect 10878 18469 10934 18476
rect 10986 18469 11042 18476
rect 11094 18469 11150 18476
rect 11202 18469 12012 18476
rect 950 18457 12012 18469
rect 950 12769 961 18457
rect 1213 18178 11749 18378
rect 1213 18015 1413 18178
rect 1481 18079 11481 18091
rect 1481 18076 1760 18079
rect 1812 18076 1868 18079
rect 1920 18076 1976 18079
rect 2028 18076 2084 18079
rect 2136 18076 2192 18079
rect 2244 18076 2300 18079
rect 2352 18076 2408 18079
rect 2460 18076 2516 18079
rect 2568 18076 2624 18079
rect 2676 18076 2732 18079
rect 2784 18076 2840 18079
rect 2892 18076 2948 18079
rect 3000 18076 3056 18079
rect 3108 18076 3164 18079
rect 3216 18076 3272 18079
rect 3324 18076 3380 18079
rect 3432 18076 3488 18079
rect 3540 18076 3596 18079
rect 3648 18076 3704 18079
rect 3756 18076 4130 18079
rect 4182 18076 4238 18079
rect 4290 18076 4346 18079
rect 4398 18076 4454 18079
rect 4506 18076 4562 18079
rect 4614 18076 4670 18079
rect 4722 18076 4778 18079
rect 4830 18076 4886 18079
rect 4938 18076 4994 18079
rect 5046 18076 5102 18079
rect 5154 18076 5210 18079
rect 5262 18076 5318 18079
rect 5370 18076 5426 18079
rect 5478 18076 5534 18079
rect 5586 18076 5642 18079
rect 5694 18076 5750 18079
rect 5802 18076 5858 18079
rect 5910 18076 5966 18079
rect 6018 18076 6074 18079
rect 6126 18076 6836 18079
rect 6888 18076 6944 18079
rect 6996 18076 7052 18079
rect 7104 18076 7160 18079
rect 7212 18076 7268 18079
rect 7320 18076 7376 18079
rect 7428 18076 7484 18079
rect 7536 18076 7592 18079
rect 7644 18076 7700 18079
rect 7752 18076 7808 18079
rect 7860 18076 7916 18079
rect 7968 18076 8024 18079
rect 8076 18076 8132 18079
rect 8184 18076 8240 18079
rect 8292 18076 8348 18079
rect 8400 18076 8456 18079
rect 8508 18076 8564 18079
rect 8616 18076 8672 18079
rect 8724 18076 8780 18079
rect 8832 18076 9206 18079
rect 9258 18076 9314 18079
rect 9366 18076 9422 18079
rect 9474 18076 9530 18079
rect 9582 18076 9638 18079
rect 9690 18076 9746 18079
rect 9798 18076 9854 18079
rect 9906 18076 9962 18079
rect 10014 18076 10070 18079
rect 10122 18076 10178 18079
rect 10230 18076 10286 18079
rect 10338 18076 10394 18079
rect 10446 18076 10502 18079
rect 10554 18076 10610 18079
rect 10662 18076 10718 18079
rect 10770 18076 10826 18079
rect 10878 18076 10934 18079
rect 10986 18076 11042 18079
rect 11094 18076 11150 18079
rect 11202 18076 11481 18079
rect 1481 18030 1494 18076
rect 11468 18030 11481 18076
rect 1481 18027 1760 18030
rect 1812 18027 1868 18030
rect 1920 18027 1976 18030
rect 2028 18027 2084 18030
rect 2136 18027 2192 18030
rect 2244 18027 2300 18030
rect 2352 18027 2408 18030
rect 2460 18027 2516 18030
rect 2568 18027 2624 18030
rect 2676 18027 2732 18030
rect 2784 18027 2840 18030
rect 2892 18027 2948 18030
rect 3000 18027 3056 18030
rect 3108 18027 3164 18030
rect 3216 18027 3272 18030
rect 3324 18027 3380 18030
rect 3432 18027 3488 18030
rect 3540 18027 3596 18030
rect 3648 18027 3704 18030
rect 3756 18027 4130 18030
rect 4182 18027 4238 18030
rect 4290 18027 4346 18030
rect 4398 18027 4454 18030
rect 4506 18027 4562 18030
rect 4614 18027 4670 18030
rect 4722 18027 4778 18030
rect 4830 18027 4886 18030
rect 4938 18027 4994 18030
rect 5046 18027 5102 18030
rect 5154 18027 5210 18030
rect 5262 18027 5318 18030
rect 5370 18027 5426 18030
rect 5478 18027 5534 18030
rect 5586 18027 5642 18030
rect 5694 18027 5750 18030
rect 5802 18027 5858 18030
rect 5910 18027 5966 18030
rect 6018 18027 6074 18030
rect 6126 18027 6836 18030
rect 6888 18027 6944 18030
rect 6996 18027 7052 18030
rect 7104 18027 7160 18030
rect 7212 18027 7268 18030
rect 7320 18027 7376 18030
rect 7428 18027 7484 18030
rect 7536 18027 7592 18030
rect 7644 18027 7700 18030
rect 7752 18027 7808 18030
rect 7860 18027 7916 18030
rect 7968 18027 8024 18030
rect 8076 18027 8132 18030
rect 8184 18027 8240 18030
rect 8292 18027 8348 18030
rect 8400 18027 8456 18030
rect 8508 18027 8564 18030
rect 8616 18027 8672 18030
rect 8724 18027 8780 18030
rect 8832 18027 9206 18030
rect 9258 18027 9314 18030
rect 9366 18027 9422 18030
rect 9474 18027 9530 18030
rect 9582 18027 9638 18030
rect 9690 18027 9746 18030
rect 9798 18027 9854 18030
rect 9906 18027 9962 18030
rect 10014 18027 10070 18030
rect 10122 18027 10178 18030
rect 10230 18027 10286 18030
rect 10338 18027 10394 18030
rect 10446 18027 10502 18030
rect 10554 18027 10610 18030
rect 10662 18027 10718 18030
rect 10770 18027 10826 18030
rect 10878 18027 10934 18030
rect 10986 18027 11042 18030
rect 11094 18027 11150 18030
rect 11202 18027 11481 18030
rect 1481 18015 11481 18027
rect 11549 18015 11749 18178
rect 1213 17963 1233 18015
rect 1285 17963 1341 18015
rect 1393 17963 1413 18015
rect 1213 17936 1413 17963
rect 1213 17907 1256 17936
rect 1213 17855 1233 17907
rect 1213 17799 1256 17855
rect 1213 17747 1233 17799
rect 1213 17691 1256 17747
rect 1213 17639 1233 17691
rect 1213 17583 1256 17639
rect 1213 17531 1233 17583
rect 1213 17475 1256 17531
rect 1213 17423 1233 17475
rect 1213 17367 1256 17423
rect 1213 17315 1233 17367
rect 1213 17259 1256 17315
rect 1213 17207 1233 17259
rect 1213 17151 1256 17207
rect 1213 17099 1233 17151
rect 1213 17043 1256 17099
rect 1213 16991 1233 17043
rect 1213 16935 1256 16991
rect 1213 16883 1233 16935
rect 1213 16827 1256 16883
rect 1213 16775 1233 16827
rect 1213 16719 1256 16775
rect 1213 16667 1233 16719
rect 1213 16611 1256 16667
rect 1213 16559 1233 16611
rect 1213 16503 1256 16559
rect 1213 16451 1233 16503
rect 1213 16395 1256 16451
rect 1213 16343 1233 16395
rect 1213 16287 1256 16343
rect 1213 16235 1233 16287
rect 1213 16179 1256 16235
rect 1213 16127 1233 16179
rect 1213 16071 1256 16127
rect 1213 16019 1233 16071
rect 1213 15963 1256 16019
rect 1213 15911 1233 15963
rect 1213 15855 1256 15911
rect 1213 15803 1233 15855
rect 1213 15747 1256 15803
rect 1213 15695 1233 15747
rect 1213 15639 1256 15695
rect 1213 15587 1233 15639
rect 1213 15531 1256 15587
rect 1213 15479 1233 15531
rect 1213 15423 1256 15479
rect 1213 15371 1233 15423
rect 1213 15315 1256 15371
rect 1213 15263 1233 15315
rect 1213 15207 1256 15263
rect 1213 15155 1233 15207
rect 1213 15099 1256 15155
rect 1213 15047 1233 15099
rect 1213 14991 1256 15047
rect 1213 14939 1233 14991
rect 1213 14883 1256 14939
rect 1213 14831 1233 14883
rect 1213 14775 1256 14831
rect 1213 14723 1233 14775
rect 1213 14667 1256 14723
rect 1213 14615 1233 14667
rect 1213 14559 1256 14615
rect 1213 14507 1233 14559
rect 1213 14451 1256 14507
rect 1213 14399 1233 14451
rect 1213 14343 1256 14399
rect 1213 14291 1233 14343
rect 1213 14235 1256 14291
rect 1213 14183 1233 14235
rect 1213 14127 1256 14183
rect 1213 14075 1233 14127
rect 1213 14019 1256 14075
rect 1213 13967 1233 14019
rect 1213 13911 1256 13967
rect 1213 13859 1233 13911
rect 1213 13803 1256 13859
rect 1213 13751 1233 13803
rect 1213 13695 1256 13751
rect 1213 13643 1233 13695
rect 1213 13587 1256 13643
rect 1213 13535 1233 13587
rect 1213 13479 1256 13535
rect 1213 13427 1233 13479
rect 1213 13371 1256 13427
rect 1213 13319 1233 13371
rect 1213 13290 1256 13319
rect 1402 13290 1413 17936
rect 11549 17963 11569 18015
rect 11621 17963 11677 18015
rect 11729 17963 11749 18015
rect 11549 17936 11749 17963
rect 1481 17835 11481 17847
rect 1481 17783 1493 17835
rect 1545 17832 1601 17835
rect 1653 17832 3863 17835
rect 3915 17832 3971 17835
rect 4023 17832 6239 17835
rect 6291 17832 6347 17835
rect 6399 17832 6455 17835
rect 6507 17832 6563 17835
rect 6615 17832 6671 17835
rect 6723 17832 8939 17835
rect 8991 17832 9047 17835
rect 9099 17832 11309 17835
rect 11361 17832 11417 17835
rect 1545 17783 1601 17786
rect 1653 17783 3863 17786
rect 3915 17783 3971 17786
rect 4023 17783 6239 17786
rect 6291 17783 6347 17786
rect 6399 17783 6455 17786
rect 6507 17783 6563 17786
rect 6615 17783 6671 17786
rect 6723 17783 8939 17786
rect 8991 17783 9047 17786
rect 9099 17783 11309 17786
rect 11361 17783 11417 17786
rect 11469 17783 11481 17835
rect 1481 17771 11481 17783
rect 1481 17591 11481 17603
rect 1481 17588 1760 17591
rect 1812 17588 1868 17591
rect 1920 17588 1976 17591
rect 2028 17588 2084 17591
rect 2136 17588 2192 17591
rect 2244 17588 2300 17591
rect 2352 17588 2408 17591
rect 2460 17588 2516 17591
rect 2568 17588 2624 17591
rect 2676 17588 2732 17591
rect 2784 17588 2840 17591
rect 2892 17588 2948 17591
rect 3000 17588 3056 17591
rect 3108 17588 3164 17591
rect 3216 17588 3272 17591
rect 3324 17588 3380 17591
rect 3432 17588 3488 17591
rect 3540 17588 3596 17591
rect 3648 17588 3704 17591
rect 3756 17588 4130 17591
rect 4182 17588 4238 17591
rect 4290 17588 4346 17591
rect 4398 17588 4454 17591
rect 4506 17588 4562 17591
rect 4614 17588 4670 17591
rect 4722 17588 4778 17591
rect 4830 17588 4886 17591
rect 4938 17588 4994 17591
rect 5046 17588 5102 17591
rect 5154 17588 5210 17591
rect 5262 17588 5318 17591
rect 5370 17588 5426 17591
rect 5478 17588 5534 17591
rect 5586 17588 5642 17591
rect 5694 17588 5750 17591
rect 5802 17588 5858 17591
rect 5910 17588 5966 17591
rect 6018 17588 6074 17591
rect 6126 17588 6836 17591
rect 6888 17588 6944 17591
rect 6996 17588 7052 17591
rect 7104 17588 7160 17591
rect 7212 17588 7268 17591
rect 7320 17588 7376 17591
rect 7428 17588 7484 17591
rect 7536 17588 7592 17591
rect 7644 17588 7700 17591
rect 7752 17588 7808 17591
rect 7860 17588 7916 17591
rect 7968 17588 8024 17591
rect 8076 17588 8132 17591
rect 8184 17588 8240 17591
rect 8292 17588 8348 17591
rect 8400 17588 8456 17591
rect 8508 17588 8564 17591
rect 8616 17588 8672 17591
rect 8724 17588 8780 17591
rect 8832 17588 9206 17591
rect 9258 17588 9314 17591
rect 9366 17588 9422 17591
rect 9474 17588 9530 17591
rect 9582 17588 9638 17591
rect 9690 17588 9746 17591
rect 9798 17588 9854 17591
rect 9906 17588 9962 17591
rect 10014 17588 10070 17591
rect 10122 17588 10178 17591
rect 10230 17588 10286 17591
rect 10338 17588 10394 17591
rect 10446 17588 10502 17591
rect 10554 17588 10610 17591
rect 10662 17588 10718 17591
rect 10770 17588 10826 17591
rect 10878 17588 10934 17591
rect 10986 17588 11042 17591
rect 11094 17588 11150 17591
rect 11202 17588 11481 17591
rect 1481 17542 1494 17588
rect 11468 17542 11481 17588
rect 1481 17539 1760 17542
rect 1812 17539 1868 17542
rect 1920 17539 1976 17542
rect 2028 17539 2084 17542
rect 2136 17539 2192 17542
rect 2244 17539 2300 17542
rect 2352 17539 2408 17542
rect 2460 17539 2516 17542
rect 2568 17539 2624 17542
rect 2676 17539 2732 17542
rect 2784 17539 2840 17542
rect 2892 17539 2948 17542
rect 3000 17539 3056 17542
rect 3108 17539 3164 17542
rect 3216 17539 3272 17542
rect 3324 17539 3380 17542
rect 3432 17539 3488 17542
rect 3540 17539 3596 17542
rect 3648 17539 3704 17542
rect 3756 17539 4130 17542
rect 4182 17539 4238 17542
rect 4290 17539 4346 17542
rect 4398 17539 4454 17542
rect 4506 17539 4562 17542
rect 4614 17539 4670 17542
rect 4722 17539 4778 17542
rect 4830 17539 4886 17542
rect 4938 17539 4994 17542
rect 5046 17539 5102 17542
rect 5154 17539 5210 17542
rect 5262 17539 5318 17542
rect 5370 17539 5426 17542
rect 5478 17539 5534 17542
rect 5586 17539 5642 17542
rect 5694 17539 5750 17542
rect 5802 17539 5858 17542
rect 5910 17539 5966 17542
rect 6018 17539 6074 17542
rect 6126 17539 6836 17542
rect 6888 17539 6944 17542
rect 6996 17539 7052 17542
rect 7104 17539 7160 17542
rect 7212 17539 7268 17542
rect 7320 17539 7376 17542
rect 7428 17539 7484 17542
rect 7536 17539 7592 17542
rect 7644 17539 7700 17542
rect 7752 17539 7808 17542
rect 7860 17539 7916 17542
rect 7968 17539 8024 17542
rect 8076 17539 8132 17542
rect 8184 17539 8240 17542
rect 8292 17539 8348 17542
rect 8400 17539 8456 17542
rect 8508 17539 8564 17542
rect 8616 17539 8672 17542
rect 8724 17539 8780 17542
rect 8832 17539 9206 17542
rect 9258 17539 9314 17542
rect 9366 17539 9422 17542
rect 9474 17539 9530 17542
rect 9582 17539 9638 17542
rect 9690 17539 9746 17542
rect 9798 17539 9854 17542
rect 9906 17539 9962 17542
rect 10014 17539 10070 17542
rect 10122 17539 10178 17542
rect 10230 17539 10286 17542
rect 10338 17539 10394 17542
rect 10446 17539 10502 17542
rect 10554 17539 10610 17542
rect 10662 17539 10718 17542
rect 10770 17539 10826 17542
rect 10878 17539 10934 17542
rect 10986 17539 11042 17542
rect 11094 17539 11150 17542
rect 11202 17539 11481 17542
rect 1481 17527 11481 17539
rect 1481 17347 11481 17359
rect 1481 17295 1493 17347
rect 1545 17344 1601 17347
rect 1653 17344 3863 17347
rect 3915 17344 3971 17347
rect 4023 17344 6239 17347
rect 6291 17344 6347 17347
rect 6399 17344 6455 17347
rect 6507 17344 6563 17347
rect 6615 17344 6671 17347
rect 6723 17344 8939 17347
rect 8991 17344 9047 17347
rect 9099 17344 11309 17347
rect 11361 17344 11417 17347
rect 1545 17295 1601 17298
rect 1653 17295 3863 17298
rect 3915 17295 3971 17298
rect 4023 17295 6239 17298
rect 6291 17295 6347 17298
rect 6399 17295 6455 17298
rect 6507 17295 6563 17298
rect 6615 17295 6671 17298
rect 6723 17295 8939 17298
rect 8991 17295 9047 17298
rect 9099 17295 11309 17298
rect 11361 17295 11417 17298
rect 11469 17295 11481 17347
rect 1481 17283 11481 17295
rect 1481 17103 11481 17115
rect 1481 17100 1760 17103
rect 1812 17100 1868 17103
rect 1920 17100 1976 17103
rect 2028 17100 2084 17103
rect 2136 17100 2192 17103
rect 2244 17100 2300 17103
rect 2352 17100 2408 17103
rect 2460 17100 2516 17103
rect 2568 17100 2624 17103
rect 2676 17100 2732 17103
rect 2784 17100 2840 17103
rect 2892 17100 2948 17103
rect 3000 17100 3056 17103
rect 3108 17100 3164 17103
rect 3216 17100 3272 17103
rect 3324 17100 3380 17103
rect 3432 17100 3488 17103
rect 3540 17100 3596 17103
rect 3648 17100 3704 17103
rect 3756 17100 4130 17103
rect 4182 17100 4238 17103
rect 4290 17100 4346 17103
rect 4398 17100 4454 17103
rect 4506 17100 4562 17103
rect 4614 17100 4670 17103
rect 4722 17100 4778 17103
rect 4830 17100 4886 17103
rect 4938 17100 4994 17103
rect 5046 17100 5102 17103
rect 5154 17100 5210 17103
rect 5262 17100 5318 17103
rect 5370 17100 5426 17103
rect 5478 17100 5534 17103
rect 5586 17100 5642 17103
rect 5694 17100 5750 17103
rect 5802 17100 5858 17103
rect 5910 17100 5966 17103
rect 6018 17100 6074 17103
rect 6126 17100 6836 17103
rect 6888 17100 6944 17103
rect 6996 17100 7052 17103
rect 7104 17100 7160 17103
rect 7212 17100 7268 17103
rect 7320 17100 7376 17103
rect 7428 17100 7484 17103
rect 7536 17100 7592 17103
rect 7644 17100 7700 17103
rect 7752 17100 7808 17103
rect 7860 17100 7916 17103
rect 7968 17100 8024 17103
rect 8076 17100 8132 17103
rect 8184 17100 8240 17103
rect 8292 17100 8348 17103
rect 8400 17100 8456 17103
rect 8508 17100 8564 17103
rect 8616 17100 8672 17103
rect 8724 17100 8780 17103
rect 8832 17100 9206 17103
rect 9258 17100 9314 17103
rect 9366 17100 9422 17103
rect 9474 17100 9530 17103
rect 9582 17100 9638 17103
rect 9690 17100 9746 17103
rect 9798 17100 9854 17103
rect 9906 17100 9962 17103
rect 10014 17100 10070 17103
rect 10122 17100 10178 17103
rect 10230 17100 10286 17103
rect 10338 17100 10394 17103
rect 10446 17100 10502 17103
rect 10554 17100 10610 17103
rect 10662 17100 10718 17103
rect 10770 17100 10826 17103
rect 10878 17100 10934 17103
rect 10986 17100 11042 17103
rect 11094 17100 11150 17103
rect 11202 17100 11481 17103
rect 1481 17054 1494 17100
rect 11468 17054 11481 17100
rect 1481 17051 1760 17054
rect 1812 17051 1868 17054
rect 1920 17051 1976 17054
rect 2028 17051 2084 17054
rect 2136 17051 2192 17054
rect 2244 17051 2300 17054
rect 2352 17051 2408 17054
rect 2460 17051 2516 17054
rect 2568 17051 2624 17054
rect 2676 17051 2732 17054
rect 2784 17051 2840 17054
rect 2892 17051 2948 17054
rect 3000 17051 3056 17054
rect 3108 17051 3164 17054
rect 3216 17051 3272 17054
rect 3324 17051 3380 17054
rect 3432 17051 3488 17054
rect 3540 17051 3596 17054
rect 3648 17051 3704 17054
rect 3756 17051 4130 17054
rect 4182 17051 4238 17054
rect 4290 17051 4346 17054
rect 4398 17051 4454 17054
rect 4506 17051 4562 17054
rect 4614 17051 4670 17054
rect 4722 17051 4778 17054
rect 4830 17051 4886 17054
rect 4938 17051 4994 17054
rect 5046 17051 5102 17054
rect 5154 17051 5210 17054
rect 5262 17051 5318 17054
rect 5370 17051 5426 17054
rect 5478 17051 5534 17054
rect 5586 17051 5642 17054
rect 5694 17051 5750 17054
rect 5802 17051 5858 17054
rect 5910 17051 5966 17054
rect 6018 17051 6074 17054
rect 6126 17051 6836 17054
rect 6888 17051 6944 17054
rect 6996 17051 7052 17054
rect 7104 17051 7160 17054
rect 7212 17051 7268 17054
rect 7320 17051 7376 17054
rect 7428 17051 7484 17054
rect 7536 17051 7592 17054
rect 7644 17051 7700 17054
rect 7752 17051 7808 17054
rect 7860 17051 7916 17054
rect 7968 17051 8024 17054
rect 8076 17051 8132 17054
rect 8184 17051 8240 17054
rect 8292 17051 8348 17054
rect 8400 17051 8456 17054
rect 8508 17051 8564 17054
rect 8616 17051 8672 17054
rect 8724 17051 8780 17054
rect 8832 17051 9206 17054
rect 9258 17051 9314 17054
rect 9366 17051 9422 17054
rect 9474 17051 9530 17054
rect 9582 17051 9638 17054
rect 9690 17051 9746 17054
rect 9798 17051 9854 17054
rect 9906 17051 9962 17054
rect 10014 17051 10070 17054
rect 10122 17051 10178 17054
rect 10230 17051 10286 17054
rect 10338 17051 10394 17054
rect 10446 17051 10502 17054
rect 10554 17051 10610 17054
rect 10662 17051 10718 17054
rect 10770 17051 10826 17054
rect 10878 17051 10934 17054
rect 10986 17051 11042 17054
rect 11094 17051 11150 17054
rect 11202 17051 11481 17054
rect 1481 17039 11481 17051
rect 1481 16859 11481 16871
rect 1481 16807 1493 16859
rect 1545 16856 1601 16859
rect 1653 16856 3863 16859
rect 3915 16856 3971 16859
rect 4023 16856 6239 16859
rect 6291 16856 6347 16859
rect 6399 16856 6455 16859
rect 6507 16856 6563 16859
rect 6615 16856 6671 16859
rect 6723 16856 8939 16859
rect 8991 16856 9047 16859
rect 9099 16856 11309 16859
rect 11361 16856 11417 16859
rect 1545 16807 1601 16810
rect 1653 16807 3863 16810
rect 3915 16807 3971 16810
rect 4023 16807 6239 16810
rect 6291 16807 6347 16810
rect 6399 16807 6455 16810
rect 6507 16807 6563 16810
rect 6615 16807 6671 16810
rect 6723 16807 8939 16810
rect 8991 16807 9047 16810
rect 9099 16807 11309 16810
rect 11361 16807 11417 16810
rect 11469 16807 11481 16859
rect 1481 16795 11481 16807
rect 1481 16615 11481 16627
rect 1481 16612 1760 16615
rect 1812 16612 1868 16615
rect 1920 16612 1976 16615
rect 2028 16612 2084 16615
rect 2136 16612 2192 16615
rect 2244 16612 2300 16615
rect 2352 16612 2408 16615
rect 2460 16612 2516 16615
rect 2568 16612 2624 16615
rect 2676 16612 2732 16615
rect 2784 16612 2840 16615
rect 2892 16612 2948 16615
rect 3000 16612 3056 16615
rect 3108 16612 3164 16615
rect 3216 16612 3272 16615
rect 3324 16612 3380 16615
rect 3432 16612 3488 16615
rect 3540 16612 3596 16615
rect 3648 16612 3704 16615
rect 3756 16612 4130 16615
rect 4182 16612 4238 16615
rect 4290 16612 4346 16615
rect 4398 16612 4454 16615
rect 4506 16612 4562 16615
rect 4614 16612 4670 16615
rect 4722 16612 4778 16615
rect 4830 16612 4886 16615
rect 4938 16612 4994 16615
rect 5046 16612 5102 16615
rect 5154 16612 5210 16615
rect 5262 16612 5318 16615
rect 5370 16612 5426 16615
rect 5478 16612 5534 16615
rect 5586 16612 5642 16615
rect 5694 16612 5750 16615
rect 5802 16612 5858 16615
rect 5910 16612 5966 16615
rect 6018 16612 6074 16615
rect 6126 16612 6836 16615
rect 6888 16612 6944 16615
rect 6996 16612 7052 16615
rect 7104 16612 7160 16615
rect 7212 16612 7268 16615
rect 7320 16612 7376 16615
rect 7428 16612 7484 16615
rect 7536 16612 7592 16615
rect 7644 16612 7700 16615
rect 7752 16612 7808 16615
rect 7860 16612 7916 16615
rect 7968 16612 8024 16615
rect 8076 16612 8132 16615
rect 8184 16612 8240 16615
rect 8292 16612 8348 16615
rect 8400 16612 8456 16615
rect 8508 16612 8564 16615
rect 8616 16612 8672 16615
rect 8724 16612 8780 16615
rect 8832 16612 9206 16615
rect 9258 16612 9314 16615
rect 9366 16612 9422 16615
rect 9474 16612 9530 16615
rect 9582 16612 9638 16615
rect 9690 16612 9746 16615
rect 9798 16612 9854 16615
rect 9906 16612 9962 16615
rect 10014 16612 10070 16615
rect 10122 16612 10178 16615
rect 10230 16612 10286 16615
rect 10338 16612 10394 16615
rect 10446 16612 10502 16615
rect 10554 16612 10610 16615
rect 10662 16612 10718 16615
rect 10770 16612 10826 16615
rect 10878 16612 10934 16615
rect 10986 16612 11042 16615
rect 11094 16612 11150 16615
rect 11202 16612 11481 16615
rect 1481 16566 1494 16612
rect 11468 16566 11481 16612
rect 1481 16563 1760 16566
rect 1812 16563 1868 16566
rect 1920 16563 1976 16566
rect 2028 16563 2084 16566
rect 2136 16563 2192 16566
rect 2244 16563 2300 16566
rect 2352 16563 2408 16566
rect 2460 16563 2516 16566
rect 2568 16563 2624 16566
rect 2676 16563 2732 16566
rect 2784 16563 2840 16566
rect 2892 16563 2948 16566
rect 3000 16563 3056 16566
rect 3108 16563 3164 16566
rect 3216 16563 3272 16566
rect 3324 16563 3380 16566
rect 3432 16563 3488 16566
rect 3540 16563 3596 16566
rect 3648 16563 3704 16566
rect 3756 16563 4130 16566
rect 4182 16563 4238 16566
rect 4290 16563 4346 16566
rect 4398 16563 4454 16566
rect 4506 16563 4562 16566
rect 4614 16563 4670 16566
rect 4722 16563 4778 16566
rect 4830 16563 4886 16566
rect 4938 16563 4994 16566
rect 5046 16563 5102 16566
rect 5154 16563 5210 16566
rect 5262 16563 5318 16566
rect 5370 16563 5426 16566
rect 5478 16563 5534 16566
rect 5586 16563 5642 16566
rect 5694 16563 5750 16566
rect 5802 16563 5858 16566
rect 5910 16563 5966 16566
rect 6018 16563 6074 16566
rect 6126 16563 6836 16566
rect 6888 16563 6944 16566
rect 6996 16563 7052 16566
rect 7104 16563 7160 16566
rect 7212 16563 7268 16566
rect 7320 16563 7376 16566
rect 7428 16563 7484 16566
rect 7536 16563 7592 16566
rect 7644 16563 7700 16566
rect 7752 16563 7808 16566
rect 7860 16563 7916 16566
rect 7968 16563 8024 16566
rect 8076 16563 8132 16566
rect 8184 16563 8240 16566
rect 8292 16563 8348 16566
rect 8400 16563 8456 16566
rect 8508 16563 8564 16566
rect 8616 16563 8672 16566
rect 8724 16563 8780 16566
rect 8832 16563 9206 16566
rect 9258 16563 9314 16566
rect 9366 16563 9422 16566
rect 9474 16563 9530 16566
rect 9582 16563 9638 16566
rect 9690 16563 9746 16566
rect 9798 16563 9854 16566
rect 9906 16563 9962 16566
rect 10014 16563 10070 16566
rect 10122 16563 10178 16566
rect 10230 16563 10286 16566
rect 10338 16563 10394 16566
rect 10446 16563 10502 16566
rect 10554 16563 10610 16566
rect 10662 16563 10718 16566
rect 10770 16563 10826 16566
rect 10878 16563 10934 16566
rect 10986 16563 11042 16566
rect 11094 16563 11150 16566
rect 11202 16563 11481 16566
rect 1481 16551 11481 16563
rect 1481 16371 11481 16383
rect 1481 16319 1493 16371
rect 1545 16368 1601 16371
rect 1653 16368 3863 16371
rect 3915 16368 3971 16371
rect 4023 16368 6239 16371
rect 6291 16368 6347 16371
rect 6399 16368 6455 16371
rect 6507 16368 6563 16371
rect 6615 16368 6671 16371
rect 6723 16368 8939 16371
rect 8991 16368 9047 16371
rect 9099 16368 11309 16371
rect 11361 16368 11417 16371
rect 1545 16319 1601 16322
rect 1653 16319 3863 16322
rect 3915 16319 3971 16322
rect 4023 16319 6239 16322
rect 6291 16319 6347 16322
rect 6399 16319 6455 16322
rect 6507 16319 6563 16322
rect 6615 16319 6671 16322
rect 6723 16319 8939 16322
rect 8991 16319 9047 16322
rect 9099 16319 11309 16322
rect 11361 16319 11417 16322
rect 11469 16319 11481 16371
rect 1481 16307 11481 16319
rect 1481 16127 11481 16139
rect 1481 16124 1760 16127
rect 1812 16124 1868 16127
rect 1920 16124 1976 16127
rect 2028 16124 2084 16127
rect 2136 16124 2192 16127
rect 2244 16124 2300 16127
rect 2352 16124 2408 16127
rect 2460 16124 2516 16127
rect 2568 16124 2624 16127
rect 2676 16124 2732 16127
rect 2784 16124 2840 16127
rect 2892 16124 2948 16127
rect 3000 16124 3056 16127
rect 3108 16124 3164 16127
rect 3216 16124 3272 16127
rect 3324 16124 3380 16127
rect 3432 16124 3488 16127
rect 3540 16124 3596 16127
rect 3648 16124 3704 16127
rect 3756 16124 4130 16127
rect 4182 16124 4238 16127
rect 4290 16124 4346 16127
rect 4398 16124 4454 16127
rect 4506 16124 4562 16127
rect 4614 16124 4670 16127
rect 4722 16124 4778 16127
rect 4830 16124 4886 16127
rect 4938 16124 4994 16127
rect 5046 16124 5102 16127
rect 5154 16124 5210 16127
rect 5262 16124 5318 16127
rect 5370 16124 5426 16127
rect 5478 16124 5534 16127
rect 5586 16124 5642 16127
rect 5694 16124 5750 16127
rect 5802 16124 5858 16127
rect 5910 16124 5966 16127
rect 6018 16124 6074 16127
rect 6126 16124 6836 16127
rect 6888 16124 6944 16127
rect 6996 16124 7052 16127
rect 7104 16124 7160 16127
rect 7212 16124 7268 16127
rect 7320 16124 7376 16127
rect 7428 16124 7484 16127
rect 7536 16124 7592 16127
rect 7644 16124 7700 16127
rect 7752 16124 7808 16127
rect 7860 16124 7916 16127
rect 7968 16124 8024 16127
rect 8076 16124 8132 16127
rect 8184 16124 8240 16127
rect 8292 16124 8348 16127
rect 8400 16124 8456 16127
rect 8508 16124 8564 16127
rect 8616 16124 8672 16127
rect 8724 16124 8780 16127
rect 8832 16124 9206 16127
rect 9258 16124 9314 16127
rect 9366 16124 9422 16127
rect 9474 16124 9530 16127
rect 9582 16124 9638 16127
rect 9690 16124 9746 16127
rect 9798 16124 9854 16127
rect 9906 16124 9962 16127
rect 10014 16124 10070 16127
rect 10122 16124 10178 16127
rect 10230 16124 10286 16127
rect 10338 16124 10394 16127
rect 10446 16124 10502 16127
rect 10554 16124 10610 16127
rect 10662 16124 10718 16127
rect 10770 16124 10826 16127
rect 10878 16124 10934 16127
rect 10986 16124 11042 16127
rect 11094 16124 11150 16127
rect 11202 16124 11481 16127
rect 1481 16078 1494 16124
rect 11468 16078 11481 16124
rect 1481 16075 1760 16078
rect 1812 16075 1868 16078
rect 1920 16075 1976 16078
rect 2028 16075 2084 16078
rect 2136 16075 2192 16078
rect 2244 16075 2300 16078
rect 2352 16075 2408 16078
rect 2460 16075 2516 16078
rect 2568 16075 2624 16078
rect 2676 16075 2732 16078
rect 2784 16075 2840 16078
rect 2892 16075 2948 16078
rect 3000 16075 3056 16078
rect 3108 16075 3164 16078
rect 3216 16075 3272 16078
rect 3324 16075 3380 16078
rect 3432 16075 3488 16078
rect 3540 16075 3596 16078
rect 3648 16075 3704 16078
rect 3756 16075 4130 16078
rect 4182 16075 4238 16078
rect 4290 16075 4346 16078
rect 4398 16075 4454 16078
rect 4506 16075 4562 16078
rect 4614 16075 4670 16078
rect 4722 16075 4778 16078
rect 4830 16075 4886 16078
rect 4938 16075 4994 16078
rect 5046 16075 5102 16078
rect 5154 16075 5210 16078
rect 5262 16075 5318 16078
rect 5370 16075 5426 16078
rect 5478 16075 5534 16078
rect 5586 16075 5642 16078
rect 5694 16075 5750 16078
rect 5802 16075 5858 16078
rect 5910 16075 5966 16078
rect 6018 16075 6074 16078
rect 6126 16075 6836 16078
rect 6888 16075 6944 16078
rect 6996 16075 7052 16078
rect 7104 16075 7160 16078
rect 7212 16075 7268 16078
rect 7320 16075 7376 16078
rect 7428 16075 7484 16078
rect 7536 16075 7592 16078
rect 7644 16075 7700 16078
rect 7752 16075 7808 16078
rect 7860 16075 7916 16078
rect 7968 16075 8024 16078
rect 8076 16075 8132 16078
rect 8184 16075 8240 16078
rect 8292 16075 8348 16078
rect 8400 16075 8456 16078
rect 8508 16075 8564 16078
rect 8616 16075 8672 16078
rect 8724 16075 8780 16078
rect 8832 16075 9206 16078
rect 9258 16075 9314 16078
rect 9366 16075 9422 16078
rect 9474 16075 9530 16078
rect 9582 16075 9638 16078
rect 9690 16075 9746 16078
rect 9798 16075 9854 16078
rect 9906 16075 9962 16078
rect 10014 16075 10070 16078
rect 10122 16075 10178 16078
rect 10230 16075 10286 16078
rect 10338 16075 10394 16078
rect 10446 16075 10502 16078
rect 10554 16075 10610 16078
rect 10662 16075 10718 16078
rect 10770 16075 10826 16078
rect 10878 16075 10934 16078
rect 10986 16075 11042 16078
rect 11094 16075 11150 16078
rect 11202 16075 11481 16078
rect 1481 16063 11481 16075
rect 1481 15883 11481 15895
rect 1481 15831 1493 15883
rect 1545 15880 1601 15883
rect 1653 15880 3863 15883
rect 3915 15880 3971 15883
rect 4023 15880 6239 15883
rect 6291 15880 6347 15883
rect 6399 15880 6455 15883
rect 6507 15880 6563 15883
rect 6615 15880 6671 15883
rect 6723 15880 8939 15883
rect 8991 15880 9047 15883
rect 9099 15880 11309 15883
rect 11361 15880 11417 15883
rect 1545 15831 1601 15834
rect 1653 15831 3863 15834
rect 3915 15831 3971 15834
rect 4023 15831 6239 15834
rect 6291 15831 6347 15834
rect 6399 15831 6455 15834
rect 6507 15831 6563 15834
rect 6615 15831 6671 15834
rect 6723 15831 8939 15834
rect 8991 15831 9047 15834
rect 9099 15831 11309 15834
rect 11361 15831 11417 15834
rect 11469 15831 11481 15883
rect 1481 15819 11481 15831
rect 1481 15639 11481 15651
rect 1481 15636 1760 15639
rect 1812 15636 1868 15639
rect 1920 15636 1976 15639
rect 2028 15636 2084 15639
rect 2136 15636 2192 15639
rect 2244 15636 2300 15639
rect 2352 15636 2408 15639
rect 2460 15636 2516 15639
rect 2568 15636 2624 15639
rect 2676 15636 2732 15639
rect 2784 15636 2840 15639
rect 2892 15636 2948 15639
rect 3000 15636 3056 15639
rect 3108 15636 3164 15639
rect 3216 15636 3272 15639
rect 3324 15636 3380 15639
rect 3432 15636 3488 15639
rect 3540 15636 3596 15639
rect 3648 15636 3704 15639
rect 3756 15636 4130 15639
rect 4182 15636 4238 15639
rect 4290 15636 4346 15639
rect 4398 15636 4454 15639
rect 4506 15636 4562 15639
rect 4614 15636 4670 15639
rect 4722 15636 4778 15639
rect 4830 15636 4886 15639
rect 4938 15636 4994 15639
rect 5046 15636 5102 15639
rect 5154 15636 5210 15639
rect 5262 15636 5318 15639
rect 5370 15636 5426 15639
rect 5478 15636 5534 15639
rect 5586 15636 5642 15639
rect 5694 15636 5750 15639
rect 5802 15636 5858 15639
rect 5910 15636 5966 15639
rect 6018 15636 6074 15639
rect 6126 15636 6836 15639
rect 6888 15636 6944 15639
rect 6996 15636 7052 15639
rect 7104 15636 7160 15639
rect 7212 15636 7268 15639
rect 7320 15636 7376 15639
rect 7428 15636 7484 15639
rect 7536 15636 7592 15639
rect 7644 15636 7700 15639
rect 7752 15636 7808 15639
rect 7860 15636 7916 15639
rect 7968 15636 8024 15639
rect 8076 15636 8132 15639
rect 8184 15636 8240 15639
rect 8292 15636 8348 15639
rect 8400 15636 8456 15639
rect 8508 15636 8564 15639
rect 8616 15636 8672 15639
rect 8724 15636 8780 15639
rect 8832 15636 9206 15639
rect 9258 15636 9314 15639
rect 9366 15636 9422 15639
rect 9474 15636 9530 15639
rect 9582 15636 9638 15639
rect 9690 15636 9746 15639
rect 9798 15636 9854 15639
rect 9906 15636 9962 15639
rect 10014 15636 10070 15639
rect 10122 15636 10178 15639
rect 10230 15636 10286 15639
rect 10338 15636 10394 15639
rect 10446 15636 10502 15639
rect 10554 15636 10610 15639
rect 10662 15636 10718 15639
rect 10770 15636 10826 15639
rect 10878 15636 10934 15639
rect 10986 15636 11042 15639
rect 11094 15636 11150 15639
rect 11202 15636 11481 15639
rect 1481 15590 1494 15636
rect 11468 15590 11481 15636
rect 1481 15587 1760 15590
rect 1812 15587 1868 15590
rect 1920 15587 1976 15590
rect 2028 15587 2084 15590
rect 2136 15587 2192 15590
rect 2244 15587 2300 15590
rect 2352 15587 2408 15590
rect 2460 15587 2516 15590
rect 2568 15587 2624 15590
rect 2676 15587 2732 15590
rect 2784 15587 2840 15590
rect 2892 15587 2948 15590
rect 3000 15587 3056 15590
rect 3108 15587 3164 15590
rect 3216 15587 3272 15590
rect 3324 15587 3380 15590
rect 3432 15587 3488 15590
rect 3540 15587 3596 15590
rect 3648 15587 3704 15590
rect 3756 15587 4130 15590
rect 4182 15587 4238 15590
rect 4290 15587 4346 15590
rect 4398 15587 4454 15590
rect 4506 15587 4562 15590
rect 4614 15587 4670 15590
rect 4722 15587 4778 15590
rect 4830 15587 4886 15590
rect 4938 15587 4994 15590
rect 5046 15587 5102 15590
rect 5154 15587 5210 15590
rect 5262 15587 5318 15590
rect 5370 15587 5426 15590
rect 5478 15587 5534 15590
rect 5586 15587 5642 15590
rect 5694 15587 5750 15590
rect 5802 15587 5858 15590
rect 5910 15587 5966 15590
rect 6018 15587 6074 15590
rect 6126 15587 6836 15590
rect 6888 15587 6944 15590
rect 6996 15587 7052 15590
rect 7104 15587 7160 15590
rect 7212 15587 7268 15590
rect 7320 15587 7376 15590
rect 7428 15587 7484 15590
rect 7536 15587 7592 15590
rect 7644 15587 7700 15590
rect 7752 15587 7808 15590
rect 7860 15587 7916 15590
rect 7968 15587 8024 15590
rect 8076 15587 8132 15590
rect 8184 15587 8240 15590
rect 8292 15587 8348 15590
rect 8400 15587 8456 15590
rect 8508 15587 8564 15590
rect 8616 15587 8672 15590
rect 8724 15587 8780 15590
rect 8832 15587 9206 15590
rect 9258 15587 9314 15590
rect 9366 15587 9422 15590
rect 9474 15587 9530 15590
rect 9582 15587 9638 15590
rect 9690 15587 9746 15590
rect 9798 15587 9854 15590
rect 9906 15587 9962 15590
rect 10014 15587 10070 15590
rect 10122 15587 10178 15590
rect 10230 15587 10286 15590
rect 10338 15587 10394 15590
rect 10446 15587 10502 15590
rect 10554 15587 10610 15590
rect 10662 15587 10718 15590
rect 10770 15587 10826 15590
rect 10878 15587 10934 15590
rect 10986 15587 11042 15590
rect 11094 15587 11150 15590
rect 11202 15587 11481 15590
rect 1481 15575 11481 15587
rect 1481 15395 11481 15407
rect 1481 15343 1493 15395
rect 1545 15392 1601 15395
rect 1653 15392 3863 15395
rect 3915 15392 3971 15395
rect 4023 15392 6239 15395
rect 6291 15392 6347 15395
rect 6399 15392 6455 15395
rect 6507 15392 6563 15395
rect 6615 15392 6671 15395
rect 6723 15392 8939 15395
rect 8991 15392 9047 15395
rect 9099 15392 11309 15395
rect 11361 15392 11417 15395
rect 1545 15343 1601 15346
rect 1653 15343 3863 15346
rect 3915 15343 3971 15346
rect 4023 15343 6239 15346
rect 6291 15343 6347 15346
rect 6399 15343 6455 15346
rect 6507 15343 6563 15346
rect 6615 15343 6671 15346
rect 6723 15343 8939 15346
rect 8991 15343 9047 15346
rect 9099 15343 11309 15346
rect 11361 15343 11417 15346
rect 11469 15343 11481 15395
rect 1481 15331 11481 15343
rect 1481 15151 11481 15163
rect 1481 15148 1760 15151
rect 1812 15148 1868 15151
rect 1920 15148 1976 15151
rect 2028 15148 2084 15151
rect 2136 15148 2192 15151
rect 2244 15148 2300 15151
rect 2352 15148 2408 15151
rect 2460 15148 2516 15151
rect 2568 15148 2624 15151
rect 2676 15148 2732 15151
rect 2784 15148 2840 15151
rect 2892 15148 2948 15151
rect 3000 15148 3056 15151
rect 3108 15148 3164 15151
rect 3216 15148 3272 15151
rect 3324 15148 3380 15151
rect 3432 15148 3488 15151
rect 3540 15148 3596 15151
rect 3648 15148 3704 15151
rect 3756 15148 4130 15151
rect 4182 15148 4238 15151
rect 4290 15148 4346 15151
rect 4398 15148 4454 15151
rect 4506 15148 4562 15151
rect 4614 15148 4670 15151
rect 4722 15148 4778 15151
rect 4830 15148 4886 15151
rect 4938 15148 4994 15151
rect 5046 15148 5102 15151
rect 5154 15148 5210 15151
rect 5262 15148 5318 15151
rect 5370 15148 5426 15151
rect 5478 15148 5534 15151
rect 5586 15148 5642 15151
rect 5694 15148 5750 15151
rect 5802 15148 5858 15151
rect 5910 15148 5966 15151
rect 6018 15148 6074 15151
rect 6126 15148 6836 15151
rect 6888 15148 6944 15151
rect 6996 15148 7052 15151
rect 7104 15148 7160 15151
rect 7212 15148 7268 15151
rect 7320 15148 7376 15151
rect 7428 15148 7484 15151
rect 7536 15148 7592 15151
rect 7644 15148 7700 15151
rect 7752 15148 7808 15151
rect 7860 15148 7916 15151
rect 7968 15148 8024 15151
rect 8076 15148 8132 15151
rect 8184 15148 8240 15151
rect 8292 15148 8348 15151
rect 8400 15148 8456 15151
rect 8508 15148 8564 15151
rect 8616 15148 8672 15151
rect 8724 15148 8780 15151
rect 8832 15148 9206 15151
rect 9258 15148 9314 15151
rect 9366 15148 9422 15151
rect 9474 15148 9530 15151
rect 9582 15148 9638 15151
rect 9690 15148 9746 15151
rect 9798 15148 9854 15151
rect 9906 15148 9962 15151
rect 10014 15148 10070 15151
rect 10122 15148 10178 15151
rect 10230 15148 10286 15151
rect 10338 15148 10394 15151
rect 10446 15148 10502 15151
rect 10554 15148 10610 15151
rect 10662 15148 10718 15151
rect 10770 15148 10826 15151
rect 10878 15148 10934 15151
rect 10986 15148 11042 15151
rect 11094 15148 11150 15151
rect 11202 15148 11481 15151
rect 1481 15102 1494 15148
rect 11468 15102 11481 15148
rect 1481 15099 1760 15102
rect 1812 15099 1868 15102
rect 1920 15099 1976 15102
rect 2028 15099 2084 15102
rect 2136 15099 2192 15102
rect 2244 15099 2300 15102
rect 2352 15099 2408 15102
rect 2460 15099 2516 15102
rect 2568 15099 2624 15102
rect 2676 15099 2732 15102
rect 2784 15099 2840 15102
rect 2892 15099 2948 15102
rect 3000 15099 3056 15102
rect 3108 15099 3164 15102
rect 3216 15099 3272 15102
rect 3324 15099 3380 15102
rect 3432 15099 3488 15102
rect 3540 15099 3596 15102
rect 3648 15099 3704 15102
rect 3756 15099 4130 15102
rect 4182 15099 4238 15102
rect 4290 15099 4346 15102
rect 4398 15099 4454 15102
rect 4506 15099 4562 15102
rect 4614 15099 4670 15102
rect 4722 15099 4778 15102
rect 4830 15099 4886 15102
rect 4938 15099 4994 15102
rect 5046 15099 5102 15102
rect 5154 15099 5210 15102
rect 5262 15099 5318 15102
rect 5370 15099 5426 15102
rect 5478 15099 5534 15102
rect 5586 15099 5642 15102
rect 5694 15099 5750 15102
rect 5802 15099 5858 15102
rect 5910 15099 5966 15102
rect 6018 15099 6074 15102
rect 6126 15099 6836 15102
rect 6888 15099 6944 15102
rect 6996 15099 7052 15102
rect 7104 15099 7160 15102
rect 7212 15099 7268 15102
rect 7320 15099 7376 15102
rect 7428 15099 7484 15102
rect 7536 15099 7592 15102
rect 7644 15099 7700 15102
rect 7752 15099 7808 15102
rect 7860 15099 7916 15102
rect 7968 15099 8024 15102
rect 8076 15099 8132 15102
rect 8184 15099 8240 15102
rect 8292 15099 8348 15102
rect 8400 15099 8456 15102
rect 8508 15099 8564 15102
rect 8616 15099 8672 15102
rect 8724 15099 8780 15102
rect 8832 15099 9206 15102
rect 9258 15099 9314 15102
rect 9366 15099 9422 15102
rect 9474 15099 9530 15102
rect 9582 15099 9638 15102
rect 9690 15099 9746 15102
rect 9798 15099 9854 15102
rect 9906 15099 9962 15102
rect 10014 15099 10070 15102
rect 10122 15099 10178 15102
rect 10230 15099 10286 15102
rect 10338 15099 10394 15102
rect 10446 15099 10502 15102
rect 10554 15099 10610 15102
rect 10662 15099 10718 15102
rect 10770 15099 10826 15102
rect 10878 15099 10934 15102
rect 10986 15099 11042 15102
rect 11094 15099 11150 15102
rect 11202 15099 11481 15102
rect 1481 15087 11481 15099
rect 1481 14907 11481 14919
rect 1481 14855 1493 14907
rect 1545 14904 1601 14907
rect 1653 14904 3863 14907
rect 3915 14904 3971 14907
rect 4023 14904 6239 14907
rect 6291 14904 6347 14907
rect 6399 14904 6455 14907
rect 6507 14904 6563 14907
rect 6615 14904 6671 14907
rect 6723 14904 8939 14907
rect 8991 14904 9047 14907
rect 9099 14904 11309 14907
rect 11361 14904 11417 14907
rect 1545 14855 1601 14858
rect 1653 14855 3863 14858
rect 3915 14855 3971 14858
rect 4023 14855 6239 14858
rect 6291 14855 6347 14858
rect 6399 14855 6455 14858
rect 6507 14855 6563 14858
rect 6615 14855 6671 14858
rect 6723 14855 8939 14858
rect 8991 14855 9047 14858
rect 9099 14855 11309 14858
rect 11361 14855 11417 14858
rect 11469 14855 11481 14907
rect 1481 14843 11481 14855
rect 1481 14663 11481 14675
rect 1481 14660 1760 14663
rect 1812 14660 1868 14663
rect 1920 14660 1976 14663
rect 2028 14660 2084 14663
rect 2136 14660 2192 14663
rect 2244 14660 2300 14663
rect 2352 14660 2408 14663
rect 2460 14660 2516 14663
rect 2568 14660 2624 14663
rect 2676 14660 2732 14663
rect 2784 14660 2840 14663
rect 2892 14660 2948 14663
rect 3000 14660 3056 14663
rect 3108 14660 3164 14663
rect 3216 14660 3272 14663
rect 3324 14660 3380 14663
rect 3432 14660 3488 14663
rect 3540 14660 3596 14663
rect 3648 14660 3704 14663
rect 3756 14660 4130 14663
rect 4182 14660 4238 14663
rect 4290 14660 4346 14663
rect 4398 14660 4454 14663
rect 4506 14660 4562 14663
rect 4614 14660 4670 14663
rect 4722 14660 4778 14663
rect 4830 14660 4886 14663
rect 4938 14660 4994 14663
rect 5046 14660 5102 14663
rect 5154 14660 5210 14663
rect 5262 14660 5318 14663
rect 5370 14660 5426 14663
rect 5478 14660 5534 14663
rect 5586 14660 5642 14663
rect 5694 14660 5750 14663
rect 5802 14660 5858 14663
rect 5910 14660 5966 14663
rect 6018 14660 6074 14663
rect 6126 14660 6836 14663
rect 6888 14660 6944 14663
rect 6996 14660 7052 14663
rect 7104 14660 7160 14663
rect 7212 14660 7268 14663
rect 7320 14660 7376 14663
rect 7428 14660 7484 14663
rect 7536 14660 7592 14663
rect 7644 14660 7700 14663
rect 7752 14660 7808 14663
rect 7860 14660 7916 14663
rect 7968 14660 8024 14663
rect 8076 14660 8132 14663
rect 8184 14660 8240 14663
rect 8292 14660 8348 14663
rect 8400 14660 8456 14663
rect 8508 14660 8564 14663
rect 8616 14660 8672 14663
rect 8724 14660 8780 14663
rect 8832 14660 9206 14663
rect 9258 14660 9314 14663
rect 9366 14660 9422 14663
rect 9474 14660 9530 14663
rect 9582 14660 9638 14663
rect 9690 14660 9746 14663
rect 9798 14660 9854 14663
rect 9906 14660 9962 14663
rect 10014 14660 10070 14663
rect 10122 14660 10178 14663
rect 10230 14660 10286 14663
rect 10338 14660 10394 14663
rect 10446 14660 10502 14663
rect 10554 14660 10610 14663
rect 10662 14660 10718 14663
rect 10770 14660 10826 14663
rect 10878 14660 10934 14663
rect 10986 14660 11042 14663
rect 11094 14660 11150 14663
rect 11202 14660 11481 14663
rect 1481 14614 1494 14660
rect 11468 14614 11481 14660
rect 1481 14611 1760 14614
rect 1812 14611 1868 14614
rect 1920 14611 1976 14614
rect 2028 14611 2084 14614
rect 2136 14611 2192 14614
rect 2244 14611 2300 14614
rect 2352 14611 2408 14614
rect 2460 14611 2516 14614
rect 2568 14611 2624 14614
rect 2676 14611 2732 14614
rect 2784 14611 2840 14614
rect 2892 14611 2948 14614
rect 3000 14611 3056 14614
rect 3108 14611 3164 14614
rect 3216 14611 3272 14614
rect 3324 14611 3380 14614
rect 3432 14611 3488 14614
rect 3540 14611 3596 14614
rect 3648 14611 3704 14614
rect 3756 14611 4130 14614
rect 4182 14611 4238 14614
rect 4290 14611 4346 14614
rect 4398 14611 4454 14614
rect 4506 14611 4562 14614
rect 4614 14611 4670 14614
rect 4722 14611 4778 14614
rect 4830 14611 4886 14614
rect 4938 14611 4994 14614
rect 5046 14611 5102 14614
rect 5154 14611 5210 14614
rect 5262 14611 5318 14614
rect 5370 14611 5426 14614
rect 5478 14611 5534 14614
rect 5586 14611 5642 14614
rect 5694 14611 5750 14614
rect 5802 14611 5858 14614
rect 5910 14611 5966 14614
rect 6018 14611 6074 14614
rect 6126 14611 6836 14614
rect 6888 14611 6944 14614
rect 6996 14611 7052 14614
rect 7104 14611 7160 14614
rect 7212 14611 7268 14614
rect 7320 14611 7376 14614
rect 7428 14611 7484 14614
rect 7536 14611 7592 14614
rect 7644 14611 7700 14614
rect 7752 14611 7808 14614
rect 7860 14611 7916 14614
rect 7968 14611 8024 14614
rect 8076 14611 8132 14614
rect 8184 14611 8240 14614
rect 8292 14611 8348 14614
rect 8400 14611 8456 14614
rect 8508 14611 8564 14614
rect 8616 14611 8672 14614
rect 8724 14611 8780 14614
rect 8832 14611 9206 14614
rect 9258 14611 9314 14614
rect 9366 14611 9422 14614
rect 9474 14611 9530 14614
rect 9582 14611 9638 14614
rect 9690 14611 9746 14614
rect 9798 14611 9854 14614
rect 9906 14611 9962 14614
rect 10014 14611 10070 14614
rect 10122 14611 10178 14614
rect 10230 14611 10286 14614
rect 10338 14611 10394 14614
rect 10446 14611 10502 14614
rect 10554 14611 10610 14614
rect 10662 14611 10718 14614
rect 10770 14611 10826 14614
rect 10878 14611 10934 14614
rect 10986 14611 11042 14614
rect 11094 14611 11150 14614
rect 11202 14611 11481 14614
rect 1481 14599 11481 14611
rect 1481 14419 11481 14431
rect 1481 14367 1493 14419
rect 1545 14416 1601 14419
rect 1653 14416 3863 14419
rect 3915 14416 3971 14419
rect 4023 14416 6239 14419
rect 6291 14416 6347 14419
rect 6399 14416 6455 14419
rect 6507 14416 6563 14419
rect 6615 14416 6671 14419
rect 6723 14416 8939 14419
rect 8991 14416 9047 14419
rect 9099 14416 11309 14419
rect 11361 14416 11417 14419
rect 1545 14367 1601 14370
rect 1653 14367 3863 14370
rect 3915 14367 3971 14370
rect 4023 14367 6239 14370
rect 6291 14367 6347 14370
rect 6399 14367 6455 14370
rect 6507 14367 6563 14370
rect 6615 14367 6671 14370
rect 6723 14367 8939 14370
rect 8991 14367 9047 14370
rect 9099 14367 11309 14370
rect 11361 14367 11417 14370
rect 11469 14367 11481 14419
rect 1481 14355 11481 14367
rect 1481 14175 11481 14187
rect 1481 14172 1760 14175
rect 1812 14172 1868 14175
rect 1920 14172 1976 14175
rect 2028 14172 2084 14175
rect 2136 14172 2192 14175
rect 2244 14172 2300 14175
rect 2352 14172 2408 14175
rect 2460 14172 2516 14175
rect 2568 14172 2624 14175
rect 2676 14172 2732 14175
rect 2784 14172 2840 14175
rect 2892 14172 2948 14175
rect 3000 14172 3056 14175
rect 3108 14172 3164 14175
rect 3216 14172 3272 14175
rect 3324 14172 3380 14175
rect 3432 14172 3488 14175
rect 3540 14172 3596 14175
rect 3648 14172 3704 14175
rect 3756 14172 4130 14175
rect 4182 14172 4238 14175
rect 4290 14172 4346 14175
rect 4398 14172 4454 14175
rect 4506 14172 4562 14175
rect 4614 14172 4670 14175
rect 4722 14172 4778 14175
rect 4830 14172 4886 14175
rect 4938 14172 4994 14175
rect 5046 14172 5102 14175
rect 5154 14172 5210 14175
rect 5262 14172 5318 14175
rect 5370 14172 5426 14175
rect 5478 14172 5534 14175
rect 5586 14172 5642 14175
rect 5694 14172 5750 14175
rect 5802 14172 5858 14175
rect 5910 14172 5966 14175
rect 6018 14172 6074 14175
rect 6126 14172 6836 14175
rect 6888 14172 6944 14175
rect 6996 14172 7052 14175
rect 7104 14172 7160 14175
rect 7212 14172 7268 14175
rect 7320 14172 7376 14175
rect 7428 14172 7484 14175
rect 7536 14172 7592 14175
rect 7644 14172 7700 14175
rect 7752 14172 7808 14175
rect 7860 14172 7916 14175
rect 7968 14172 8024 14175
rect 8076 14172 8132 14175
rect 8184 14172 8240 14175
rect 8292 14172 8348 14175
rect 8400 14172 8456 14175
rect 8508 14172 8564 14175
rect 8616 14172 8672 14175
rect 8724 14172 8780 14175
rect 8832 14172 9206 14175
rect 9258 14172 9314 14175
rect 9366 14172 9422 14175
rect 9474 14172 9530 14175
rect 9582 14172 9638 14175
rect 9690 14172 9746 14175
rect 9798 14172 9854 14175
rect 9906 14172 9962 14175
rect 10014 14172 10070 14175
rect 10122 14172 10178 14175
rect 10230 14172 10286 14175
rect 10338 14172 10394 14175
rect 10446 14172 10502 14175
rect 10554 14172 10610 14175
rect 10662 14172 10718 14175
rect 10770 14172 10826 14175
rect 10878 14172 10934 14175
rect 10986 14172 11042 14175
rect 11094 14172 11150 14175
rect 11202 14172 11481 14175
rect 1481 14126 1494 14172
rect 11468 14126 11481 14172
rect 1481 14123 1760 14126
rect 1812 14123 1868 14126
rect 1920 14123 1976 14126
rect 2028 14123 2084 14126
rect 2136 14123 2192 14126
rect 2244 14123 2300 14126
rect 2352 14123 2408 14126
rect 2460 14123 2516 14126
rect 2568 14123 2624 14126
rect 2676 14123 2732 14126
rect 2784 14123 2840 14126
rect 2892 14123 2948 14126
rect 3000 14123 3056 14126
rect 3108 14123 3164 14126
rect 3216 14123 3272 14126
rect 3324 14123 3380 14126
rect 3432 14123 3488 14126
rect 3540 14123 3596 14126
rect 3648 14123 3704 14126
rect 3756 14123 4130 14126
rect 4182 14123 4238 14126
rect 4290 14123 4346 14126
rect 4398 14123 4454 14126
rect 4506 14123 4562 14126
rect 4614 14123 4670 14126
rect 4722 14123 4778 14126
rect 4830 14123 4886 14126
rect 4938 14123 4994 14126
rect 5046 14123 5102 14126
rect 5154 14123 5210 14126
rect 5262 14123 5318 14126
rect 5370 14123 5426 14126
rect 5478 14123 5534 14126
rect 5586 14123 5642 14126
rect 5694 14123 5750 14126
rect 5802 14123 5858 14126
rect 5910 14123 5966 14126
rect 6018 14123 6074 14126
rect 6126 14123 6836 14126
rect 6888 14123 6944 14126
rect 6996 14123 7052 14126
rect 7104 14123 7160 14126
rect 7212 14123 7268 14126
rect 7320 14123 7376 14126
rect 7428 14123 7484 14126
rect 7536 14123 7592 14126
rect 7644 14123 7700 14126
rect 7752 14123 7808 14126
rect 7860 14123 7916 14126
rect 7968 14123 8024 14126
rect 8076 14123 8132 14126
rect 8184 14123 8240 14126
rect 8292 14123 8348 14126
rect 8400 14123 8456 14126
rect 8508 14123 8564 14126
rect 8616 14123 8672 14126
rect 8724 14123 8780 14126
rect 8832 14123 9206 14126
rect 9258 14123 9314 14126
rect 9366 14123 9422 14126
rect 9474 14123 9530 14126
rect 9582 14123 9638 14126
rect 9690 14123 9746 14126
rect 9798 14123 9854 14126
rect 9906 14123 9962 14126
rect 10014 14123 10070 14126
rect 10122 14123 10178 14126
rect 10230 14123 10286 14126
rect 10338 14123 10394 14126
rect 10446 14123 10502 14126
rect 10554 14123 10610 14126
rect 10662 14123 10718 14126
rect 10770 14123 10826 14126
rect 10878 14123 10934 14126
rect 10986 14123 11042 14126
rect 11094 14123 11150 14126
rect 11202 14123 11481 14126
rect 1481 14111 11481 14123
rect 1481 13931 11481 13943
rect 1481 13879 1493 13931
rect 1545 13928 1601 13931
rect 1653 13928 3863 13931
rect 3915 13928 3971 13931
rect 4023 13928 6239 13931
rect 6291 13928 6347 13931
rect 6399 13928 6455 13931
rect 6507 13928 6563 13931
rect 6615 13928 6671 13931
rect 6723 13928 8939 13931
rect 8991 13928 9047 13931
rect 9099 13928 11309 13931
rect 11361 13928 11417 13931
rect 1545 13879 1601 13882
rect 1653 13879 3863 13882
rect 3915 13879 3971 13882
rect 4023 13879 6239 13882
rect 6291 13879 6347 13882
rect 6399 13879 6455 13882
rect 6507 13879 6563 13882
rect 6615 13879 6671 13882
rect 6723 13879 8939 13882
rect 8991 13879 9047 13882
rect 9099 13879 11309 13882
rect 11361 13879 11417 13882
rect 11469 13879 11481 13931
rect 1481 13867 11481 13879
rect 1481 13687 11481 13699
rect 1481 13684 1760 13687
rect 1812 13684 1868 13687
rect 1920 13684 1976 13687
rect 2028 13684 2084 13687
rect 2136 13684 2192 13687
rect 2244 13684 2300 13687
rect 2352 13684 2408 13687
rect 2460 13684 2516 13687
rect 2568 13684 2624 13687
rect 2676 13684 2732 13687
rect 2784 13684 2840 13687
rect 2892 13684 2948 13687
rect 3000 13684 3056 13687
rect 3108 13684 3164 13687
rect 3216 13684 3272 13687
rect 3324 13684 3380 13687
rect 3432 13684 3488 13687
rect 3540 13684 3596 13687
rect 3648 13684 3704 13687
rect 3756 13684 4130 13687
rect 4182 13684 4238 13687
rect 4290 13684 4346 13687
rect 4398 13684 4454 13687
rect 4506 13684 4562 13687
rect 4614 13684 4670 13687
rect 4722 13684 4778 13687
rect 4830 13684 4886 13687
rect 4938 13684 4994 13687
rect 5046 13684 5102 13687
rect 5154 13684 5210 13687
rect 5262 13684 5318 13687
rect 5370 13684 5426 13687
rect 5478 13684 5534 13687
rect 5586 13684 5642 13687
rect 5694 13684 5750 13687
rect 5802 13684 5858 13687
rect 5910 13684 5966 13687
rect 6018 13684 6074 13687
rect 6126 13684 6836 13687
rect 6888 13684 6944 13687
rect 6996 13684 7052 13687
rect 7104 13684 7160 13687
rect 7212 13684 7268 13687
rect 7320 13684 7376 13687
rect 7428 13684 7484 13687
rect 7536 13684 7592 13687
rect 7644 13684 7700 13687
rect 7752 13684 7808 13687
rect 7860 13684 7916 13687
rect 7968 13684 8024 13687
rect 8076 13684 8132 13687
rect 8184 13684 8240 13687
rect 8292 13684 8348 13687
rect 8400 13684 8456 13687
rect 8508 13684 8564 13687
rect 8616 13684 8672 13687
rect 8724 13684 8780 13687
rect 8832 13684 9206 13687
rect 9258 13684 9314 13687
rect 9366 13684 9422 13687
rect 9474 13684 9530 13687
rect 9582 13684 9638 13687
rect 9690 13684 9746 13687
rect 9798 13684 9854 13687
rect 9906 13684 9962 13687
rect 10014 13684 10070 13687
rect 10122 13684 10178 13687
rect 10230 13684 10286 13687
rect 10338 13684 10394 13687
rect 10446 13684 10502 13687
rect 10554 13684 10610 13687
rect 10662 13684 10718 13687
rect 10770 13684 10826 13687
rect 10878 13684 10934 13687
rect 10986 13684 11042 13687
rect 11094 13684 11150 13687
rect 11202 13684 11481 13687
rect 1481 13638 1494 13684
rect 11468 13638 11481 13684
rect 1481 13635 1760 13638
rect 1812 13635 1868 13638
rect 1920 13635 1976 13638
rect 2028 13635 2084 13638
rect 2136 13635 2192 13638
rect 2244 13635 2300 13638
rect 2352 13635 2408 13638
rect 2460 13635 2516 13638
rect 2568 13635 2624 13638
rect 2676 13635 2732 13638
rect 2784 13635 2840 13638
rect 2892 13635 2948 13638
rect 3000 13635 3056 13638
rect 3108 13635 3164 13638
rect 3216 13635 3272 13638
rect 3324 13635 3380 13638
rect 3432 13635 3488 13638
rect 3540 13635 3596 13638
rect 3648 13635 3704 13638
rect 3756 13635 4130 13638
rect 4182 13635 4238 13638
rect 4290 13635 4346 13638
rect 4398 13635 4454 13638
rect 4506 13635 4562 13638
rect 4614 13635 4670 13638
rect 4722 13635 4778 13638
rect 4830 13635 4886 13638
rect 4938 13635 4994 13638
rect 5046 13635 5102 13638
rect 5154 13635 5210 13638
rect 5262 13635 5318 13638
rect 5370 13635 5426 13638
rect 5478 13635 5534 13638
rect 5586 13635 5642 13638
rect 5694 13635 5750 13638
rect 5802 13635 5858 13638
rect 5910 13635 5966 13638
rect 6018 13635 6074 13638
rect 6126 13635 6836 13638
rect 6888 13635 6944 13638
rect 6996 13635 7052 13638
rect 7104 13635 7160 13638
rect 7212 13635 7268 13638
rect 7320 13635 7376 13638
rect 7428 13635 7484 13638
rect 7536 13635 7592 13638
rect 7644 13635 7700 13638
rect 7752 13635 7808 13638
rect 7860 13635 7916 13638
rect 7968 13635 8024 13638
rect 8076 13635 8132 13638
rect 8184 13635 8240 13638
rect 8292 13635 8348 13638
rect 8400 13635 8456 13638
rect 8508 13635 8564 13638
rect 8616 13635 8672 13638
rect 8724 13635 8780 13638
rect 8832 13635 9206 13638
rect 9258 13635 9314 13638
rect 9366 13635 9422 13638
rect 9474 13635 9530 13638
rect 9582 13635 9638 13638
rect 9690 13635 9746 13638
rect 9798 13635 9854 13638
rect 9906 13635 9962 13638
rect 10014 13635 10070 13638
rect 10122 13635 10178 13638
rect 10230 13635 10286 13638
rect 10338 13635 10394 13638
rect 10446 13635 10502 13638
rect 10554 13635 10610 13638
rect 10662 13635 10718 13638
rect 10770 13635 10826 13638
rect 10878 13635 10934 13638
rect 10986 13635 11042 13638
rect 11094 13635 11150 13638
rect 11202 13635 11481 13638
rect 1481 13623 11481 13635
rect 1481 13443 11481 13455
rect 1481 13391 1493 13443
rect 1545 13440 1601 13443
rect 1653 13440 3863 13443
rect 3915 13440 3971 13443
rect 4023 13440 6239 13443
rect 6291 13440 6347 13443
rect 6399 13440 6455 13443
rect 6507 13440 6563 13443
rect 6615 13440 6671 13443
rect 6723 13440 8939 13443
rect 8991 13440 9047 13443
rect 9099 13440 11309 13443
rect 11361 13440 11417 13443
rect 1545 13391 1601 13394
rect 1653 13391 3863 13394
rect 3915 13391 3971 13394
rect 4023 13391 6239 13394
rect 6291 13391 6347 13394
rect 6399 13391 6455 13394
rect 6507 13391 6563 13394
rect 6615 13391 6671 13394
rect 6723 13391 8939 13394
rect 8991 13391 9047 13394
rect 9099 13391 11309 13394
rect 11361 13391 11417 13394
rect 11469 13391 11481 13443
rect 1481 13379 11481 13391
rect 1213 13263 1413 13290
rect 1213 13211 1233 13263
rect 1285 13211 1341 13263
rect 1393 13211 1413 13263
rect 11549 13290 11560 17936
rect 11706 17907 11749 17936
rect 11729 17855 11749 17907
rect 11706 17799 11749 17855
rect 11729 17747 11749 17799
rect 11706 17691 11749 17747
rect 11729 17639 11749 17691
rect 11706 17583 11749 17639
rect 11729 17531 11749 17583
rect 11706 17475 11749 17531
rect 11729 17423 11749 17475
rect 11706 17367 11749 17423
rect 11729 17315 11749 17367
rect 11706 17259 11749 17315
rect 11729 17207 11749 17259
rect 11706 17151 11749 17207
rect 11729 17099 11749 17151
rect 11706 17043 11749 17099
rect 11729 16991 11749 17043
rect 11706 16935 11749 16991
rect 11729 16883 11749 16935
rect 11706 16827 11749 16883
rect 11729 16775 11749 16827
rect 11706 16719 11749 16775
rect 11729 16667 11749 16719
rect 11706 16611 11749 16667
rect 11729 16559 11749 16611
rect 11706 16503 11749 16559
rect 11729 16451 11749 16503
rect 11706 16395 11749 16451
rect 11729 16343 11749 16395
rect 11706 16287 11749 16343
rect 11729 16235 11749 16287
rect 11706 16179 11749 16235
rect 11729 16127 11749 16179
rect 11706 16071 11749 16127
rect 11729 16019 11749 16071
rect 11706 15963 11749 16019
rect 11729 15911 11749 15963
rect 11706 15855 11749 15911
rect 11729 15803 11749 15855
rect 11706 15747 11749 15803
rect 11729 15695 11749 15747
rect 11706 15639 11749 15695
rect 11729 15587 11749 15639
rect 11706 15531 11749 15587
rect 11729 15479 11749 15531
rect 11706 15423 11749 15479
rect 11729 15371 11749 15423
rect 11706 15315 11749 15371
rect 11729 15263 11749 15315
rect 11706 15207 11749 15263
rect 11729 15155 11749 15207
rect 11706 15099 11749 15155
rect 11729 15047 11749 15099
rect 11706 14991 11749 15047
rect 11729 14939 11749 14991
rect 11706 14883 11749 14939
rect 11729 14831 11749 14883
rect 11706 14775 11749 14831
rect 11729 14723 11749 14775
rect 11706 14667 11749 14723
rect 11729 14615 11749 14667
rect 11706 14559 11749 14615
rect 11729 14507 11749 14559
rect 11706 14451 11749 14507
rect 11729 14399 11749 14451
rect 11706 14343 11749 14399
rect 11729 14291 11749 14343
rect 11706 14235 11749 14291
rect 11729 14183 11749 14235
rect 11706 14127 11749 14183
rect 11729 14075 11749 14127
rect 11706 14019 11749 14075
rect 11729 13967 11749 14019
rect 11706 13911 11749 13967
rect 11729 13859 11749 13911
rect 11706 13803 11749 13859
rect 11729 13751 11749 13803
rect 11706 13695 11749 13751
rect 11729 13643 11749 13695
rect 11706 13587 11749 13643
rect 11729 13535 11749 13587
rect 11706 13479 11749 13535
rect 11729 13427 11749 13479
rect 11706 13371 11749 13427
rect 11729 13319 11749 13371
rect 11706 13290 11749 13319
rect 11549 13263 11749 13290
rect 11549 13211 11569 13263
rect 11621 13211 11677 13263
rect 11729 13211 11749 13263
rect 1213 13048 1413 13211
rect 1481 13199 11481 13211
rect 1481 13196 1760 13199
rect 1812 13196 1868 13199
rect 1920 13196 1976 13199
rect 2028 13196 2084 13199
rect 2136 13196 2192 13199
rect 2244 13196 2300 13199
rect 2352 13196 2408 13199
rect 2460 13196 2516 13199
rect 2568 13196 2624 13199
rect 2676 13196 2732 13199
rect 2784 13196 2840 13199
rect 2892 13196 2948 13199
rect 3000 13196 3056 13199
rect 3108 13196 3164 13199
rect 3216 13196 3272 13199
rect 3324 13196 3380 13199
rect 3432 13196 3488 13199
rect 3540 13196 3596 13199
rect 3648 13196 3704 13199
rect 3756 13196 4130 13199
rect 4182 13196 4238 13199
rect 4290 13196 4346 13199
rect 4398 13196 4454 13199
rect 4506 13196 4562 13199
rect 4614 13196 4670 13199
rect 4722 13196 4778 13199
rect 4830 13196 4886 13199
rect 4938 13196 4994 13199
rect 5046 13196 5102 13199
rect 5154 13196 5210 13199
rect 5262 13196 5318 13199
rect 5370 13196 5426 13199
rect 5478 13196 5534 13199
rect 5586 13196 5642 13199
rect 5694 13196 5750 13199
rect 5802 13196 5858 13199
rect 5910 13196 5966 13199
rect 6018 13196 6074 13199
rect 6126 13196 6836 13199
rect 6888 13196 6944 13199
rect 6996 13196 7052 13199
rect 7104 13196 7160 13199
rect 7212 13196 7268 13199
rect 7320 13196 7376 13199
rect 7428 13196 7484 13199
rect 7536 13196 7592 13199
rect 7644 13196 7700 13199
rect 7752 13196 7808 13199
rect 7860 13196 7916 13199
rect 7968 13196 8024 13199
rect 8076 13196 8132 13199
rect 8184 13196 8240 13199
rect 8292 13196 8348 13199
rect 8400 13196 8456 13199
rect 8508 13196 8564 13199
rect 8616 13196 8672 13199
rect 8724 13196 8780 13199
rect 8832 13196 9206 13199
rect 9258 13196 9314 13199
rect 9366 13196 9422 13199
rect 9474 13196 9530 13199
rect 9582 13196 9638 13199
rect 9690 13196 9746 13199
rect 9798 13196 9854 13199
rect 9906 13196 9962 13199
rect 10014 13196 10070 13199
rect 10122 13196 10178 13199
rect 10230 13196 10286 13199
rect 10338 13196 10394 13199
rect 10446 13196 10502 13199
rect 10554 13196 10610 13199
rect 10662 13196 10718 13199
rect 10770 13196 10826 13199
rect 10878 13196 10934 13199
rect 10986 13196 11042 13199
rect 11094 13196 11150 13199
rect 11202 13196 11481 13199
rect 1481 13150 1494 13196
rect 11468 13150 11481 13196
rect 1481 13147 1760 13150
rect 1812 13147 1868 13150
rect 1920 13147 1976 13150
rect 2028 13147 2084 13150
rect 2136 13147 2192 13150
rect 2244 13147 2300 13150
rect 2352 13147 2408 13150
rect 2460 13147 2516 13150
rect 2568 13147 2624 13150
rect 2676 13147 2732 13150
rect 2784 13147 2840 13150
rect 2892 13147 2948 13150
rect 3000 13147 3056 13150
rect 3108 13147 3164 13150
rect 3216 13147 3272 13150
rect 3324 13147 3380 13150
rect 3432 13147 3488 13150
rect 3540 13147 3596 13150
rect 3648 13147 3704 13150
rect 3756 13147 4130 13150
rect 4182 13147 4238 13150
rect 4290 13147 4346 13150
rect 4398 13147 4454 13150
rect 4506 13147 4562 13150
rect 4614 13147 4670 13150
rect 4722 13147 4778 13150
rect 4830 13147 4886 13150
rect 4938 13147 4994 13150
rect 5046 13147 5102 13150
rect 5154 13147 5210 13150
rect 5262 13147 5318 13150
rect 5370 13147 5426 13150
rect 5478 13147 5534 13150
rect 5586 13147 5642 13150
rect 5694 13147 5750 13150
rect 5802 13147 5858 13150
rect 5910 13147 5966 13150
rect 6018 13147 6074 13150
rect 6126 13147 6836 13150
rect 6888 13147 6944 13150
rect 6996 13147 7052 13150
rect 7104 13147 7160 13150
rect 7212 13147 7268 13150
rect 7320 13147 7376 13150
rect 7428 13147 7484 13150
rect 7536 13147 7592 13150
rect 7644 13147 7700 13150
rect 7752 13147 7808 13150
rect 7860 13147 7916 13150
rect 7968 13147 8024 13150
rect 8076 13147 8132 13150
rect 8184 13147 8240 13150
rect 8292 13147 8348 13150
rect 8400 13147 8456 13150
rect 8508 13147 8564 13150
rect 8616 13147 8672 13150
rect 8724 13147 8780 13150
rect 8832 13147 9206 13150
rect 9258 13147 9314 13150
rect 9366 13147 9422 13150
rect 9474 13147 9530 13150
rect 9582 13147 9638 13150
rect 9690 13147 9746 13150
rect 9798 13147 9854 13150
rect 9906 13147 9962 13150
rect 10014 13147 10070 13150
rect 10122 13147 10178 13150
rect 10230 13147 10286 13150
rect 10338 13147 10394 13150
rect 10446 13147 10502 13150
rect 10554 13147 10610 13150
rect 10662 13147 10718 13150
rect 10770 13147 10826 13150
rect 10878 13147 10934 13150
rect 10986 13147 11042 13150
rect 11094 13147 11150 13150
rect 11202 13147 11481 13150
rect 1481 13135 11481 13147
rect 11549 13048 11749 13211
rect 1213 12848 11749 13048
rect 12001 12769 12012 18457
rect 950 12757 12012 12769
rect 950 12750 1760 12757
rect 1812 12750 1868 12757
rect 1920 12750 1976 12757
rect 2028 12750 2084 12757
rect 2136 12750 2192 12757
rect 2244 12750 2300 12757
rect 2352 12750 2408 12757
rect 2460 12750 2516 12757
rect 2568 12750 2624 12757
rect 2676 12750 2732 12757
rect 2784 12750 2840 12757
rect 2892 12750 2948 12757
rect 3000 12750 3056 12757
rect 3108 12750 3164 12757
rect 3216 12750 3272 12757
rect 3324 12750 3380 12757
rect 3432 12750 3488 12757
rect 3540 12750 3596 12757
rect 3648 12750 3704 12757
rect 3756 12750 4130 12757
rect 4182 12750 4238 12757
rect 4290 12750 4346 12757
rect 4398 12750 4454 12757
rect 4506 12750 4562 12757
rect 4614 12750 4670 12757
rect 4722 12750 4778 12757
rect 4830 12750 4886 12757
rect 4938 12750 4994 12757
rect 5046 12750 5102 12757
rect 5154 12750 5210 12757
rect 5262 12750 5318 12757
rect 5370 12750 5426 12757
rect 5478 12750 5534 12757
rect 5586 12750 5642 12757
rect 5694 12750 5750 12757
rect 5802 12750 5858 12757
rect 5910 12750 5966 12757
rect 6018 12750 6074 12757
rect 6126 12750 6836 12757
rect 6888 12750 6944 12757
rect 6996 12750 7052 12757
rect 7104 12750 7160 12757
rect 7212 12750 7268 12757
rect 7320 12750 7376 12757
rect 7428 12750 7484 12757
rect 7536 12750 7592 12757
rect 7644 12750 7700 12757
rect 7752 12750 7808 12757
rect 7860 12750 7916 12757
rect 7968 12750 8024 12757
rect 8076 12750 8132 12757
rect 8184 12750 8240 12757
rect 8292 12750 8348 12757
rect 8400 12750 8456 12757
rect 8508 12750 8564 12757
rect 8616 12750 8672 12757
rect 8724 12750 8780 12757
rect 8832 12750 9206 12757
rect 9258 12750 9314 12757
rect 9366 12750 9422 12757
rect 9474 12750 9530 12757
rect 9582 12750 9638 12757
rect 9690 12750 9746 12757
rect 9798 12750 9854 12757
rect 9906 12750 9962 12757
rect 10014 12750 10070 12757
rect 10122 12750 10178 12757
rect 10230 12750 10286 12757
rect 10338 12750 10394 12757
rect 10446 12750 10502 12757
rect 10554 12750 10610 12757
rect 10662 12750 10718 12757
rect 10770 12750 10826 12757
rect 10878 12750 10934 12757
rect 10986 12750 11042 12757
rect 11094 12750 11150 12757
rect 11202 12750 12012 12757
rect 950 12604 1058 12750
rect 11904 12604 12012 12750
rect 950 12597 1760 12604
rect 1812 12597 1868 12604
rect 1920 12597 1976 12604
rect 2028 12597 2084 12604
rect 2136 12597 2192 12604
rect 2244 12597 2300 12604
rect 2352 12597 2408 12604
rect 2460 12597 2516 12604
rect 2568 12597 2624 12604
rect 2676 12597 2732 12604
rect 2784 12597 2840 12604
rect 2892 12597 2948 12604
rect 3000 12597 3056 12604
rect 3108 12597 3164 12604
rect 3216 12597 3272 12604
rect 3324 12597 3380 12604
rect 3432 12597 3488 12604
rect 3540 12597 3596 12604
rect 3648 12597 3704 12604
rect 3756 12597 4130 12604
rect 4182 12597 4238 12604
rect 4290 12597 4346 12604
rect 4398 12597 4454 12604
rect 4506 12597 4562 12604
rect 4614 12597 4670 12604
rect 4722 12597 4778 12604
rect 4830 12597 4886 12604
rect 4938 12597 4994 12604
rect 5046 12597 5102 12604
rect 5154 12597 5210 12604
rect 5262 12597 5318 12604
rect 5370 12597 5426 12604
rect 5478 12597 5534 12604
rect 5586 12597 5642 12604
rect 5694 12597 5750 12604
rect 5802 12597 5858 12604
rect 5910 12597 5966 12604
rect 6018 12597 6074 12604
rect 6126 12597 6836 12604
rect 6888 12597 6944 12604
rect 6996 12597 7052 12604
rect 7104 12597 7160 12604
rect 7212 12597 7268 12604
rect 7320 12597 7376 12604
rect 7428 12597 7484 12604
rect 7536 12597 7592 12604
rect 7644 12597 7700 12604
rect 7752 12597 7808 12604
rect 7860 12597 7916 12604
rect 7968 12597 8024 12604
rect 8076 12597 8132 12604
rect 8184 12597 8240 12604
rect 8292 12597 8348 12604
rect 8400 12597 8456 12604
rect 8508 12597 8564 12604
rect 8616 12597 8672 12604
rect 8724 12597 8780 12604
rect 8832 12597 9206 12604
rect 9258 12597 9314 12604
rect 9366 12597 9422 12604
rect 9474 12597 9530 12604
rect 9582 12597 9638 12604
rect 9690 12597 9746 12604
rect 9798 12597 9854 12604
rect 9906 12597 9962 12604
rect 10014 12597 10070 12604
rect 10122 12597 10178 12604
rect 10230 12597 10286 12604
rect 10338 12597 10394 12604
rect 10446 12597 10502 12604
rect 10554 12597 10610 12604
rect 10662 12597 10718 12604
rect 10770 12597 10826 12604
rect 10878 12597 10934 12604
rect 10986 12597 11042 12604
rect 11094 12597 11150 12604
rect 11202 12597 12012 12604
rect 950 12585 12012 12597
rect 950 6897 961 12585
rect 1213 12306 11749 12506
rect 1213 12143 1413 12306
rect 1481 12207 11481 12219
rect 1481 12204 1760 12207
rect 1812 12204 1868 12207
rect 1920 12204 1976 12207
rect 2028 12204 2084 12207
rect 2136 12204 2192 12207
rect 2244 12204 2300 12207
rect 2352 12204 2408 12207
rect 2460 12204 2516 12207
rect 2568 12204 2624 12207
rect 2676 12204 2732 12207
rect 2784 12204 2840 12207
rect 2892 12204 2948 12207
rect 3000 12204 3056 12207
rect 3108 12204 3164 12207
rect 3216 12204 3272 12207
rect 3324 12204 3380 12207
rect 3432 12204 3488 12207
rect 3540 12204 3596 12207
rect 3648 12204 3704 12207
rect 3756 12204 4130 12207
rect 4182 12204 4238 12207
rect 4290 12204 4346 12207
rect 4398 12204 4454 12207
rect 4506 12204 4562 12207
rect 4614 12204 4670 12207
rect 4722 12204 4778 12207
rect 4830 12204 4886 12207
rect 4938 12204 4994 12207
rect 5046 12204 5102 12207
rect 5154 12204 5210 12207
rect 5262 12204 5318 12207
rect 5370 12204 5426 12207
rect 5478 12204 5534 12207
rect 5586 12204 5642 12207
rect 5694 12204 5750 12207
rect 5802 12204 5858 12207
rect 5910 12204 5966 12207
rect 6018 12204 6074 12207
rect 6126 12204 6836 12207
rect 6888 12204 6944 12207
rect 6996 12204 7052 12207
rect 7104 12204 7160 12207
rect 7212 12204 7268 12207
rect 7320 12204 7376 12207
rect 7428 12204 7484 12207
rect 7536 12204 7592 12207
rect 7644 12204 7700 12207
rect 7752 12204 7808 12207
rect 7860 12204 7916 12207
rect 7968 12204 8024 12207
rect 8076 12204 8132 12207
rect 8184 12204 8240 12207
rect 8292 12204 8348 12207
rect 8400 12204 8456 12207
rect 8508 12204 8564 12207
rect 8616 12204 8672 12207
rect 8724 12204 8780 12207
rect 8832 12204 9206 12207
rect 9258 12204 9314 12207
rect 9366 12204 9422 12207
rect 9474 12204 9530 12207
rect 9582 12204 9638 12207
rect 9690 12204 9746 12207
rect 9798 12204 9854 12207
rect 9906 12204 9962 12207
rect 10014 12204 10070 12207
rect 10122 12204 10178 12207
rect 10230 12204 10286 12207
rect 10338 12204 10394 12207
rect 10446 12204 10502 12207
rect 10554 12204 10610 12207
rect 10662 12204 10718 12207
rect 10770 12204 10826 12207
rect 10878 12204 10934 12207
rect 10986 12204 11042 12207
rect 11094 12204 11150 12207
rect 11202 12204 11481 12207
rect 1481 12158 1494 12204
rect 11468 12158 11481 12204
rect 1481 12155 1760 12158
rect 1812 12155 1868 12158
rect 1920 12155 1976 12158
rect 2028 12155 2084 12158
rect 2136 12155 2192 12158
rect 2244 12155 2300 12158
rect 2352 12155 2408 12158
rect 2460 12155 2516 12158
rect 2568 12155 2624 12158
rect 2676 12155 2732 12158
rect 2784 12155 2840 12158
rect 2892 12155 2948 12158
rect 3000 12155 3056 12158
rect 3108 12155 3164 12158
rect 3216 12155 3272 12158
rect 3324 12155 3380 12158
rect 3432 12155 3488 12158
rect 3540 12155 3596 12158
rect 3648 12155 3704 12158
rect 3756 12155 4130 12158
rect 4182 12155 4238 12158
rect 4290 12155 4346 12158
rect 4398 12155 4454 12158
rect 4506 12155 4562 12158
rect 4614 12155 4670 12158
rect 4722 12155 4778 12158
rect 4830 12155 4886 12158
rect 4938 12155 4994 12158
rect 5046 12155 5102 12158
rect 5154 12155 5210 12158
rect 5262 12155 5318 12158
rect 5370 12155 5426 12158
rect 5478 12155 5534 12158
rect 5586 12155 5642 12158
rect 5694 12155 5750 12158
rect 5802 12155 5858 12158
rect 5910 12155 5966 12158
rect 6018 12155 6074 12158
rect 6126 12155 6836 12158
rect 6888 12155 6944 12158
rect 6996 12155 7052 12158
rect 7104 12155 7160 12158
rect 7212 12155 7268 12158
rect 7320 12155 7376 12158
rect 7428 12155 7484 12158
rect 7536 12155 7592 12158
rect 7644 12155 7700 12158
rect 7752 12155 7808 12158
rect 7860 12155 7916 12158
rect 7968 12155 8024 12158
rect 8076 12155 8132 12158
rect 8184 12155 8240 12158
rect 8292 12155 8348 12158
rect 8400 12155 8456 12158
rect 8508 12155 8564 12158
rect 8616 12155 8672 12158
rect 8724 12155 8780 12158
rect 8832 12155 9206 12158
rect 9258 12155 9314 12158
rect 9366 12155 9422 12158
rect 9474 12155 9530 12158
rect 9582 12155 9638 12158
rect 9690 12155 9746 12158
rect 9798 12155 9854 12158
rect 9906 12155 9962 12158
rect 10014 12155 10070 12158
rect 10122 12155 10178 12158
rect 10230 12155 10286 12158
rect 10338 12155 10394 12158
rect 10446 12155 10502 12158
rect 10554 12155 10610 12158
rect 10662 12155 10718 12158
rect 10770 12155 10826 12158
rect 10878 12155 10934 12158
rect 10986 12155 11042 12158
rect 11094 12155 11150 12158
rect 11202 12155 11481 12158
rect 1481 12143 11481 12155
rect 11549 12143 11749 12306
rect 1213 12091 1233 12143
rect 1285 12091 1341 12143
rect 1393 12091 1413 12143
rect 1213 12064 1413 12091
rect 1213 12035 1256 12064
rect 1213 11983 1233 12035
rect 1213 11927 1256 11983
rect 1213 11875 1233 11927
rect 1213 11819 1256 11875
rect 1213 11767 1233 11819
rect 1213 11711 1256 11767
rect 1213 11659 1233 11711
rect 1213 11603 1256 11659
rect 1213 11551 1233 11603
rect 1213 11495 1256 11551
rect 1213 11443 1233 11495
rect 1213 11387 1256 11443
rect 1213 11335 1233 11387
rect 1213 11279 1256 11335
rect 1213 11227 1233 11279
rect 1213 11171 1256 11227
rect 1213 11119 1233 11171
rect 1213 11063 1256 11119
rect 1213 11011 1233 11063
rect 1213 10955 1256 11011
rect 1213 10903 1233 10955
rect 1213 10847 1256 10903
rect 1213 10795 1233 10847
rect 1213 10739 1256 10795
rect 1213 10687 1233 10739
rect 1213 10631 1256 10687
rect 1213 10579 1233 10631
rect 1213 10523 1256 10579
rect 1213 10471 1233 10523
rect 1213 10415 1256 10471
rect 1213 10363 1233 10415
rect 1213 10307 1256 10363
rect 1213 10255 1233 10307
rect 1213 10199 1256 10255
rect 1213 10147 1233 10199
rect 1213 10091 1256 10147
rect 1213 10039 1233 10091
rect 1213 9983 1256 10039
rect 1213 9931 1233 9983
rect 1213 9875 1256 9931
rect 1213 9823 1233 9875
rect 1213 9767 1256 9823
rect 1213 9715 1233 9767
rect 1213 9659 1256 9715
rect 1213 9607 1233 9659
rect 1213 9551 1256 9607
rect 1213 9499 1233 9551
rect 1213 9443 1256 9499
rect 1213 9391 1233 9443
rect 1213 9335 1256 9391
rect 1213 9283 1233 9335
rect 1213 9227 1256 9283
rect 1213 9175 1233 9227
rect 1213 9119 1256 9175
rect 1213 9067 1233 9119
rect 1213 9011 1256 9067
rect 1213 8959 1233 9011
rect 1213 8903 1256 8959
rect 1213 8851 1233 8903
rect 1213 8795 1256 8851
rect 1213 8743 1233 8795
rect 1213 8687 1256 8743
rect 1213 8635 1233 8687
rect 1213 8579 1256 8635
rect 1213 8527 1233 8579
rect 1213 8471 1256 8527
rect 1213 8419 1233 8471
rect 1213 8363 1256 8419
rect 1213 8311 1233 8363
rect 1213 8255 1256 8311
rect 1213 8203 1233 8255
rect 1213 8147 1256 8203
rect 1213 8095 1233 8147
rect 1213 8039 1256 8095
rect 1213 7987 1233 8039
rect 1213 7931 1256 7987
rect 1213 7879 1233 7931
rect 1213 7823 1256 7879
rect 1213 7771 1233 7823
rect 1213 7715 1256 7771
rect 1213 7663 1233 7715
rect 1213 7607 1256 7663
rect 1213 7555 1233 7607
rect 1213 7499 1256 7555
rect 1213 7447 1233 7499
rect 1213 7418 1256 7447
rect 1402 7418 1413 12064
rect 11549 12091 11569 12143
rect 11621 12091 11677 12143
rect 11729 12091 11749 12143
rect 11549 12064 11749 12091
rect 1481 11963 11481 11975
rect 1481 11911 1493 11963
rect 1545 11960 1601 11963
rect 1653 11960 3863 11963
rect 3915 11960 3971 11963
rect 4023 11960 6239 11963
rect 6291 11960 6347 11963
rect 6399 11960 6455 11963
rect 6507 11960 6563 11963
rect 6615 11960 6671 11963
rect 6723 11960 8939 11963
rect 8991 11960 9047 11963
rect 9099 11960 11309 11963
rect 11361 11960 11417 11963
rect 1545 11911 1601 11914
rect 1653 11911 3863 11914
rect 3915 11911 3971 11914
rect 4023 11911 6239 11914
rect 6291 11911 6347 11914
rect 6399 11911 6455 11914
rect 6507 11911 6563 11914
rect 6615 11911 6671 11914
rect 6723 11911 8939 11914
rect 8991 11911 9047 11914
rect 9099 11911 11309 11914
rect 11361 11911 11417 11914
rect 11469 11911 11481 11963
rect 1481 11899 11481 11911
rect 1481 11719 11481 11731
rect 1481 11716 1760 11719
rect 1812 11716 1868 11719
rect 1920 11716 1976 11719
rect 2028 11716 2084 11719
rect 2136 11716 2192 11719
rect 2244 11716 2300 11719
rect 2352 11716 2408 11719
rect 2460 11716 2516 11719
rect 2568 11716 2624 11719
rect 2676 11716 2732 11719
rect 2784 11716 2840 11719
rect 2892 11716 2948 11719
rect 3000 11716 3056 11719
rect 3108 11716 3164 11719
rect 3216 11716 3272 11719
rect 3324 11716 3380 11719
rect 3432 11716 3488 11719
rect 3540 11716 3596 11719
rect 3648 11716 3704 11719
rect 3756 11716 4130 11719
rect 4182 11716 4238 11719
rect 4290 11716 4346 11719
rect 4398 11716 4454 11719
rect 4506 11716 4562 11719
rect 4614 11716 4670 11719
rect 4722 11716 4778 11719
rect 4830 11716 4886 11719
rect 4938 11716 4994 11719
rect 5046 11716 5102 11719
rect 5154 11716 5210 11719
rect 5262 11716 5318 11719
rect 5370 11716 5426 11719
rect 5478 11716 5534 11719
rect 5586 11716 5642 11719
rect 5694 11716 5750 11719
rect 5802 11716 5858 11719
rect 5910 11716 5966 11719
rect 6018 11716 6074 11719
rect 6126 11716 6836 11719
rect 6888 11716 6944 11719
rect 6996 11716 7052 11719
rect 7104 11716 7160 11719
rect 7212 11716 7268 11719
rect 7320 11716 7376 11719
rect 7428 11716 7484 11719
rect 7536 11716 7592 11719
rect 7644 11716 7700 11719
rect 7752 11716 7808 11719
rect 7860 11716 7916 11719
rect 7968 11716 8024 11719
rect 8076 11716 8132 11719
rect 8184 11716 8240 11719
rect 8292 11716 8348 11719
rect 8400 11716 8456 11719
rect 8508 11716 8564 11719
rect 8616 11716 8672 11719
rect 8724 11716 8780 11719
rect 8832 11716 9206 11719
rect 9258 11716 9314 11719
rect 9366 11716 9422 11719
rect 9474 11716 9530 11719
rect 9582 11716 9638 11719
rect 9690 11716 9746 11719
rect 9798 11716 9854 11719
rect 9906 11716 9962 11719
rect 10014 11716 10070 11719
rect 10122 11716 10178 11719
rect 10230 11716 10286 11719
rect 10338 11716 10394 11719
rect 10446 11716 10502 11719
rect 10554 11716 10610 11719
rect 10662 11716 10718 11719
rect 10770 11716 10826 11719
rect 10878 11716 10934 11719
rect 10986 11716 11042 11719
rect 11094 11716 11150 11719
rect 11202 11716 11481 11719
rect 1481 11670 1494 11716
rect 11468 11670 11481 11716
rect 1481 11667 1760 11670
rect 1812 11667 1868 11670
rect 1920 11667 1976 11670
rect 2028 11667 2084 11670
rect 2136 11667 2192 11670
rect 2244 11667 2300 11670
rect 2352 11667 2408 11670
rect 2460 11667 2516 11670
rect 2568 11667 2624 11670
rect 2676 11667 2732 11670
rect 2784 11667 2840 11670
rect 2892 11667 2948 11670
rect 3000 11667 3056 11670
rect 3108 11667 3164 11670
rect 3216 11667 3272 11670
rect 3324 11667 3380 11670
rect 3432 11667 3488 11670
rect 3540 11667 3596 11670
rect 3648 11667 3704 11670
rect 3756 11667 4130 11670
rect 4182 11667 4238 11670
rect 4290 11667 4346 11670
rect 4398 11667 4454 11670
rect 4506 11667 4562 11670
rect 4614 11667 4670 11670
rect 4722 11667 4778 11670
rect 4830 11667 4886 11670
rect 4938 11667 4994 11670
rect 5046 11667 5102 11670
rect 5154 11667 5210 11670
rect 5262 11667 5318 11670
rect 5370 11667 5426 11670
rect 5478 11667 5534 11670
rect 5586 11667 5642 11670
rect 5694 11667 5750 11670
rect 5802 11667 5858 11670
rect 5910 11667 5966 11670
rect 6018 11667 6074 11670
rect 6126 11667 6836 11670
rect 6888 11667 6944 11670
rect 6996 11667 7052 11670
rect 7104 11667 7160 11670
rect 7212 11667 7268 11670
rect 7320 11667 7376 11670
rect 7428 11667 7484 11670
rect 7536 11667 7592 11670
rect 7644 11667 7700 11670
rect 7752 11667 7808 11670
rect 7860 11667 7916 11670
rect 7968 11667 8024 11670
rect 8076 11667 8132 11670
rect 8184 11667 8240 11670
rect 8292 11667 8348 11670
rect 8400 11667 8456 11670
rect 8508 11667 8564 11670
rect 8616 11667 8672 11670
rect 8724 11667 8780 11670
rect 8832 11667 9206 11670
rect 9258 11667 9314 11670
rect 9366 11667 9422 11670
rect 9474 11667 9530 11670
rect 9582 11667 9638 11670
rect 9690 11667 9746 11670
rect 9798 11667 9854 11670
rect 9906 11667 9962 11670
rect 10014 11667 10070 11670
rect 10122 11667 10178 11670
rect 10230 11667 10286 11670
rect 10338 11667 10394 11670
rect 10446 11667 10502 11670
rect 10554 11667 10610 11670
rect 10662 11667 10718 11670
rect 10770 11667 10826 11670
rect 10878 11667 10934 11670
rect 10986 11667 11042 11670
rect 11094 11667 11150 11670
rect 11202 11667 11481 11670
rect 1481 11655 11481 11667
rect 1481 11475 11481 11487
rect 1481 11423 1493 11475
rect 1545 11472 1601 11475
rect 1653 11472 3863 11475
rect 3915 11472 3971 11475
rect 4023 11472 6239 11475
rect 6291 11472 6347 11475
rect 6399 11472 6455 11475
rect 6507 11472 6563 11475
rect 6615 11472 6671 11475
rect 6723 11472 8939 11475
rect 8991 11472 9047 11475
rect 9099 11472 11309 11475
rect 11361 11472 11417 11475
rect 1545 11423 1601 11426
rect 1653 11423 3863 11426
rect 3915 11423 3971 11426
rect 4023 11423 6239 11426
rect 6291 11423 6347 11426
rect 6399 11423 6455 11426
rect 6507 11423 6563 11426
rect 6615 11423 6671 11426
rect 6723 11423 8939 11426
rect 8991 11423 9047 11426
rect 9099 11423 11309 11426
rect 11361 11423 11417 11426
rect 11469 11423 11481 11475
rect 1481 11411 11481 11423
rect 1481 11231 11481 11243
rect 1481 11228 1760 11231
rect 1812 11228 1868 11231
rect 1920 11228 1976 11231
rect 2028 11228 2084 11231
rect 2136 11228 2192 11231
rect 2244 11228 2300 11231
rect 2352 11228 2408 11231
rect 2460 11228 2516 11231
rect 2568 11228 2624 11231
rect 2676 11228 2732 11231
rect 2784 11228 2840 11231
rect 2892 11228 2948 11231
rect 3000 11228 3056 11231
rect 3108 11228 3164 11231
rect 3216 11228 3272 11231
rect 3324 11228 3380 11231
rect 3432 11228 3488 11231
rect 3540 11228 3596 11231
rect 3648 11228 3704 11231
rect 3756 11228 4130 11231
rect 4182 11228 4238 11231
rect 4290 11228 4346 11231
rect 4398 11228 4454 11231
rect 4506 11228 4562 11231
rect 4614 11228 4670 11231
rect 4722 11228 4778 11231
rect 4830 11228 4886 11231
rect 4938 11228 4994 11231
rect 5046 11228 5102 11231
rect 5154 11228 5210 11231
rect 5262 11228 5318 11231
rect 5370 11228 5426 11231
rect 5478 11228 5534 11231
rect 5586 11228 5642 11231
rect 5694 11228 5750 11231
rect 5802 11228 5858 11231
rect 5910 11228 5966 11231
rect 6018 11228 6074 11231
rect 6126 11228 6836 11231
rect 6888 11228 6944 11231
rect 6996 11228 7052 11231
rect 7104 11228 7160 11231
rect 7212 11228 7268 11231
rect 7320 11228 7376 11231
rect 7428 11228 7484 11231
rect 7536 11228 7592 11231
rect 7644 11228 7700 11231
rect 7752 11228 7808 11231
rect 7860 11228 7916 11231
rect 7968 11228 8024 11231
rect 8076 11228 8132 11231
rect 8184 11228 8240 11231
rect 8292 11228 8348 11231
rect 8400 11228 8456 11231
rect 8508 11228 8564 11231
rect 8616 11228 8672 11231
rect 8724 11228 8780 11231
rect 8832 11228 9206 11231
rect 9258 11228 9314 11231
rect 9366 11228 9422 11231
rect 9474 11228 9530 11231
rect 9582 11228 9638 11231
rect 9690 11228 9746 11231
rect 9798 11228 9854 11231
rect 9906 11228 9962 11231
rect 10014 11228 10070 11231
rect 10122 11228 10178 11231
rect 10230 11228 10286 11231
rect 10338 11228 10394 11231
rect 10446 11228 10502 11231
rect 10554 11228 10610 11231
rect 10662 11228 10718 11231
rect 10770 11228 10826 11231
rect 10878 11228 10934 11231
rect 10986 11228 11042 11231
rect 11094 11228 11150 11231
rect 11202 11228 11481 11231
rect 1481 11182 1494 11228
rect 11468 11182 11481 11228
rect 1481 11179 1760 11182
rect 1812 11179 1868 11182
rect 1920 11179 1976 11182
rect 2028 11179 2084 11182
rect 2136 11179 2192 11182
rect 2244 11179 2300 11182
rect 2352 11179 2408 11182
rect 2460 11179 2516 11182
rect 2568 11179 2624 11182
rect 2676 11179 2732 11182
rect 2784 11179 2840 11182
rect 2892 11179 2948 11182
rect 3000 11179 3056 11182
rect 3108 11179 3164 11182
rect 3216 11179 3272 11182
rect 3324 11179 3380 11182
rect 3432 11179 3488 11182
rect 3540 11179 3596 11182
rect 3648 11179 3704 11182
rect 3756 11179 4130 11182
rect 4182 11179 4238 11182
rect 4290 11179 4346 11182
rect 4398 11179 4454 11182
rect 4506 11179 4562 11182
rect 4614 11179 4670 11182
rect 4722 11179 4778 11182
rect 4830 11179 4886 11182
rect 4938 11179 4994 11182
rect 5046 11179 5102 11182
rect 5154 11179 5210 11182
rect 5262 11179 5318 11182
rect 5370 11179 5426 11182
rect 5478 11179 5534 11182
rect 5586 11179 5642 11182
rect 5694 11179 5750 11182
rect 5802 11179 5858 11182
rect 5910 11179 5966 11182
rect 6018 11179 6074 11182
rect 6126 11179 6836 11182
rect 6888 11179 6944 11182
rect 6996 11179 7052 11182
rect 7104 11179 7160 11182
rect 7212 11179 7268 11182
rect 7320 11179 7376 11182
rect 7428 11179 7484 11182
rect 7536 11179 7592 11182
rect 7644 11179 7700 11182
rect 7752 11179 7808 11182
rect 7860 11179 7916 11182
rect 7968 11179 8024 11182
rect 8076 11179 8132 11182
rect 8184 11179 8240 11182
rect 8292 11179 8348 11182
rect 8400 11179 8456 11182
rect 8508 11179 8564 11182
rect 8616 11179 8672 11182
rect 8724 11179 8780 11182
rect 8832 11179 9206 11182
rect 9258 11179 9314 11182
rect 9366 11179 9422 11182
rect 9474 11179 9530 11182
rect 9582 11179 9638 11182
rect 9690 11179 9746 11182
rect 9798 11179 9854 11182
rect 9906 11179 9962 11182
rect 10014 11179 10070 11182
rect 10122 11179 10178 11182
rect 10230 11179 10286 11182
rect 10338 11179 10394 11182
rect 10446 11179 10502 11182
rect 10554 11179 10610 11182
rect 10662 11179 10718 11182
rect 10770 11179 10826 11182
rect 10878 11179 10934 11182
rect 10986 11179 11042 11182
rect 11094 11179 11150 11182
rect 11202 11179 11481 11182
rect 1481 11167 11481 11179
rect 1481 10987 11481 10999
rect 1481 10935 1493 10987
rect 1545 10984 1601 10987
rect 1653 10984 3863 10987
rect 3915 10984 3971 10987
rect 4023 10984 6239 10987
rect 6291 10984 6347 10987
rect 6399 10984 6455 10987
rect 6507 10984 6563 10987
rect 6615 10984 6671 10987
rect 6723 10984 8939 10987
rect 8991 10984 9047 10987
rect 9099 10984 11309 10987
rect 11361 10984 11417 10987
rect 1545 10935 1601 10938
rect 1653 10935 3863 10938
rect 3915 10935 3971 10938
rect 4023 10935 6239 10938
rect 6291 10935 6347 10938
rect 6399 10935 6455 10938
rect 6507 10935 6563 10938
rect 6615 10935 6671 10938
rect 6723 10935 8939 10938
rect 8991 10935 9047 10938
rect 9099 10935 11309 10938
rect 11361 10935 11417 10938
rect 11469 10935 11481 10987
rect 1481 10923 11481 10935
rect 1481 10743 11481 10755
rect 1481 10740 1760 10743
rect 1812 10740 1868 10743
rect 1920 10740 1976 10743
rect 2028 10740 2084 10743
rect 2136 10740 2192 10743
rect 2244 10740 2300 10743
rect 2352 10740 2408 10743
rect 2460 10740 2516 10743
rect 2568 10740 2624 10743
rect 2676 10740 2732 10743
rect 2784 10740 2840 10743
rect 2892 10740 2948 10743
rect 3000 10740 3056 10743
rect 3108 10740 3164 10743
rect 3216 10740 3272 10743
rect 3324 10740 3380 10743
rect 3432 10740 3488 10743
rect 3540 10740 3596 10743
rect 3648 10740 3704 10743
rect 3756 10740 4130 10743
rect 4182 10740 4238 10743
rect 4290 10740 4346 10743
rect 4398 10740 4454 10743
rect 4506 10740 4562 10743
rect 4614 10740 4670 10743
rect 4722 10740 4778 10743
rect 4830 10740 4886 10743
rect 4938 10740 4994 10743
rect 5046 10740 5102 10743
rect 5154 10740 5210 10743
rect 5262 10740 5318 10743
rect 5370 10740 5426 10743
rect 5478 10740 5534 10743
rect 5586 10740 5642 10743
rect 5694 10740 5750 10743
rect 5802 10740 5858 10743
rect 5910 10740 5966 10743
rect 6018 10740 6074 10743
rect 6126 10740 6836 10743
rect 6888 10740 6944 10743
rect 6996 10740 7052 10743
rect 7104 10740 7160 10743
rect 7212 10740 7268 10743
rect 7320 10740 7376 10743
rect 7428 10740 7484 10743
rect 7536 10740 7592 10743
rect 7644 10740 7700 10743
rect 7752 10740 7808 10743
rect 7860 10740 7916 10743
rect 7968 10740 8024 10743
rect 8076 10740 8132 10743
rect 8184 10740 8240 10743
rect 8292 10740 8348 10743
rect 8400 10740 8456 10743
rect 8508 10740 8564 10743
rect 8616 10740 8672 10743
rect 8724 10740 8780 10743
rect 8832 10740 9206 10743
rect 9258 10740 9314 10743
rect 9366 10740 9422 10743
rect 9474 10740 9530 10743
rect 9582 10740 9638 10743
rect 9690 10740 9746 10743
rect 9798 10740 9854 10743
rect 9906 10740 9962 10743
rect 10014 10740 10070 10743
rect 10122 10740 10178 10743
rect 10230 10740 10286 10743
rect 10338 10740 10394 10743
rect 10446 10740 10502 10743
rect 10554 10740 10610 10743
rect 10662 10740 10718 10743
rect 10770 10740 10826 10743
rect 10878 10740 10934 10743
rect 10986 10740 11042 10743
rect 11094 10740 11150 10743
rect 11202 10740 11481 10743
rect 1481 10694 1494 10740
rect 11468 10694 11481 10740
rect 1481 10691 1760 10694
rect 1812 10691 1868 10694
rect 1920 10691 1976 10694
rect 2028 10691 2084 10694
rect 2136 10691 2192 10694
rect 2244 10691 2300 10694
rect 2352 10691 2408 10694
rect 2460 10691 2516 10694
rect 2568 10691 2624 10694
rect 2676 10691 2732 10694
rect 2784 10691 2840 10694
rect 2892 10691 2948 10694
rect 3000 10691 3056 10694
rect 3108 10691 3164 10694
rect 3216 10691 3272 10694
rect 3324 10691 3380 10694
rect 3432 10691 3488 10694
rect 3540 10691 3596 10694
rect 3648 10691 3704 10694
rect 3756 10691 4130 10694
rect 4182 10691 4238 10694
rect 4290 10691 4346 10694
rect 4398 10691 4454 10694
rect 4506 10691 4562 10694
rect 4614 10691 4670 10694
rect 4722 10691 4778 10694
rect 4830 10691 4886 10694
rect 4938 10691 4994 10694
rect 5046 10691 5102 10694
rect 5154 10691 5210 10694
rect 5262 10691 5318 10694
rect 5370 10691 5426 10694
rect 5478 10691 5534 10694
rect 5586 10691 5642 10694
rect 5694 10691 5750 10694
rect 5802 10691 5858 10694
rect 5910 10691 5966 10694
rect 6018 10691 6074 10694
rect 6126 10691 6836 10694
rect 6888 10691 6944 10694
rect 6996 10691 7052 10694
rect 7104 10691 7160 10694
rect 7212 10691 7268 10694
rect 7320 10691 7376 10694
rect 7428 10691 7484 10694
rect 7536 10691 7592 10694
rect 7644 10691 7700 10694
rect 7752 10691 7808 10694
rect 7860 10691 7916 10694
rect 7968 10691 8024 10694
rect 8076 10691 8132 10694
rect 8184 10691 8240 10694
rect 8292 10691 8348 10694
rect 8400 10691 8456 10694
rect 8508 10691 8564 10694
rect 8616 10691 8672 10694
rect 8724 10691 8780 10694
rect 8832 10691 9206 10694
rect 9258 10691 9314 10694
rect 9366 10691 9422 10694
rect 9474 10691 9530 10694
rect 9582 10691 9638 10694
rect 9690 10691 9746 10694
rect 9798 10691 9854 10694
rect 9906 10691 9962 10694
rect 10014 10691 10070 10694
rect 10122 10691 10178 10694
rect 10230 10691 10286 10694
rect 10338 10691 10394 10694
rect 10446 10691 10502 10694
rect 10554 10691 10610 10694
rect 10662 10691 10718 10694
rect 10770 10691 10826 10694
rect 10878 10691 10934 10694
rect 10986 10691 11042 10694
rect 11094 10691 11150 10694
rect 11202 10691 11481 10694
rect 1481 10679 11481 10691
rect 1481 10499 11481 10511
rect 1481 10447 1493 10499
rect 1545 10496 1601 10499
rect 1653 10496 3863 10499
rect 3915 10496 3971 10499
rect 4023 10496 6239 10499
rect 6291 10496 6347 10499
rect 6399 10496 6455 10499
rect 6507 10496 6563 10499
rect 6615 10496 6671 10499
rect 6723 10496 8939 10499
rect 8991 10496 9047 10499
rect 9099 10496 11309 10499
rect 11361 10496 11417 10499
rect 1545 10447 1601 10450
rect 1653 10447 3863 10450
rect 3915 10447 3971 10450
rect 4023 10447 6239 10450
rect 6291 10447 6347 10450
rect 6399 10447 6455 10450
rect 6507 10447 6563 10450
rect 6615 10447 6671 10450
rect 6723 10447 8939 10450
rect 8991 10447 9047 10450
rect 9099 10447 11309 10450
rect 11361 10447 11417 10450
rect 11469 10447 11481 10499
rect 1481 10435 11481 10447
rect 1481 10255 11481 10267
rect 1481 10252 1760 10255
rect 1812 10252 1868 10255
rect 1920 10252 1976 10255
rect 2028 10252 2084 10255
rect 2136 10252 2192 10255
rect 2244 10252 2300 10255
rect 2352 10252 2408 10255
rect 2460 10252 2516 10255
rect 2568 10252 2624 10255
rect 2676 10252 2732 10255
rect 2784 10252 2840 10255
rect 2892 10252 2948 10255
rect 3000 10252 3056 10255
rect 3108 10252 3164 10255
rect 3216 10252 3272 10255
rect 3324 10252 3380 10255
rect 3432 10252 3488 10255
rect 3540 10252 3596 10255
rect 3648 10252 3704 10255
rect 3756 10252 4130 10255
rect 4182 10252 4238 10255
rect 4290 10252 4346 10255
rect 4398 10252 4454 10255
rect 4506 10252 4562 10255
rect 4614 10252 4670 10255
rect 4722 10252 4778 10255
rect 4830 10252 4886 10255
rect 4938 10252 4994 10255
rect 5046 10252 5102 10255
rect 5154 10252 5210 10255
rect 5262 10252 5318 10255
rect 5370 10252 5426 10255
rect 5478 10252 5534 10255
rect 5586 10252 5642 10255
rect 5694 10252 5750 10255
rect 5802 10252 5858 10255
rect 5910 10252 5966 10255
rect 6018 10252 6074 10255
rect 6126 10252 6836 10255
rect 6888 10252 6944 10255
rect 6996 10252 7052 10255
rect 7104 10252 7160 10255
rect 7212 10252 7268 10255
rect 7320 10252 7376 10255
rect 7428 10252 7484 10255
rect 7536 10252 7592 10255
rect 7644 10252 7700 10255
rect 7752 10252 7808 10255
rect 7860 10252 7916 10255
rect 7968 10252 8024 10255
rect 8076 10252 8132 10255
rect 8184 10252 8240 10255
rect 8292 10252 8348 10255
rect 8400 10252 8456 10255
rect 8508 10252 8564 10255
rect 8616 10252 8672 10255
rect 8724 10252 8780 10255
rect 8832 10252 9206 10255
rect 9258 10252 9314 10255
rect 9366 10252 9422 10255
rect 9474 10252 9530 10255
rect 9582 10252 9638 10255
rect 9690 10252 9746 10255
rect 9798 10252 9854 10255
rect 9906 10252 9962 10255
rect 10014 10252 10070 10255
rect 10122 10252 10178 10255
rect 10230 10252 10286 10255
rect 10338 10252 10394 10255
rect 10446 10252 10502 10255
rect 10554 10252 10610 10255
rect 10662 10252 10718 10255
rect 10770 10252 10826 10255
rect 10878 10252 10934 10255
rect 10986 10252 11042 10255
rect 11094 10252 11150 10255
rect 11202 10252 11481 10255
rect 1481 10206 1494 10252
rect 11468 10206 11481 10252
rect 1481 10203 1760 10206
rect 1812 10203 1868 10206
rect 1920 10203 1976 10206
rect 2028 10203 2084 10206
rect 2136 10203 2192 10206
rect 2244 10203 2300 10206
rect 2352 10203 2408 10206
rect 2460 10203 2516 10206
rect 2568 10203 2624 10206
rect 2676 10203 2732 10206
rect 2784 10203 2840 10206
rect 2892 10203 2948 10206
rect 3000 10203 3056 10206
rect 3108 10203 3164 10206
rect 3216 10203 3272 10206
rect 3324 10203 3380 10206
rect 3432 10203 3488 10206
rect 3540 10203 3596 10206
rect 3648 10203 3704 10206
rect 3756 10203 4130 10206
rect 4182 10203 4238 10206
rect 4290 10203 4346 10206
rect 4398 10203 4454 10206
rect 4506 10203 4562 10206
rect 4614 10203 4670 10206
rect 4722 10203 4778 10206
rect 4830 10203 4886 10206
rect 4938 10203 4994 10206
rect 5046 10203 5102 10206
rect 5154 10203 5210 10206
rect 5262 10203 5318 10206
rect 5370 10203 5426 10206
rect 5478 10203 5534 10206
rect 5586 10203 5642 10206
rect 5694 10203 5750 10206
rect 5802 10203 5858 10206
rect 5910 10203 5966 10206
rect 6018 10203 6074 10206
rect 6126 10203 6836 10206
rect 6888 10203 6944 10206
rect 6996 10203 7052 10206
rect 7104 10203 7160 10206
rect 7212 10203 7268 10206
rect 7320 10203 7376 10206
rect 7428 10203 7484 10206
rect 7536 10203 7592 10206
rect 7644 10203 7700 10206
rect 7752 10203 7808 10206
rect 7860 10203 7916 10206
rect 7968 10203 8024 10206
rect 8076 10203 8132 10206
rect 8184 10203 8240 10206
rect 8292 10203 8348 10206
rect 8400 10203 8456 10206
rect 8508 10203 8564 10206
rect 8616 10203 8672 10206
rect 8724 10203 8780 10206
rect 8832 10203 9206 10206
rect 9258 10203 9314 10206
rect 9366 10203 9422 10206
rect 9474 10203 9530 10206
rect 9582 10203 9638 10206
rect 9690 10203 9746 10206
rect 9798 10203 9854 10206
rect 9906 10203 9962 10206
rect 10014 10203 10070 10206
rect 10122 10203 10178 10206
rect 10230 10203 10286 10206
rect 10338 10203 10394 10206
rect 10446 10203 10502 10206
rect 10554 10203 10610 10206
rect 10662 10203 10718 10206
rect 10770 10203 10826 10206
rect 10878 10203 10934 10206
rect 10986 10203 11042 10206
rect 11094 10203 11150 10206
rect 11202 10203 11481 10206
rect 1481 10191 11481 10203
rect 1481 10011 11481 10023
rect 1481 9959 1493 10011
rect 1545 10008 1601 10011
rect 1653 10008 3863 10011
rect 3915 10008 3971 10011
rect 4023 10008 6239 10011
rect 6291 10008 6347 10011
rect 6399 10008 6455 10011
rect 6507 10008 6563 10011
rect 6615 10008 6671 10011
rect 6723 10008 8939 10011
rect 8991 10008 9047 10011
rect 9099 10008 11309 10011
rect 11361 10008 11417 10011
rect 1545 9959 1601 9962
rect 1653 9959 3863 9962
rect 3915 9959 3971 9962
rect 4023 9959 6239 9962
rect 6291 9959 6347 9962
rect 6399 9959 6455 9962
rect 6507 9959 6563 9962
rect 6615 9959 6671 9962
rect 6723 9959 8939 9962
rect 8991 9959 9047 9962
rect 9099 9959 11309 9962
rect 11361 9959 11417 9962
rect 11469 9959 11481 10011
rect 1481 9947 11481 9959
rect 1481 9767 11481 9779
rect 1481 9764 1760 9767
rect 1812 9764 1868 9767
rect 1920 9764 1976 9767
rect 2028 9764 2084 9767
rect 2136 9764 2192 9767
rect 2244 9764 2300 9767
rect 2352 9764 2408 9767
rect 2460 9764 2516 9767
rect 2568 9764 2624 9767
rect 2676 9764 2732 9767
rect 2784 9764 2840 9767
rect 2892 9764 2948 9767
rect 3000 9764 3056 9767
rect 3108 9764 3164 9767
rect 3216 9764 3272 9767
rect 3324 9764 3380 9767
rect 3432 9764 3488 9767
rect 3540 9764 3596 9767
rect 3648 9764 3704 9767
rect 3756 9764 4130 9767
rect 4182 9764 4238 9767
rect 4290 9764 4346 9767
rect 4398 9764 4454 9767
rect 4506 9764 4562 9767
rect 4614 9764 4670 9767
rect 4722 9764 4778 9767
rect 4830 9764 4886 9767
rect 4938 9764 4994 9767
rect 5046 9764 5102 9767
rect 5154 9764 5210 9767
rect 5262 9764 5318 9767
rect 5370 9764 5426 9767
rect 5478 9764 5534 9767
rect 5586 9764 5642 9767
rect 5694 9764 5750 9767
rect 5802 9764 5858 9767
rect 5910 9764 5966 9767
rect 6018 9764 6074 9767
rect 6126 9764 6836 9767
rect 6888 9764 6944 9767
rect 6996 9764 7052 9767
rect 7104 9764 7160 9767
rect 7212 9764 7268 9767
rect 7320 9764 7376 9767
rect 7428 9764 7484 9767
rect 7536 9764 7592 9767
rect 7644 9764 7700 9767
rect 7752 9764 7808 9767
rect 7860 9764 7916 9767
rect 7968 9764 8024 9767
rect 8076 9764 8132 9767
rect 8184 9764 8240 9767
rect 8292 9764 8348 9767
rect 8400 9764 8456 9767
rect 8508 9764 8564 9767
rect 8616 9764 8672 9767
rect 8724 9764 8780 9767
rect 8832 9764 9206 9767
rect 9258 9764 9314 9767
rect 9366 9764 9422 9767
rect 9474 9764 9530 9767
rect 9582 9764 9638 9767
rect 9690 9764 9746 9767
rect 9798 9764 9854 9767
rect 9906 9764 9962 9767
rect 10014 9764 10070 9767
rect 10122 9764 10178 9767
rect 10230 9764 10286 9767
rect 10338 9764 10394 9767
rect 10446 9764 10502 9767
rect 10554 9764 10610 9767
rect 10662 9764 10718 9767
rect 10770 9764 10826 9767
rect 10878 9764 10934 9767
rect 10986 9764 11042 9767
rect 11094 9764 11150 9767
rect 11202 9764 11481 9767
rect 1481 9718 1494 9764
rect 11468 9718 11481 9764
rect 1481 9715 1760 9718
rect 1812 9715 1868 9718
rect 1920 9715 1976 9718
rect 2028 9715 2084 9718
rect 2136 9715 2192 9718
rect 2244 9715 2300 9718
rect 2352 9715 2408 9718
rect 2460 9715 2516 9718
rect 2568 9715 2624 9718
rect 2676 9715 2732 9718
rect 2784 9715 2840 9718
rect 2892 9715 2948 9718
rect 3000 9715 3056 9718
rect 3108 9715 3164 9718
rect 3216 9715 3272 9718
rect 3324 9715 3380 9718
rect 3432 9715 3488 9718
rect 3540 9715 3596 9718
rect 3648 9715 3704 9718
rect 3756 9715 4130 9718
rect 4182 9715 4238 9718
rect 4290 9715 4346 9718
rect 4398 9715 4454 9718
rect 4506 9715 4562 9718
rect 4614 9715 4670 9718
rect 4722 9715 4778 9718
rect 4830 9715 4886 9718
rect 4938 9715 4994 9718
rect 5046 9715 5102 9718
rect 5154 9715 5210 9718
rect 5262 9715 5318 9718
rect 5370 9715 5426 9718
rect 5478 9715 5534 9718
rect 5586 9715 5642 9718
rect 5694 9715 5750 9718
rect 5802 9715 5858 9718
rect 5910 9715 5966 9718
rect 6018 9715 6074 9718
rect 6126 9715 6836 9718
rect 6888 9715 6944 9718
rect 6996 9715 7052 9718
rect 7104 9715 7160 9718
rect 7212 9715 7268 9718
rect 7320 9715 7376 9718
rect 7428 9715 7484 9718
rect 7536 9715 7592 9718
rect 7644 9715 7700 9718
rect 7752 9715 7808 9718
rect 7860 9715 7916 9718
rect 7968 9715 8024 9718
rect 8076 9715 8132 9718
rect 8184 9715 8240 9718
rect 8292 9715 8348 9718
rect 8400 9715 8456 9718
rect 8508 9715 8564 9718
rect 8616 9715 8672 9718
rect 8724 9715 8780 9718
rect 8832 9715 9206 9718
rect 9258 9715 9314 9718
rect 9366 9715 9422 9718
rect 9474 9715 9530 9718
rect 9582 9715 9638 9718
rect 9690 9715 9746 9718
rect 9798 9715 9854 9718
rect 9906 9715 9962 9718
rect 10014 9715 10070 9718
rect 10122 9715 10178 9718
rect 10230 9715 10286 9718
rect 10338 9715 10394 9718
rect 10446 9715 10502 9718
rect 10554 9715 10610 9718
rect 10662 9715 10718 9718
rect 10770 9715 10826 9718
rect 10878 9715 10934 9718
rect 10986 9715 11042 9718
rect 11094 9715 11150 9718
rect 11202 9715 11481 9718
rect 1481 9703 11481 9715
rect 1481 9523 11481 9535
rect 1481 9471 1493 9523
rect 1545 9520 1601 9523
rect 1653 9520 3863 9523
rect 3915 9520 3971 9523
rect 4023 9520 6239 9523
rect 6291 9520 6347 9523
rect 6399 9520 6455 9523
rect 6507 9520 6563 9523
rect 6615 9520 6671 9523
rect 6723 9520 8939 9523
rect 8991 9520 9047 9523
rect 9099 9520 11309 9523
rect 11361 9520 11417 9523
rect 1545 9471 1601 9474
rect 1653 9471 3863 9474
rect 3915 9471 3971 9474
rect 4023 9471 6239 9474
rect 6291 9471 6347 9474
rect 6399 9471 6455 9474
rect 6507 9471 6563 9474
rect 6615 9471 6671 9474
rect 6723 9471 8939 9474
rect 8991 9471 9047 9474
rect 9099 9471 11309 9474
rect 11361 9471 11417 9474
rect 11469 9471 11481 9523
rect 1481 9459 11481 9471
rect 1481 9279 11481 9291
rect 1481 9276 1760 9279
rect 1812 9276 1868 9279
rect 1920 9276 1976 9279
rect 2028 9276 2084 9279
rect 2136 9276 2192 9279
rect 2244 9276 2300 9279
rect 2352 9276 2408 9279
rect 2460 9276 2516 9279
rect 2568 9276 2624 9279
rect 2676 9276 2732 9279
rect 2784 9276 2840 9279
rect 2892 9276 2948 9279
rect 3000 9276 3056 9279
rect 3108 9276 3164 9279
rect 3216 9276 3272 9279
rect 3324 9276 3380 9279
rect 3432 9276 3488 9279
rect 3540 9276 3596 9279
rect 3648 9276 3704 9279
rect 3756 9276 4130 9279
rect 4182 9276 4238 9279
rect 4290 9276 4346 9279
rect 4398 9276 4454 9279
rect 4506 9276 4562 9279
rect 4614 9276 4670 9279
rect 4722 9276 4778 9279
rect 4830 9276 4886 9279
rect 4938 9276 4994 9279
rect 5046 9276 5102 9279
rect 5154 9276 5210 9279
rect 5262 9276 5318 9279
rect 5370 9276 5426 9279
rect 5478 9276 5534 9279
rect 5586 9276 5642 9279
rect 5694 9276 5750 9279
rect 5802 9276 5858 9279
rect 5910 9276 5966 9279
rect 6018 9276 6074 9279
rect 6126 9276 6836 9279
rect 6888 9276 6944 9279
rect 6996 9276 7052 9279
rect 7104 9276 7160 9279
rect 7212 9276 7268 9279
rect 7320 9276 7376 9279
rect 7428 9276 7484 9279
rect 7536 9276 7592 9279
rect 7644 9276 7700 9279
rect 7752 9276 7808 9279
rect 7860 9276 7916 9279
rect 7968 9276 8024 9279
rect 8076 9276 8132 9279
rect 8184 9276 8240 9279
rect 8292 9276 8348 9279
rect 8400 9276 8456 9279
rect 8508 9276 8564 9279
rect 8616 9276 8672 9279
rect 8724 9276 8780 9279
rect 8832 9276 9206 9279
rect 9258 9276 9314 9279
rect 9366 9276 9422 9279
rect 9474 9276 9530 9279
rect 9582 9276 9638 9279
rect 9690 9276 9746 9279
rect 9798 9276 9854 9279
rect 9906 9276 9962 9279
rect 10014 9276 10070 9279
rect 10122 9276 10178 9279
rect 10230 9276 10286 9279
rect 10338 9276 10394 9279
rect 10446 9276 10502 9279
rect 10554 9276 10610 9279
rect 10662 9276 10718 9279
rect 10770 9276 10826 9279
rect 10878 9276 10934 9279
rect 10986 9276 11042 9279
rect 11094 9276 11150 9279
rect 11202 9276 11481 9279
rect 1481 9230 1494 9276
rect 11468 9230 11481 9276
rect 1481 9227 1760 9230
rect 1812 9227 1868 9230
rect 1920 9227 1976 9230
rect 2028 9227 2084 9230
rect 2136 9227 2192 9230
rect 2244 9227 2300 9230
rect 2352 9227 2408 9230
rect 2460 9227 2516 9230
rect 2568 9227 2624 9230
rect 2676 9227 2732 9230
rect 2784 9227 2840 9230
rect 2892 9227 2948 9230
rect 3000 9227 3056 9230
rect 3108 9227 3164 9230
rect 3216 9227 3272 9230
rect 3324 9227 3380 9230
rect 3432 9227 3488 9230
rect 3540 9227 3596 9230
rect 3648 9227 3704 9230
rect 3756 9227 4130 9230
rect 4182 9227 4238 9230
rect 4290 9227 4346 9230
rect 4398 9227 4454 9230
rect 4506 9227 4562 9230
rect 4614 9227 4670 9230
rect 4722 9227 4778 9230
rect 4830 9227 4886 9230
rect 4938 9227 4994 9230
rect 5046 9227 5102 9230
rect 5154 9227 5210 9230
rect 5262 9227 5318 9230
rect 5370 9227 5426 9230
rect 5478 9227 5534 9230
rect 5586 9227 5642 9230
rect 5694 9227 5750 9230
rect 5802 9227 5858 9230
rect 5910 9227 5966 9230
rect 6018 9227 6074 9230
rect 6126 9227 6836 9230
rect 6888 9227 6944 9230
rect 6996 9227 7052 9230
rect 7104 9227 7160 9230
rect 7212 9227 7268 9230
rect 7320 9227 7376 9230
rect 7428 9227 7484 9230
rect 7536 9227 7592 9230
rect 7644 9227 7700 9230
rect 7752 9227 7808 9230
rect 7860 9227 7916 9230
rect 7968 9227 8024 9230
rect 8076 9227 8132 9230
rect 8184 9227 8240 9230
rect 8292 9227 8348 9230
rect 8400 9227 8456 9230
rect 8508 9227 8564 9230
rect 8616 9227 8672 9230
rect 8724 9227 8780 9230
rect 8832 9227 9206 9230
rect 9258 9227 9314 9230
rect 9366 9227 9422 9230
rect 9474 9227 9530 9230
rect 9582 9227 9638 9230
rect 9690 9227 9746 9230
rect 9798 9227 9854 9230
rect 9906 9227 9962 9230
rect 10014 9227 10070 9230
rect 10122 9227 10178 9230
rect 10230 9227 10286 9230
rect 10338 9227 10394 9230
rect 10446 9227 10502 9230
rect 10554 9227 10610 9230
rect 10662 9227 10718 9230
rect 10770 9227 10826 9230
rect 10878 9227 10934 9230
rect 10986 9227 11042 9230
rect 11094 9227 11150 9230
rect 11202 9227 11481 9230
rect 1481 9215 11481 9227
rect 1481 9035 11481 9047
rect 1481 8983 1493 9035
rect 1545 9032 1601 9035
rect 1653 9032 3863 9035
rect 3915 9032 3971 9035
rect 4023 9032 6239 9035
rect 6291 9032 6347 9035
rect 6399 9032 6455 9035
rect 6507 9032 6563 9035
rect 6615 9032 6671 9035
rect 6723 9032 8939 9035
rect 8991 9032 9047 9035
rect 9099 9032 11309 9035
rect 11361 9032 11417 9035
rect 1545 8983 1601 8986
rect 1653 8983 3863 8986
rect 3915 8983 3971 8986
rect 4023 8983 6239 8986
rect 6291 8983 6347 8986
rect 6399 8983 6455 8986
rect 6507 8983 6563 8986
rect 6615 8983 6671 8986
rect 6723 8983 8939 8986
rect 8991 8983 9047 8986
rect 9099 8983 11309 8986
rect 11361 8983 11417 8986
rect 11469 8983 11481 9035
rect 1481 8971 11481 8983
rect 1481 8791 11481 8803
rect 1481 8788 1760 8791
rect 1812 8788 1868 8791
rect 1920 8788 1976 8791
rect 2028 8788 2084 8791
rect 2136 8788 2192 8791
rect 2244 8788 2300 8791
rect 2352 8788 2408 8791
rect 2460 8788 2516 8791
rect 2568 8788 2624 8791
rect 2676 8788 2732 8791
rect 2784 8788 2840 8791
rect 2892 8788 2948 8791
rect 3000 8788 3056 8791
rect 3108 8788 3164 8791
rect 3216 8788 3272 8791
rect 3324 8788 3380 8791
rect 3432 8788 3488 8791
rect 3540 8788 3596 8791
rect 3648 8788 3704 8791
rect 3756 8788 4130 8791
rect 4182 8788 4238 8791
rect 4290 8788 4346 8791
rect 4398 8788 4454 8791
rect 4506 8788 4562 8791
rect 4614 8788 4670 8791
rect 4722 8788 4778 8791
rect 4830 8788 4886 8791
rect 4938 8788 4994 8791
rect 5046 8788 5102 8791
rect 5154 8788 5210 8791
rect 5262 8788 5318 8791
rect 5370 8788 5426 8791
rect 5478 8788 5534 8791
rect 5586 8788 5642 8791
rect 5694 8788 5750 8791
rect 5802 8788 5858 8791
rect 5910 8788 5966 8791
rect 6018 8788 6074 8791
rect 6126 8788 6836 8791
rect 6888 8788 6944 8791
rect 6996 8788 7052 8791
rect 7104 8788 7160 8791
rect 7212 8788 7268 8791
rect 7320 8788 7376 8791
rect 7428 8788 7484 8791
rect 7536 8788 7592 8791
rect 7644 8788 7700 8791
rect 7752 8788 7808 8791
rect 7860 8788 7916 8791
rect 7968 8788 8024 8791
rect 8076 8788 8132 8791
rect 8184 8788 8240 8791
rect 8292 8788 8348 8791
rect 8400 8788 8456 8791
rect 8508 8788 8564 8791
rect 8616 8788 8672 8791
rect 8724 8788 8780 8791
rect 8832 8788 9206 8791
rect 9258 8788 9314 8791
rect 9366 8788 9422 8791
rect 9474 8788 9530 8791
rect 9582 8788 9638 8791
rect 9690 8788 9746 8791
rect 9798 8788 9854 8791
rect 9906 8788 9962 8791
rect 10014 8788 10070 8791
rect 10122 8788 10178 8791
rect 10230 8788 10286 8791
rect 10338 8788 10394 8791
rect 10446 8788 10502 8791
rect 10554 8788 10610 8791
rect 10662 8788 10718 8791
rect 10770 8788 10826 8791
rect 10878 8788 10934 8791
rect 10986 8788 11042 8791
rect 11094 8788 11150 8791
rect 11202 8788 11481 8791
rect 1481 8742 1494 8788
rect 11468 8742 11481 8788
rect 1481 8739 1760 8742
rect 1812 8739 1868 8742
rect 1920 8739 1976 8742
rect 2028 8739 2084 8742
rect 2136 8739 2192 8742
rect 2244 8739 2300 8742
rect 2352 8739 2408 8742
rect 2460 8739 2516 8742
rect 2568 8739 2624 8742
rect 2676 8739 2732 8742
rect 2784 8739 2840 8742
rect 2892 8739 2948 8742
rect 3000 8739 3056 8742
rect 3108 8739 3164 8742
rect 3216 8739 3272 8742
rect 3324 8739 3380 8742
rect 3432 8739 3488 8742
rect 3540 8739 3596 8742
rect 3648 8739 3704 8742
rect 3756 8739 4130 8742
rect 4182 8739 4238 8742
rect 4290 8739 4346 8742
rect 4398 8739 4454 8742
rect 4506 8739 4562 8742
rect 4614 8739 4670 8742
rect 4722 8739 4778 8742
rect 4830 8739 4886 8742
rect 4938 8739 4994 8742
rect 5046 8739 5102 8742
rect 5154 8739 5210 8742
rect 5262 8739 5318 8742
rect 5370 8739 5426 8742
rect 5478 8739 5534 8742
rect 5586 8739 5642 8742
rect 5694 8739 5750 8742
rect 5802 8739 5858 8742
rect 5910 8739 5966 8742
rect 6018 8739 6074 8742
rect 6126 8739 6836 8742
rect 6888 8739 6944 8742
rect 6996 8739 7052 8742
rect 7104 8739 7160 8742
rect 7212 8739 7268 8742
rect 7320 8739 7376 8742
rect 7428 8739 7484 8742
rect 7536 8739 7592 8742
rect 7644 8739 7700 8742
rect 7752 8739 7808 8742
rect 7860 8739 7916 8742
rect 7968 8739 8024 8742
rect 8076 8739 8132 8742
rect 8184 8739 8240 8742
rect 8292 8739 8348 8742
rect 8400 8739 8456 8742
rect 8508 8739 8564 8742
rect 8616 8739 8672 8742
rect 8724 8739 8780 8742
rect 8832 8739 9206 8742
rect 9258 8739 9314 8742
rect 9366 8739 9422 8742
rect 9474 8739 9530 8742
rect 9582 8739 9638 8742
rect 9690 8739 9746 8742
rect 9798 8739 9854 8742
rect 9906 8739 9962 8742
rect 10014 8739 10070 8742
rect 10122 8739 10178 8742
rect 10230 8739 10286 8742
rect 10338 8739 10394 8742
rect 10446 8739 10502 8742
rect 10554 8739 10610 8742
rect 10662 8739 10718 8742
rect 10770 8739 10826 8742
rect 10878 8739 10934 8742
rect 10986 8739 11042 8742
rect 11094 8739 11150 8742
rect 11202 8739 11481 8742
rect 1481 8727 11481 8739
rect 1481 8547 11481 8559
rect 1481 8495 1493 8547
rect 1545 8544 1601 8547
rect 1653 8544 3863 8547
rect 3915 8544 3971 8547
rect 4023 8544 6239 8547
rect 6291 8544 6347 8547
rect 6399 8544 6455 8547
rect 6507 8544 6563 8547
rect 6615 8544 6671 8547
rect 6723 8544 8939 8547
rect 8991 8544 9047 8547
rect 9099 8544 11309 8547
rect 11361 8544 11417 8547
rect 1545 8495 1601 8498
rect 1653 8495 3863 8498
rect 3915 8495 3971 8498
rect 4023 8495 6239 8498
rect 6291 8495 6347 8498
rect 6399 8495 6455 8498
rect 6507 8495 6563 8498
rect 6615 8495 6671 8498
rect 6723 8495 8939 8498
rect 8991 8495 9047 8498
rect 9099 8495 11309 8498
rect 11361 8495 11417 8498
rect 11469 8495 11481 8547
rect 1481 8483 11481 8495
rect 1481 8303 11481 8315
rect 1481 8300 1760 8303
rect 1812 8300 1868 8303
rect 1920 8300 1976 8303
rect 2028 8300 2084 8303
rect 2136 8300 2192 8303
rect 2244 8300 2300 8303
rect 2352 8300 2408 8303
rect 2460 8300 2516 8303
rect 2568 8300 2624 8303
rect 2676 8300 2732 8303
rect 2784 8300 2840 8303
rect 2892 8300 2948 8303
rect 3000 8300 3056 8303
rect 3108 8300 3164 8303
rect 3216 8300 3272 8303
rect 3324 8300 3380 8303
rect 3432 8300 3488 8303
rect 3540 8300 3596 8303
rect 3648 8300 3704 8303
rect 3756 8300 4130 8303
rect 4182 8300 4238 8303
rect 4290 8300 4346 8303
rect 4398 8300 4454 8303
rect 4506 8300 4562 8303
rect 4614 8300 4670 8303
rect 4722 8300 4778 8303
rect 4830 8300 4886 8303
rect 4938 8300 4994 8303
rect 5046 8300 5102 8303
rect 5154 8300 5210 8303
rect 5262 8300 5318 8303
rect 5370 8300 5426 8303
rect 5478 8300 5534 8303
rect 5586 8300 5642 8303
rect 5694 8300 5750 8303
rect 5802 8300 5858 8303
rect 5910 8300 5966 8303
rect 6018 8300 6074 8303
rect 6126 8300 6836 8303
rect 6888 8300 6944 8303
rect 6996 8300 7052 8303
rect 7104 8300 7160 8303
rect 7212 8300 7268 8303
rect 7320 8300 7376 8303
rect 7428 8300 7484 8303
rect 7536 8300 7592 8303
rect 7644 8300 7700 8303
rect 7752 8300 7808 8303
rect 7860 8300 7916 8303
rect 7968 8300 8024 8303
rect 8076 8300 8132 8303
rect 8184 8300 8240 8303
rect 8292 8300 8348 8303
rect 8400 8300 8456 8303
rect 8508 8300 8564 8303
rect 8616 8300 8672 8303
rect 8724 8300 8780 8303
rect 8832 8300 9206 8303
rect 9258 8300 9314 8303
rect 9366 8300 9422 8303
rect 9474 8300 9530 8303
rect 9582 8300 9638 8303
rect 9690 8300 9746 8303
rect 9798 8300 9854 8303
rect 9906 8300 9962 8303
rect 10014 8300 10070 8303
rect 10122 8300 10178 8303
rect 10230 8300 10286 8303
rect 10338 8300 10394 8303
rect 10446 8300 10502 8303
rect 10554 8300 10610 8303
rect 10662 8300 10718 8303
rect 10770 8300 10826 8303
rect 10878 8300 10934 8303
rect 10986 8300 11042 8303
rect 11094 8300 11150 8303
rect 11202 8300 11481 8303
rect 1481 8254 1494 8300
rect 11468 8254 11481 8300
rect 1481 8251 1760 8254
rect 1812 8251 1868 8254
rect 1920 8251 1976 8254
rect 2028 8251 2084 8254
rect 2136 8251 2192 8254
rect 2244 8251 2300 8254
rect 2352 8251 2408 8254
rect 2460 8251 2516 8254
rect 2568 8251 2624 8254
rect 2676 8251 2732 8254
rect 2784 8251 2840 8254
rect 2892 8251 2948 8254
rect 3000 8251 3056 8254
rect 3108 8251 3164 8254
rect 3216 8251 3272 8254
rect 3324 8251 3380 8254
rect 3432 8251 3488 8254
rect 3540 8251 3596 8254
rect 3648 8251 3704 8254
rect 3756 8251 4130 8254
rect 4182 8251 4238 8254
rect 4290 8251 4346 8254
rect 4398 8251 4454 8254
rect 4506 8251 4562 8254
rect 4614 8251 4670 8254
rect 4722 8251 4778 8254
rect 4830 8251 4886 8254
rect 4938 8251 4994 8254
rect 5046 8251 5102 8254
rect 5154 8251 5210 8254
rect 5262 8251 5318 8254
rect 5370 8251 5426 8254
rect 5478 8251 5534 8254
rect 5586 8251 5642 8254
rect 5694 8251 5750 8254
rect 5802 8251 5858 8254
rect 5910 8251 5966 8254
rect 6018 8251 6074 8254
rect 6126 8251 6836 8254
rect 6888 8251 6944 8254
rect 6996 8251 7052 8254
rect 7104 8251 7160 8254
rect 7212 8251 7268 8254
rect 7320 8251 7376 8254
rect 7428 8251 7484 8254
rect 7536 8251 7592 8254
rect 7644 8251 7700 8254
rect 7752 8251 7808 8254
rect 7860 8251 7916 8254
rect 7968 8251 8024 8254
rect 8076 8251 8132 8254
rect 8184 8251 8240 8254
rect 8292 8251 8348 8254
rect 8400 8251 8456 8254
rect 8508 8251 8564 8254
rect 8616 8251 8672 8254
rect 8724 8251 8780 8254
rect 8832 8251 9206 8254
rect 9258 8251 9314 8254
rect 9366 8251 9422 8254
rect 9474 8251 9530 8254
rect 9582 8251 9638 8254
rect 9690 8251 9746 8254
rect 9798 8251 9854 8254
rect 9906 8251 9962 8254
rect 10014 8251 10070 8254
rect 10122 8251 10178 8254
rect 10230 8251 10286 8254
rect 10338 8251 10394 8254
rect 10446 8251 10502 8254
rect 10554 8251 10610 8254
rect 10662 8251 10718 8254
rect 10770 8251 10826 8254
rect 10878 8251 10934 8254
rect 10986 8251 11042 8254
rect 11094 8251 11150 8254
rect 11202 8251 11481 8254
rect 1481 8239 11481 8251
rect 1481 8059 11481 8071
rect 1481 8007 1493 8059
rect 1545 8056 1601 8059
rect 1653 8056 3863 8059
rect 3915 8056 3971 8059
rect 4023 8056 6239 8059
rect 6291 8056 6347 8059
rect 6399 8056 6455 8059
rect 6507 8056 6563 8059
rect 6615 8056 6671 8059
rect 6723 8056 8939 8059
rect 8991 8056 9047 8059
rect 9099 8056 11309 8059
rect 11361 8056 11417 8059
rect 1545 8007 1601 8010
rect 1653 8007 3863 8010
rect 3915 8007 3971 8010
rect 4023 8007 6239 8010
rect 6291 8007 6347 8010
rect 6399 8007 6455 8010
rect 6507 8007 6563 8010
rect 6615 8007 6671 8010
rect 6723 8007 8939 8010
rect 8991 8007 9047 8010
rect 9099 8007 11309 8010
rect 11361 8007 11417 8010
rect 11469 8007 11481 8059
rect 1481 7995 11481 8007
rect 1481 7815 11481 7827
rect 1481 7812 1760 7815
rect 1812 7812 1868 7815
rect 1920 7812 1976 7815
rect 2028 7812 2084 7815
rect 2136 7812 2192 7815
rect 2244 7812 2300 7815
rect 2352 7812 2408 7815
rect 2460 7812 2516 7815
rect 2568 7812 2624 7815
rect 2676 7812 2732 7815
rect 2784 7812 2840 7815
rect 2892 7812 2948 7815
rect 3000 7812 3056 7815
rect 3108 7812 3164 7815
rect 3216 7812 3272 7815
rect 3324 7812 3380 7815
rect 3432 7812 3488 7815
rect 3540 7812 3596 7815
rect 3648 7812 3704 7815
rect 3756 7812 4130 7815
rect 4182 7812 4238 7815
rect 4290 7812 4346 7815
rect 4398 7812 4454 7815
rect 4506 7812 4562 7815
rect 4614 7812 4670 7815
rect 4722 7812 4778 7815
rect 4830 7812 4886 7815
rect 4938 7812 4994 7815
rect 5046 7812 5102 7815
rect 5154 7812 5210 7815
rect 5262 7812 5318 7815
rect 5370 7812 5426 7815
rect 5478 7812 5534 7815
rect 5586 7812 5642 7815
rect 5694 7812 5750 7815
rect 5802 7812 5858 7815
rect 5910 7812 5966 7815
rect 6018 7812 6074 7815
rect 6126 7812 6836 7815
rect 6888 7812 6944 7815
rect 6996 7812 7052 7815
rect 7104 7812 7160 7815
rect 7212 7812 7268 7815
rect 7320 7812 7376 7815
rect 7428 7812 7484 7815
rect 7536 7812 7592 7815
rect 7644 7812 7700 7815
rect 7752 7812 7808 7815
rect 7860 7812 7916 7815
rect 7968 7812 8024 7815
rect 8076 7812 8132 7815
rect 8184 7812 8240 7815
rect 8292 7812 8348 7815
rect 8400 7812 8456 7815
rect 8508 7812 8564 7815
rect 8616 7812 8672 7815
rect 8724 7812 8780 7815
rect 8832 7812 9206 7815
rect 9258 7812 9314 7815
rect 9366 7812 9422 7815
rect 9474 7812 9530 7815
rect 9582 7812 9638 7815
rect 9690 7812 9746 7815
rect 9798 7812 9854 7815
rect 9906 7812 9962 7815
rect 10014 7812 10070 7815
rect 10122 7812 10178 7815
rect 10230 7812 10286 7815
rect 10338 7812 10394 7815
rect 10446 7812 10502 7815
rect 10554 7812 10610 7815
rect 10662 7812 10718 7815
rect 10770 7812 10826 7815
rect 10878 7812 10934 7815
rect 10986 7812 11042 7815
rect 11094 7812 11150 7815
rect 11202 7812 11481 7815
rect 1481 7766 1494 7812
rect 11468 7766 11481 7812
rect 1481 7763 1760 7766
rect 1812 7763 1868 7766
rect 1920 7763 1976 7766
rect 2028 7763 2084 7766
rect 2136 7763 2192 7766
rect 2244 7763 2300 7766
rect 2352 7763 2408 7766
rect 2460 7763 2516 7766
rect 2568 7763 2624 7766
rect 2676 7763 2732 7766
rect 2784 7763 2840 7766
rect 2892 7763 2948 7766
rect 3000 7763 3056 7766
rect 3108 7763 3164 7766
rect 3216 7763 3272 7766
rect 3324 7763 3380 7766
rect 3432 7763 3488 7766
rect 3540 7763 3596 7766
rect 3648 7763 3704 7766
rect 3756 7763 4130 7766
rect 4182 7763 4238 7766
rect 4290 7763 4346 7766
rect 4398 7763 4454 7766
rect 4506 7763 4562 7766
rect 4614 7763 4670 7766
rect 4722 7763 4778 7766
rect 4830 7763 4886 7766
rect 4938 7763 4994 7766
rect 5046 7763 5102 7766
rect 5154 7763 5210 7766
rect 5262 7763 5318 7766
rect 5370 7763 5426 7766
rect 5478 7763 5534 7766
rect 5586 7763 5642 7766
rect 5694 7763 5750 7766
rect 5802 7763 5858 7766
rect 5910 7763 5966 7766
rect 6018 7763 6074 7766
rect 6126 7763 6836 7766
rect 6888 7763 6944 7766
rect 6996 7763 7052 7766
rect 7104 7763 7160 7766
rect 7212 7763 7268 7766
rect 7320 7763 7376 7766
rect 7428 7763 7484 7766
rect 7536 7763 7592 7766
rect 7644 7763 7700 7766
rect 7752 7763 7808 7766
rect 7860 7763 7916 7766
rect 7968 7763 8024 7766
rect 8076 7763 8132 7766
rect 8184 7763 8240 7766
rect 8292 7763 8348 7766
rect 8400 7763 8456 7766
rect 8508 7763 8564 7766
rect 8616 7763 8672 7766
rect 8724 7763 8780 7766
rect 8832 7763 9206 7766
rect 9258 7763 9314 7766
rect 9366 7763 9422 7766
rect 9474 7763 9530 7766
rect 9582 7763 9638 7766
rect 9690 7763 9746 7766
rect 9798 7763 9854 7766
rect 9906 7763 9962 7766
rect 10014 7763 10070 7766
rect 10122 7763 10178 7766
rect 10230 7763 10286 7766
rect 10338 7763 10394 7766
rect 10446 7763 10502 7766
rect 10554 7763 10610 7766
rect 10662 7763 10718 7766
rect 10770 7763 10826 7766
rect 10878 7763 10934 7766
rect 10986 7763 11042 7766
rect 11094 7763 11150 7766
rect 11202 7763 11481 7766
rect 1481 7751 11481 7763
rect 1481 7571 11481 7583
rect 1481 7519 1493 7571
rect 1545 7568 1601 7571
rect 1653 7568 3863 7571
rect 3915 7568 3971 7571
rect 4023 7568 6239 7571
rect 6291 7568 6347 7571
rect 6399 7568 6455 7571
rect 6507 7568 6563 7571
rect 6615 7568 6671 7571
rect 6723 7568 8939 7571
rect 8991 7568 9047 7571
rect 9099 7568 11309 7571
rect 11361 7568 11417 7571
rect 1545 7519 1601 7522
rect 1653 7519 3863 7522
rect 3915 7519 3971 7522
rect 4023 7519 6239 7522
rect 6291 7519 6347 7522
rect 6399 7519 6455 7522
rect 6507 7519 6563 7522
rect 6615 7519 6671 7522
rect 6723 7519 8939 7522
rect 8991 7519 9047 7522
rect 9099 7519 11309 7522
rect 11361 7519 11417 7522
rect 11469 7519 11481 7571
rect 1481 7507 11481 7519
rect 1213 7391 1413 7418
rect 1213 7339 1233 7391
rect 1285 7339 1341 7391
rect 1393 7339 1413 7391
rect 11549 7418 11560 12064
rect 11706 12035 11749 12064
rect 11729 11983 11749 12035
rect 11706 11927 11749 11983
rect 11729 11875 11749 11927
rect 11706 11819 11749 11875
rect 11729 11767 11749 11819
rect 11706 11711 11749 11767
rect 11729 11659 11749 11711
rect 11706 11603 11749 11659
rect 11729 11551 11749 11603
rect 11706 11495 11749 11551
rect 11729 11443 11749 11495
rect 11706 11387 11749 11443
rect 11729 11335 11749 11387
rect 11706 11279 11749 11335
rect 11729 11227 11749 11279
rect 11706 11171 11749 11227
rect 11729 11119 11749 11171
rect 11706 11063 11749 11119
rect 11729 11011 11749 11063
rect 11706 10955 11749 11011
rect 11729 10903 11749 10955
rect 11706 10847 11749 10903
rect 11729 10795 11749 10847
rect 11706 10739 11749 10795
rect 11729 10687 11749 10739
rect 11706 10631 11749 10687
rect 11729 10579 11749 10631
rect 11706 10523 11749 10579
rect 11729 10471 11749 10523
rect 11706 10415 11749 10471
rect 11729 10363 11749 10415
rect 11706 10307 11749 10363
rect 11729 10255 11749 10307
rect 11706 10199 11749 10255
rect 11729 10147 11749 10199
rect 11706 10091 11749 10147
rect 11729 10039 11749 10091
rect 11706 9983 11749 10039
rect 11729 9931 11749 9983
rect 11706 9875 11749 9931
rect 11729 9823 11749 9875
rect 11706 9767 11749 9823
rect 11729 9715 11749 9767
rect 11706 9659 11749 9715
rect 11729 9607 11749 9659
rect 11706 9551 11749 9607
rect 11729 9499 11749 9551
rect 11706 9443 11749 9499
rect 11729 9391 11749 9443
rect 11706 9335 11749 9391
rect 11729 9283 11749 9335
rect 11706 9227 11749 9283
rect 11729 9175 11749 9227
rect 11706 9119 11749 9175
rect 11729 9067 11749 9119
rect 11706 9011 11749 9067
rect 11729 8959 11749 9011
rect 11706 8903 11749 8959
rect 11729 8851 11749 8903
rect 11706 8795 11749 8851
rect 11729 8743 11749 8795
rect 11706 8687 11749 8743
rect 11729 8635 11749 8687
rect 11706 8579 11749 8635
rect 11729 8527 11749 8579
rect 11706 8471 11749 8527
rect 11729 8419 11749 8471
rect 11706 8363 11749 8419
rect 11729 8311 11749 8363
rect 11706 8255 11749 8311
rect 11729 8203 11749 8255
rect 11706 8147 11749 8203
rect 11729 8095 11749 8147
rect 11706 8039 11749 8095
rect 11729 7987 11749 8039
rect 11706 7931 11749 7987
rect 11729 7879 11749 7931
rect 11706 7823 11749 7879
rect 11729 7771 11749 7823
rect 11706 7715 11749 7771
rect 11729 7663 11749 7715
rect 11706 7607 11749 7663
rect 11729 7555 11749 7607
rect 11706 7499 11749 7555
rect 11729 7447 11749 7499
rect 11706 7418 11749 7447
rect 11549 7391 11749 7418
rect 11549 7339 11569 7391
rect 11621 7339 11677 7391
rect 11729 7339 11749 7391
rect 1213 7176 1413 7339
rect 1481 7327 11481 7339
rect 1481 7324 1760 7327
rect 1812 7324 1868 7327
rect 1920 7324 1976 7327
rect 2028 7324 2084 7327
rect 2136 7324 2192 7327
rect 2244 7324 2300 7327
rect 2352 7324 2408 7327
rect 2460 7324 2516 7327
rect 2568 7324 2624 7327
rect 2676 7324 2732 7327
rect 2784 7324 2840 7327
rect 2892 7324 2948 7327
rect 3000 7324 3056 7327
rect 3108 7324 3164 7327
rect 3216 7324 3272 7327
rect 3324 7324 3380 7327
rect 3432 7324 3488 7327
rect 3540 7324 3596 7327
rect 3648 7324 3704 7327
rect 3756 7324 4130 7327
rect 4182 7324 4238 7327
rect 4290 7324 4346 7327
rect 4398 7324 4454 7327
rect 4506 7324 4562 7327
rect 4614 7324 4670 7327
rect 4722 7324 4778 7327
rect 4830 7324 4886 7327
rect 4938 7324 4994 7327
rect 5046 7324 5102 7327
rect 5154 7324 5210 7327
rect 5262 7324 5318 7327
rect 5370 7324 5426 7327
rect 5478 7324 5534 7327
rect 5586 7324 5642 7327
rect 5694 7324 5750 7327
rect 5802 7324 5858 7327
rect 5910 7324 5966 7327
rect 6018 7324 6074 7327
rect 6126 7324 6836 7327
rect 6888 7324 6944 7327
rect 6996 7324 7052 7327
rect 7104 7324 7160 7327
rect 7212 7324 7268 7327
rect 7320 7324 7376 7327
rect 7428 7324 7484 7327
rect 7536 7324 7592 7327
rect 7644 7324 7700 7327
rect 7752 7324 7808 7327
rect 7860 7324 7916 7327
rect 7968 7324 8024 7327
rect 8076 7324 8132 7327
rect 8184 7324 8240 7327
rect 8292 7324 8348 7327
rect 8400 7324 8456 7327
rect 8508 7324 8564 7327
rect 8616 7324 8672 7327
rect 8724 7324 8780 7327
rect 8832 7324 9206 7327
rect 9258 7324 9314 7327
rect 9366 7324 9422 7327
rect 9474 7324 9530 7327
rect 9582 7324 9638 7327
rect 9690 7324 9746 7327
rect 9798 7324 9854 7327
rect 9906 7324 9962 7327
rect 10014 7324 10070 7327
rect 10122 7324 10178 7327
rect 10230 7324 10286 7327
rect 10338 7324 10394 7327
rect 10446 7324 10502 7327
rect 10554 7324 10610 7327
rect 10662 7324 10718 7327
rect 10770 7324 10826 7327
rect 10878 7324 10934 7327
rect 10986 7324 11042 7327
rect 11094 7324 11150 7327
rect 11202 7324 11481 7327
rect 1481 7278 1494 7324
rect 11468 7278 11481 7324
rect 1481 7275 1760 7278
rect 1812 7275 1868 7278
rect 1920 7275 1976 7278
rect 2028 7275 2084 7278
rect 2136 7275 2192 7278
rect 2244 7275 2300 7278
rect 2352 7275 2408 7278
rect 2460 7275 2516 7278
rect 2568 7275 2624 7278
rect 2676 7275 2732 7278
rect 2784 7275 2840 7278
rect 2892 7275 2948 7278
rect 3000 7275 3056 7278
rect 3108 7275 3164 7278
rect 3216 7275 3272 7278
rect 3324 7275 3380 7278
rect 3432 7275 3488 7278
rect 3540 7275 3596 7278
rect 3648 7275 3704 7278
rect 3756 7275 4130 7278
rect 4182 7275 4238 7278
rect 4290 7275 4346 7278
rect 4398 7275 4454 7278
rect 4506 7275 4562 7278
rect 4614 7275 4670 7278
rect 4722 7275 4778 7278
rect 4830 7275 4886 7278
rect 4938 7275 4994 7278
rect 5046 7275 5102 7278
rect 5154 7275 5210 7278
rect 5262 7275 5318 7278
rect 5370 7275 5426 7278
rect 5478 7275 5534 7278
rect 5586 7275 5642 7278
rect 5694 7275 5750 7278
rect 5802 7275 5858 7278
rect 5910 7275 5966 7278
rect 6018 7275 6074 7278
rect 6126 7275 6836 7278
rect 6888 7275 6944 7278
rect 6996 7275 7052 7278
rect 7104 7275 7160 7278
rect 7212 7275 7268 7278
rect 7320 7275 7376 7278
rect 7428 7275 7484 7278
rect 7536 7275 7592 7278
rect 7644 7275 7700 7278
rect 7752 7275 7808 7278
rect 7860 7275 7916 7278
rect 7968 7275 8024 7278
rect 8076 7275 8132 7278
rect 8184 7275 8240 7278
rect 8292 7275 8348 7278
rect 8400 7275 8456 7278
rect 8508 7275 8564 7278
rect 8616 7275 8672 7278
rect 8724 7275 8780 7278
rect 8832 7275 9206 7278
rect 9258 7275 9314 7278
rect 9366 7275 9422 7278
rect 9474 7275 9530 7278
rect 9582 7275 9638 7278
rect 9690 7275 9746 7278
rect 9798 7275 9854 7278
rect 9906 7275 9962 7278
rect 10014 7275 10070 7278
rect 10122 7275 10178 7278
rect 10230 7275 10286 7278
rect 10338 7275 10394 7278
rect 10446 7275 10502 7278
rect 10554 7275 10610 7278
rect 10662 7275 10718 7278
rect 10770 7275 10826 7278
rect 10878 7275 10934 7278
rect 10986 7275 11042 7278
rect 11094 7275 11150 7278
rect 11202 7275 11481 7278
rect 1481 7263 11481 7275
rect 11549 7176 11749 7339
rect 1213 6976 11749 7176
rect 12001 6897 12012 12585
rect 950 6885 12012 6897
rect 950 6878 1760 6885
rect 1812 6878 1868 6885
rect 1920 6878 1976 6885
rect 2028 6878 2084 6885
rect 2136 6878 2192 6885
rect 2244 6878 2300 6885
rect 2352 6878 2408 6885
rect 2460 6878 2516 6885
rect 2568 6878 2624 6885
rect 2676 6878 2732 6885
rect 2784 6878 2840 6885
rect 2892 6878 2948 6885
rect 3000 6878 3056 6885
rect 3108 6878 3164 6885
rect 3216 6878 3272 6885
rect 3324 6878 3380 6885
rect 3432 6878 3488 6885
rect 3540 6878 3596 6885
rect 3648 6878 3704 6885
rect 3756 6878 4130 6885
rect 4182 6878 4238 6885
rect 4290 6878 4346 6885
rect 4398 6878 4454 6885
rect 4506 6878 4562 6885
rect 4614 6878 4670 6885
rect 4722 6878 4778 6885
rect 4830 6878 4886 6885
rect 4938 6878 4994 6885
rect 5046 6878 5102 6885
rect 5154 6878 5210 6885
rect 5262 6878 5318 6885
rect 5370 6878 5426 6885
rect 5478 6878 5534 6885
rect 5586 6878 5642 6885
rect 5694 6878 5750 6885
rect 5802 6878 5858 6885
rect 5910 6878 5966 6885
rect 6018 6878 6074 6885
rect 6126 6878 6836 6885
rect 6888 6878 6944 6885
rect 6996 6878 7052 6885
rect 7104 6878 7160 6885
rect 7212 6878 7268 6885
rect 7320 6878 7376 6885
rect 7428 6878 7484 6885
rect 7536 6878 7592 6885
rect 7644 6878 7700 6885
rect 7752 6878 7808 6885
rect 7860 6878 7916 6885
rect 7968 6878 8024 6885
rect 8076 6878 8132 6885
rect 8184 6878 8240 6885
rect 8292 6878 8348 6885
rect 8400 6878 8456 6885
rect 8508 6878 8564 6885
rect 8616 6878 8672 6885
rect 8724 6878 8780 6885
rect 8832 6878 9206 6885
rect 9258 6878 9314 6885
rect 9366 6878 9422 6885
rect 9474 6878 9530 6885
rect 9582 6878 9638 6885
rect 9690 6878 9746 6885
rect 9798 6878 9854 6885
rect 9906 6878 9962 6885
rect 10014 6878 10070 6885
rect 10122 6878 10178 6885
rect 10230 6878 10286 6885
rect 10338 6878 10394 6885
rect 10446 6878 10502 6885
rect 10554 6878 10610 6885
rect 10662 6878 10718 6885
rect 10770 6878 10826 6885
rect 10878 6878 10934 6885
rect 10986 6878 11042 6885
rect 11094 6878 11150 6885
rect 11202 6878 12012 6885
rect 950 6732 1058 6878
rect 11904 6732 12012 6878
rect 950 6725 1760 6732
rect 1812 6725 1868 6732
rect 1920 6725 1976 6732
rect 2028 6725 2084 6732
rect 2136 6725 2192 6732
rect 2244 6725 2300 6732
rect 2352 6725 2408 6732
rect 2460 6725 2516 6732
rect 2568 6725 2624 6732
rect 2676 6725 2732 6732
rect 2784 6725 2840 6732
rect 2892 6725 2948 6732
rect 3000 6725 3056 6732
rect 3108 6725 3164 6732
rect 3216 6725 3272 6732
rect 3324 6725 3380 6732
rect 3432 6725 3488 6732
rect 3540 6725 3596 6732
rect 3648 6725 3704 6732
rect 3756 6725 4130 6732
rect 4182 6725 4238 6732
rect 4290 6725 4346 6732
rect 4398 6725 4454 6732
rect 4506 6725 4562 6732
rect 4614 6725 4670 6732
rect 4722 6725 4778 6732
rect 4830 6725 4886 6732
rect 4938 6725 4994 6732
rect 5046 6725 5102 6732
rect 5154 6725 5210 6732
rect 5262 6725 5318 6732
rect 5370 6725 5426 6732
rect 5478 6725 5534 6732
rect 5586 6725 5642 6732
rect 5694 6725 5750 6732
rect 5802 6725 5858 6732
rect 5910 6725 5966 6732
rect 6018 6725 6074 6732
rect 6126 6725 6836 6732
rect 6888 6725 6944 6732
rect 6996 6725 7052 6732
rect 7104 6725 7160 6732
rect 7212 6725 7268 6732
rect 7320 6725 7376 6732
rect 7428 6725 7484 6732
rect 7536 6725 7592 6732
rect 7644 6725 7700 6732
rect 7752 6725 7808 6732
rect 7860 6725 7916 6732
rect 7968 6725 8024 6732
rect 8076 6725 8132 6732
rect 8184 6725 8240 6732
rect 8292 6725 8348 6732
rect 8400 6725 8456 6732
rect 8508 6725 8564 6732
rect 8616 6725 8672 6732
rect 8724 6725 8780 6732
rect 8832 6725 9206 6732
rect 9258 6725 9314 6732
rect 9366 6725 9422 6732
rect 9474 6725 9530 6732
rect 9582 6725 9638 6732
rect 9690 6725 9746 6732
rect 9798 6725 9854 6732
rect 9906 6725 9962 6732
rect 10014 6725 10070 6732
rect 10122 6725 10178 6732
rect 10230 6725 10286 6732
rect 10338 6725 10394 6732
rect 10446 6725 10502 6732
rect 10554 6725 10610 6732
rect 10662 6725 10718 6732
rect 10770 6725 10826 6732
rect 10878 6725 10934 6732
rect 10986 6725 11042 6732
rect 11094 6725 11150 6732
rect 11202 6725 12012 6732
rect 950 6713 12012 6725
rect 950 1011 961 6713
rect 1213 6434 11749 6634
rect 1213 6271 1413 6434
rect 1481 6335 11481 6347
rect 1481 6332 1760 6335
rect 1812 6332 1868 6335
rect 1920 6332 1976 6335
rect 2028 6332 2084 6335
rect 2136 6332 2192 6335
rect 2244 6332 2300 6335
rect 2352 6332 2408 6335
rect 2460 6332 2516 6335
rect 2568 6332 2624 6335
rect 2676 6332 2732 6335
rect 2784 6332 2840 6335
rect 2892 6332 2948 6335
rect 3000 6332 3056 6335
rect 3108 6332 3164 6335
rect 3216 6332 3272 6335
rect 3324 6332 3380 6335
rect 3432 6332 3488 6335
rect 3540 6332 3596 6335
rect 3648 6332 3704 6335
rect 3756 6332 4130 6335
rect 4182 6332 4238 6335
rect 4290 6332 4346 6335
rect 4398 6332 4454 6335
rect 4506 6332 4562 6335
rect 4614 6332 4670 6335
rect 4722 6332 4778 6335
rect 4830 6332 4886 6335
rect 4938 6332 4994 6335
rect 5046 6332 5102 6335
rect 5154 6332 5210 6335
rect 5262 6332 5318 6335
rect 5370 6332 5426 6335
rect 5478 6332 5534 6335
rect 5586 6332 5642 6335
rect 5694 6332 5750 6335
rect 5802 6332 5858 6335
rect 5910 6332 5966 6335
rect 6018 6332 6074 6335
rect 6126 6332 6836 6335
rect 6888 6332 6944 6335
rect 6996 6332 7052 6335
rect 7104 6332 7160 6335
rect 7212 6332 7268 6335
rect 7320 6332 7376 6335
rect 7428 6332 7484 6335
rect 7536 6332 7592 6335
rect 7644 6332 7700 6335
rect 7752 6332 7808 6335
rect 7860 6332 7916 6335
rect 7968 6332 8024 6335
rect 8076 6332 8132 6335
rect 8184 6332 8240 6335
rect 8292 6332 8348 6335
rect 8400 6332 8456 6335
rect 8508 6332 8564 6335
rect 8616 6332 8672 6335
rect 8724 6332 8780 6335
rect 8832 6332 9206 6335
rect 9258 6332 9314 6335
rect 9366 6332 9422 6335
rect 9474 6332 9530 6335
rect 9582 6332 9638 6335
rect 9690 6332 9746 6335
rect 9798 6332 9854 6335
rect 9906 6332 9962 6335
rect 10014 6332 10070 6335
rect 10122 6332 10178 6335
rect 10230 6332 10286 6335
rect 10338 6332 10394 6335
rect 10446 6332 10502 6335
rect 10554 6332 10610 6335
rect 10662 6332 10718 6335
rect 10770 6332 10826 6335
rect 10878 6332 10934 6335
rect 10986 6332 11042 6335
rect 11094 6332 11150 6335
rect 11202 6332 11481 6335
rect 1481 6286 1494 6332
rect 11468 6286 11481 6332
rect 1481 6283 1760 6286
rect 1812 6283 1868 6286
rect 1920 6283 1976 6286
rect 2028 6283 2084 6286
rect 2136 6283 2192 6286
rect 2244 6283 2300 6286
rect 2352 6283 2408 6286
rect 2460 6283 2516 6286
rect 2568 6283 2624 6286
rect 2676 6283 2732 6286
rect 2784 6283 2840 6286
rect 2892 6283 2948 6286
rect 3000 6283 3056 6286
rect 3108 6283 3164 6286
rect 3216 6283 3272 6286
rect 3324 6283 3380 6286
rect 3432 6283 3488 6286
rect 3540 6283 3596 6286
rect 3648 6283 3704 6286
rect 3756 6283 4130 6286
rect 4182 6283 4238 6286
rect 4290 6283 4346 6286
rect 4398 6283 4454 6286
rect 4506 6283 4562 6286
rect 4614 6283 4670 6286
rect 4722 6283 4778 6286
rect 4830 6283 4886 6286
rect 4938 6283 4994 6286
rect 5046 6283 5102 6286
rect 5154 6283 5210 6286
rect 5262 6283 5318 6286
rect 5370 6283 5426 6286
rect 5478 6283 5534 6286
rect 5586 6283 5642 6286
rect 5694 6283 5750 6286
rect 5802 6283 5858 6286
rect 5910 6283 5966 6286
rect 6018 6283 6074 6286
rect 6126 6283 6836 6286
rect 6888 6283 6944 6286
rect 6996 6283 7052 6286
rect 7104 6283 7160 6286
rect 7212 6283 7268 6286
rect 7320 6283 7376 6286
rect 7428 6283 7484 6286
rect 7536 6283 7592 6286
rect 7644 6283 7700 6286
rect 7752 6283 7808 6286
rect 7860 6283 7916 6286
rect 7968 6283 8024 6286
rect 8076 6283 8132 6286
rect 8184 6283 8240 6286
rect 8292 6283 8348 6286
rect 8400 6283 8456 6286
rect 8508 6283 8564 6286
rect 8616 6283 8672 6286
rect 8724 6283 8780 6286
rect 8832 6283 9206 6286
rect 9258 6283 9314 6286
rect 9366 6283 9422 6286
rect 9474 6283 9530 6286
rect 9582 6283 9638 6286
rect 9690 6283 9746 6286
rect 9798 6283 9854 6286
rect 9906 6283 9962 6286
rect 10014 6283 10070 6286
rect 10122 6283 10178 6286
rect 10230 6283 10286 6286
rect 10338 6283 10394 6286
rect 10446 6283 10502 6286
rect 10554 6283 10610 6286
rect 10662 6283 10718 6286
rect 10770 6283 10826 6286
rect 10878 6283 10934 6286
rect 10986 6283 11042 6286
rect 11094 6283 11150 6286
rect 11202 6283 11481 6286
rect 1481 6271 11481 6283
rect 11549 6271 11749 6434
rect 1213 6219 1233 6271
rect 1285 6219 1341 6271
rect 1393 6219 1413 6271
rect 1213 6192 1413 6219
rect 1213 6163 1256 6192
rect 1213 6111 1233 6163
rect 1213 6055 1256 6111
rect 1213 6003 1233 6055
rect 1213 5947 1256 6003
rect 1213 5895 1233 5947
rect 1213 5839 1256 5895
rect 1213 5787 1233 5839
rect 1213 5731 1256 5787
rect 1213 5679 1233 5731
rect 1213 5623 1256 5679
rect 1213 5571 1233 5623
rect 1213 5515 1256 5571
rect 1213 5463 1233 5515
rect 1213 5407 1256 5463
rect 1213 5355 1233 5407
rect 1213 5299 1256 5355
rect 1213 5247 1233 5299
rect 1213 5191 1256 5247
rect 1213 5139 1233 5191
rect 1213 5083 1256 5139
rect 1213 5031 1233 5083
rect 1213 4975 1256 5031
rect 1213 4923 1233 4975
rect 1213 4867 1256 4923
rect 1213 4815 1233 4867
rect 1213 4759 1256 4815
rect 1213 4707 1233 4759
rect 1213 4651 1256 4707
rect 1213 4599 1233 4651
rect 1213 4543 1256 4599
rect 1213 4491 1233 4543
rect 1213 4435 1256 4491
rect 1213 4383 1233 4435
rect 1213 4327 1256 4383
rect 1213 4275 1233 4327
rect 1213 4219 1256 4275
rect 1213 4167 1233 4219
rect 1213 4111 1256 4167
rect 1213 4059 1233 4111
rect 1213 4003 1256 4059
rect 1213 3951 1233 4003
rect 1213 3895 1256 3951
rect 1213 3843 1233 3895
rect 1213 3787 1256 3843
rect 1213 3735 1233 3787
rect 1213 3679 1256 3735
rect 1213 3627 1233 3679
rect 1213 3571 1256 3627
rect 1213 3519 1233 3571
rect 1213 3463 1256 3519
rect 1213 3411 1233 3463
rect 1213 3355 1256 3411
rect 1213 3303 1233 3355
rect 1213 3247 1256 3303
rect 1213 3195 1233 3247
rect 1213 3139 1256 3195
rect 1213 3087 1233 3139
rect 1213 3031 1256 3087
rect 1213 2979 1233 3031
rect 1213 2923 1256 2979
rect 1213 2871 1233 2923
rect 1213 2815 1256 2871
rect 1213 2763 1233 2815
rect 1213 2707 1256 2763
rect 1213 2655 1233 2707
rect 1213 2599 1256 2655
rect 1213 2547 1233 2599
rect 1213 2491 1256 2547
rect 1213 2439 1233 2491
rect 1213 2383 1256 2439
rect 1213 2331 1233 2383
rect 1213 2275 1256 2331
rect 1213 2223 1233 2275
rect 1213 2167 1256 2223
rect 1213 2115 1233 2167
rect 1213 2059 1256 2115
rect 1213 2007 1233 2059
rect 1213 1951 1256 2007
rect 1213 1899 1233 1951
rect 1213 1843 1256 1899
rect 1213 1791 1233 1843
rect 1213 1735 1256 1791
rect 1213 1683 1233 1735
rect 1213 1627 1256 1683
rect 1213 1575 1233 1627
rect 1213 1546 1256 1575
rect 1402 1546 1413 6192
rect 11549 6219 11569 6271
rect 11621 6219 11677 6271
rect 11729 6219 11749 6271
rect 11549 6192 11749 6219
rect 1481 6091 11481 6103
rect 1481 6039 1493 6091
rect 1545 6088 1601 6091
rect 1653 6088 3863 6091
rect 3915 6088 3971 6091
rect 4023 6088 6239 6091
rect 6291 6088 6347 6091
rect 6399 6088 6455 6091
rect 6507 6088 6563 6091
rect 6615 6088 6671 6091
rect 6723 6088 8939 6091
rect 8991 6088 9047 6091
rect 9099 6088 11309 6091
rect 11361 6088 11417 6091
rect 1545 6039 1601 6042
rect 1653 6039 3863 6042
rect 3915 6039 3971 6042
rect 4023 6039 6239 6042
rect 6291 6039 6347 6042
rect 6399 6039 6455 6042
rect 6507 6039 6563 6042
rect 6615 6039 6671 6042
rect 6723 6039 8939 6042
rect 8991 6039 9047 6042
rect 9099 6039 11309 6042
rect 11361 6039 11417 6042
rect 11469 6039 11481 6091
rect 1481 6027 11481 6039
rect 1481 5847 11481 5859
rect 1481 5844 1760 5847
rect 1812 5844 1868 5847
rect 1920 5844 1976 5847
rect 2028 5844 2084 5847
rect 2136 5844 2192 5847
rect 2244 5844 2300 5847
rect 2352 5844 2408 5847
rect 2460 5844 2516 5847
rect 2568 5844 2624 5847
rect 2676 5844 2732 5847
rect 2784 5844 2840 5847
rect 2892 5844 2948 5847
rect 3000 5844 3056 5847
rect 3108 5844 3164 5847
rect 3216 5844 3272 5847
rect 3324 5844 3380 5847
rect 3432 5844 3488 5847
rect 3540 5844 3596 5847
rect 3648 5844 3704 5847
rect 3756 5844 4130 5847
rect 4182 5844 4238 5847
rect 4290 5844 4346 5847
rect 4398 5844 4454 5847
rect 4506 5844 4562 5847
rect 4614 5844 4670 5847
rect 4722 5844 4778 5847
rect 4830 5844 4886 5847
rect 4938 5844 4994 5847
rect 5046 5844 5102 5847
rect 5154 5844 5210 5847
rect 5262 5844 5318 5847
rect 5370 5844 5426 5847
rect 5478 5844 5534 5847
rect 5586 5844 5642 5847
rect 5694 5844 5750 5847
rect 5802 5844 5858 5847
rect 5910 5844 5966 5847
rect 6018 5844 6074 5847
rect 6126 5844 6836 5847
rect 6888 5844 6944 5847
rect 6996 5844 7052 5847
rect 7104 5844 7160 5847
rect 7212 5844 7268 5847
rect 7320 5844 7376 5847
rect 7428 5844 7484 5847
rect 7536 5844 7592 5847
rect 7644 5844 7700 5847
rect 7752 5844 7808 5847
rect 7860 5844 7916 5847
rect 7968 5844 8024 5847
rect 8076 5844 8132 5847
rect 8184 5844 8240 5847
rect 8292 5844 8348 5847
rect 8400 5844 8456 5847
rect 8508 5844 8564 5847
rect 8616 5844 8672 5847
rect 8724 5844 8780 5847
rect 8832 5844 9206 5847
rect 9258 5844 9314 5847
rect 9366 5844 9422 5847
rect 9474 5844 9530 5847
rect 9582 5844 9638 5847
rect 9690 5844 9746 5847
rect 9798 5844 9854 5847
rect 9906 5844 9962 5847
rect 10014 5844 10070 5847
rect 10122 5844 10178 5847
rect 10230 5844 10286 5847
rect 10338 5844 10394 5847
rect 10446 5844 10502 5847
rect 10554 5844 10610 5847
rect 10662 5844 10718 5847
rect 10770 5844 10826 5847
rect 10878 5844 10934 5847
rect 10986 5844 11042 5847
rect 11094 5844 11150 5847
rect 11202 5844 11481 5847
rect 1481 5798 1494 5844
rect 11468 5798 11481 5844
rect 1481 5795 1760 5798
rect 1812 5795 1868 5798
rect 1920 5795 1976 5798
rect 2028 5795 2084 5798
rect 2136 5795 2192 5798
rect 2244 5795 2300 5798
rect 2352 5795 2408 5798
rect 2460 5795 2516 5798
rect 2568 5795 2624 5798
rect 2676 5795 2732 5798
rect 2784 5795 2840 5798
rect 2892 5795 2948 5798
rect 3000 5795 3056 5798
rect 3108 5795 3164 5798
rect 3216 5795 3272 5798
rect 3324 5795 3380 5798
rect 3432 5795 3488 5798
rect 3540 5795 3596 5798
rect 3648 5795 3704 5798
rect 3756 5795 4130 5798
rect 4182 5795 4238 5798
rect 4290 5795 4346 5798
rect 4398 5795 4454 5798
rect 4506 5795 4562 5798
rect 4614 5795 4670 5798
rect 4722 5795 4778 5798
rect 4830 5795 4886 5798
rect 4938 5795 4994 5798
rect 5046 5795 5102 5798
rect 5154 5795 5210 5798
rect 5262 5795 5318 5798
rect 5370 5795 5426 5798
rect 5478 5795 5534 5798
rect 5586 5795 5642 5798
rect 5694 5795 5750 5798
rect 5802 5795 5858 5798
rect 5910 5795 5966 5798
rect 6018 5795 6074 5798
rect 6126 5795 6836 5798
rect 6888 5795 6944 5798
rect 6996 5795 7052 5798
rect 7104 5795 7160 5798
rect 7212 5795 7268 5798
rect 7320 5795 7376 5798
rect 7428 5795 7484 5798
rect 7536 5795 7592 5798
rect 7644 5795 7700 5798
rect 7752 5795 7808 5798
rect 7860 5795 7916 5798
rect 7968 5795 8024 5798
rect 8076 5795 8132 5798
rect 8184 5795 8240 5798
rect 8292 5795 8348 5798
rect 8400 5795 8456 5798
rect 8508 5795 8564 5798
rect 8616 5795 8672 5798
rect 8724 5795 8780 5798
rect 8832 5795 9206 5798
rect 9258 5795 9314 5798
rect 9366 5795 9422 5798
rect 9474 5795 9530 5798
rect 9582 5795 9638 5798
rect 9690 5795 9746 5798
rect 9798 5795 9854 5798
rect 9906 5795 9962 5798
rect 10014 5795 10070 5798
rect 10122 5795 10178 5798
rect 10230 5795 10286 5798
rect 10338 5795 10394 5798
rect 10446 5795 10502 5798
rect 10554 5795 10610 5798
rect 10662 5795 10718 5798
rect 10770 5795 10826 5798
rect 10878 5795 10934 5798
rect 10986 5795 11042 5798
rect 11094 5795 11150 5798
rect 11202 5795 11481 5798
rect 1481 5783 11481 5795
rect 1481 5603 11481 5615
rect 1481 5551 1493 5603
rect 1545 5600 1601 5603
rect 1653 5600 3863 5603
rect 3915 5600 3971 5603
rect 4023 5600 6239 5603
rect 6291 5600 6347 5603
rect 6399 5600 6455 5603
rect 6507 5600 6563 5603
rect 6615 5600 6671 5603
rect 6723 5600 8939 5603
rect 8991 5600 9047 5603
rect 9099 5600 11309 5603
rect 11361 5600 11417 5603
rect 1545 5551 1601 5554
rect 1653 5551 3863 5554
rect 3915 5551 3971 5554
rect 4023 5551 6239 5554
rect 6291 5551 6347 5554
rect 6399 5551 6455 5554
rect 6507 5551 6563 5554
rect 6615 5551 6671 5554
rect 6723 5551 8939 5554
rect 8991 5551 9047 5554
rect 9099 5551 11309 5554
rect 11361 5551 11417 5554
rect 11469 5551 11481 5603
rect 1481 5539 11481 5551
rect 1481 5359 11481 5371
rect 1481 5356 1760 5359
rect 1812 5356 1868 5359
rect 1920 5356 1976 5359
rect 2028 5356 2084 5359
rect 2136 5356 2192 5359
rect 2244 5356 2300 5359
rect 2352 5356 2408 5359
rect 2460 5356 2516 5359
rect 2568 5356 2624 5359
rect 2676 5356 2732 5359
rect 2784 5356 2840 5359
rect 2892 5356 2948 5359
rect 3000 5356 3056 5359
rect 3108 5356 3164 5359
rect 3216 5356 3272 5359
rect 3324 5356 3380 5359
rect 3432 5356 3488 5359
rect 3540 5356 3596 5359
rect 3648 5356 3704 5359
rect 3756 5356 4130 5359
rect 4182 5356 4238 5359
rect 4290 5356 4346 5359
rect 4398 5356 4454 5359
rect 4506 5356 4562 5359
rect 4614 5356 4670 5359
rect 4722 5356 4778 5359
rect 4830 5356 4886 5359
rect 4938 5356 4994 5359
rect 5046 5356 5102 5359
rect 5154 5356 5210 5359
rect 5262 5356 5318 5359
rect 5370 5356 5426 5359
rect 5478 5356 5534 5359
rect 5586 5356 5642 5359
rect 5694 5356 5750 5359
rect 5802 5356 5858 5359
rect 5910 5356 5966 5359
rect 6018 5356 6074 5359
rect 6126 5356 6836 5359
rect 6888 5356 6944 5359
rect 6996 5356 7052 5359
rect 7104 5356 7160 5359
rect 7212 5356 7268 5359
rect 7320 5356 7376 5359
rect 7428 5356 7484 5359
rect 7536 5356 7592 5359
rect 7644 5356 7700 5359
rect 7752 5356 7808 5359
rect 7860 5356 7916 5359
rect 7968 5356 8024 5359
rect 8076 5356 8132 5359
rect 8184 5356 8240 5359
rect 8292 5356 8348 5359
rect 8400 5356 8456 5359
rect 8508 5356 8564 5359
rect 8616 5356 8672 5359
rect 8724 5356 8780 5359
rect 8832 5356 9206 5359
rect 9258 5356 9314 5359
rect 9366 5356 9422 5359
rect 9474 5356 9530 5359
rect 9582 5356 9638 5359
rect 9690 5356 9746 5359
rect 9798 5356 9854 5359
rect 9906 5356 9962 5359
rect 10014 5356 10070 5359
rect 10122 5356 10178 5359
rect 10230 5356 10286 5359
rect 10338 5356 10394 5359
rect 10446 5356 10502 5359
rect 10554 5356 10610 5359
rect 10662 5356 10718 5359
rect 10770 5356 10826 5359
rect 10878 5356 10934 5359
rect 10986 5356 11042 5359
rect 11094 5356 11150 5359
rect 11202 5356 11481 5359
rect 1481 5310 1494 5356
rect 11468 5310 11481 5356
rect 1481 5307 1760 5310
rect 1812 5307 1868 5310
rect 1920 5307 1976 5310
rect 2028 5307 2084 5310
rect 2136 5307 2192 5310
rect 2244 5307 2300 5310
rect 2352 5307 2408 5310
rect 2460 5307 2516 5310
rect 2568 5307 2624 5310
rect 2676 5307 2732 5310
rect 2784 5307 2840 5310
rect 2892 5307 2948 5310
rect 3000 5307 3056 5310
rect 3108 5307 3164 5310
rect 3216 5307 3272 5310
rect 3324 5307 3380 5310
rect 3432 5307 3488 5310
rect 3540 5307 3596 5310
rect 3648 5307 3704 5310
rect 3756 5307 4130 5310
rect 4182 5307 4238 5310
rect 4290 5307 4346 5310
rect 4398 5307 4454 5310
rect 4506 5307 4562 5310
rect 4614 5307 4670 5310
rect 4722 5307 4778 5310
rect 4830 5307 4886 5310
rect 4938 5307 4994 5310
rect 5046 5307 5102 5310
rect 5154 5307 5210 5310
rect 5262 5307 5318 5310
rect 5370 5307 5426 5310
rect 5478 5307 5534 5310
rect 5586 5307 5642 5310
rect 5694 5307 5750 5310
rect 5802 5307 5858 5310
rect 5910 5307 5966 5310
rect 6018 5307 6074 5310
rect 6126 5307 6836 5310
rect 6888 5307 6944 5310
rect 6996 5307 7052 5310
rect 7104 5307 7160 5310
rect 7212 5307 7268 5310
rect 7320 5307 7376 5310
rect 7428 5307 7484 5310
rect 7536 5307 7592 5310
rect 7644 5307 7700 5310
rect 7752 5307 7808 5310
rect 7860 5307 7916 5310
rect 7968 5307 8024 5310
rect 8076 5307 8132 5310
rect 8184 5307 8240 5310
rect 8292 5307 8348 5310
rect 8400 5307 8456 5310
rect 8508 5307 8564 5310
rect 8616 5307 8672 5310
rect 8724 5307 8780 5310
rect 8832 5307 9206 5310
rect 9258 5307 9314 5310
rect 9366 5307 9422 5310
rect 9474 5307 9530 5310
rect 9582 5307 9638 5310
rect 9690 5307 9746 5310
rect 9798 5307 9854 5310
rect 9906 5307 9962 5310
rect 10014 5307 10070 5310
rect 10122 5307 10178 5310
rect 10230 5307 10286 5310
rect 10338 5307 10394 5310
rect 10446 5307 10502 5310
rect 10554 5307 10610 5310
rect 10662 5307 10718 5310
rect 10770 5307 10826 5310
rect 10878 5307 10934 5310
rect 10986 5307 11042 5310
rect 11094 5307 11150 5310
rect 11202 5307 11481 5310
rect 1481 5295 11481 5307
rect 1481 5115 11481 5127
rect 1481 5063 1493 5115
rect 1545 5112 1601 5115
rect 1653 5112 3863 5115
rect 3915 5112 3971 5115
rect 4023 5112 6239 5115
rect 6291 5112 6347 5115
rect 6399 5112 6455 5115
rect 6507 5112 6563 5115
rect 6615 5112 6671 5115
rect 6723 5112 8939 5115
rect 8991 5112 9047 5115
rect 9099 5112 11309 5115
rect 11361 5112 11417 5115
rect 1545 5063 1601 5066
rect 1653 5063 3863 5066
rect 3915 5063 3971 5066
rect 4023 5063 6239 5066
rect 6291 5063 6347 5066
rect 6399 5063 6455 5066
rect 6507 5063 6563 5066
rect 6615 5063 6671 5066
rect 6723 5063 8939 5066
rect 8991 5063 9047 5066
rect 9099 5063 11309 5066
rect 11361 5063 11417 5066
rect 11469 5063 11481 5115
rect 1481 5051 11481 5063
rect 1481 4871 11481 4883
rect 1481 4868 1760 4871
rect 1812 4868 1868 4871
rect 1920 4868 1976 4871
rect 2028 4868 2084 4871
rect 2136 4868 2192 4871
rect 2244 4868 2300 4871
rect 2352 4868 2408 4871
rect 2460 4868 2516 4871
rect 2568 4868 2624 4871
rect 2676 4868 2732 4871
rect 2784 4868 2840 4871
rect 2892 4868 2948 4871
rect 3000 4868 3056 4871
rect 3108 4868 3164 4871
rect 3216 4868 3272 4871
rect 3324 4868 3380 4871
rect 3432 4868 3488 4871
rect 3540 4868 3596 4871
rect 3648 4868 3704 4871
rect 3756 4868 4130 4871
rect 4182 4868 4238 4871
rect 4290 4868 4346 4871
rect 4398 4868 4454 4871
rect 4506 4868 4562 4871
rect 4614 4868 4670 4871
rect 4722 4868 4778 4871
rect 4830 4868 4886 4871
rect 4938 4868 4994 4871
rect 5046 4868 5102 4871
rect 5154 4868 5210 4871
rect 5262 4868 5318 4871
rect 5370 4868 5426 4871
rect 5478 4868 5534 4871
rect 5586 4868 5642 4871
rect 5694 4868 5750 4871
rect 5802 4868 5858 4871
rect 5910 4868 5966 4871
rect 6018 4868 6074 4871
rect 6126 4868 6836 4871
rect 6888 4868 6944 4871
rect 6996 4868 7052 4871
rect 7104 4868 7160 4871
rect 7212 4868 7268 4871
rect 7320 4868 7376 4871
rect 7428 4868 7484 4871
rect 7536 4868 7592 4871
rect 7644 4868 7700 4871
rect 7752 4868 7808 4871
rect 7860 4868 7916 4871
rect 7968 4868 8024 4871
rect 8076 4868 8132 4871
rect 8184 4868 8240 4871
rect 8292 4868 8348 4871
rect 8400 4868 8456 4871
rect 8508 4868 8564 4871
rect 8616 4868 8672 4871
rect 8724 4868 8780 4871
rect 8832 4868 9206 4871
rect 9258 4868 9314 4871
rect 9366 4868 9422 4871
rect 9474 4868 9530 4871
rect 9582 4868 9638 4871
rect 9690 4868 9746 4871
rect 9798 4868 9854 4871
rect 9906 4868 9962 4871
rect 10014 4868 10070 4871
rect 10122 4868 10178 4871
rect 10230 4868 10286 4871
rect 10338 4868 10394 4871
rect 10446 4868 10502 4871
rect 10554 4868 10610 4871
rect 10662 4868 10718 4871
rect 10770 4868 10826 4871
rect 10878 4868 10934 4871
rect 10986 4868 11042 4871
rect 11094 4868 11150 4871
rect 11202 4868 11481 4871
rect 1481 4822 1494 4868
rect 11468 4822 11481 4868
rect 1481 4819 1760 4822
rect 1812 4819 1868 4822
rect 1920 4819 1976 4822
rect 2028 4819 2084 4822
rect 2136 4819 2192 4822
rect 2244 4819 2300 4822
rect 2352 4819 2408 4822
rect 2460 4819 2516 4822
rect 2568 4819 2624 4822
rect 2676 4819 2732 4822
rect 2784 4819 2840 4822
rect 2892 4819 2948 4822
rect 3000 4819 3056 4822
rect 3108 4819 3164 4822
rect 3216 4819 3272 4822
rect 3324 4819 3380 4822
rect 3432 4819 3488 4822
rect 3540 4819 3596 4822
rect 3648 4819 3704 4822
rect 3756 4819 4130 4822
rect 4182 4819 4238 4822
rect 4290 4819 4346 4822
rect 4398 4819 4454 4822
rect 4506 4819 4562 4822
rect 4614 4819 4670 4822
rect 4722 4819 4778 4822
rect 4830 4819 4886 4822
rect 4938 4819 4994 4822
rect 5046 4819 5102 4822
rect 5154 4819 5210 4822
rect 5262 4819 5318 4822
rect 5370 4819 5426 4822
rect 5478 4819 5534 4822
rect 5586 4819 5642 4822
rect 5694 4819 5750 4822
rect 5802 4819 5858 4822
rect 5910 4819 5966 4822
rect 6018 4819 6074 4822
rect 6126 4819 6836 4822
rect 6888 4819 6944 4822
rect 6996 4819 7052 4822
rect 7104 4819 7160 4822
rect 7212 4819 7268 4822
rect 7320 4819 7376 4822
rect 7428 4819 7484 4822
rect 7536 4819 7592 4822
rect 7644 4819 7700 4822
rect 7752 4819 7808 4822
rect 7860 4819 7916 4822
rect 7968 4819 8024 4822
rect 8076 4819 8132 4822
rect 8184 4819 8240 4822
rect 8292 4819 8348 4822
rect 8400 4819 8456 4822
rect 8508 4819 8564 4822
rect 8616 4819 8672 4822
rect 8724 4819 8780 4822
rect 8832 4819 9206 4822
rect 9258 4819 9314 4822
rect 9366 4819 9422 4822
rect 9474 4819 9530 4822
rect 9582 4819 9638 4822
rect 9690 4819 9746 4822
rect 9798 4819 9854 4822
rect 9906 4819 9962 4822
rect 10014 4819 10070 4822
rect 10122 4819 10178 4822
rect 10230 4819 10286 4822
rect 10338 4819 10394 4822
rect 10446 4819 10502 4822
rect 10554 4819 10610 4822
rect 10662 4819 10718 4822
rect 10770 4819 10826 4822
rect 10878 4819 10934 4822
rect 10986 4819 11042 4822
rect 11094 4819 11150 4822
rect 11202 4819 11481 4822
rect 1481 4807 11481 4819
rect 1481 4627 11481 4639
rect 1481 4575 1493 4627
rect 1545 4624 1601 4627
rect 1653 4624 3863 4627
rect 3915 4624 3971 4627
rect 4023 4624 6239 4627
rect 6291 4624 6347 4627
rect 6399 4624 6455 4627
rect 6507 4624 6563 4627
rect 6615 4624 6671 4627
rect 6723 4624 8939 4627
rect 8991 4624 9047 4627
rect 9099 4624 11309 4627
rect 11361 4624 11417 4627
rect 1545 4575 1601 4578
rect 1653 4575 3863 4578
rect 3915 4575 3971 4578
rect 4023 4575 6239 4578
rect 6291 4575 6347 4578
rect 6399 4575 6455 4578
rect 6507 4575 6563 4578
rect 6615 4575 6671 4578
rect 6723 4575 8939 4578
rect 8991 4575 9047 4578
rect 9099 4575 11309 4578
rect 11361 4575 11417 4578
rect 11469 4575 11481 4627
rect 1481 4563 11481 4575
rect 1481 4383 11481 4395
rect 1481 4380 1760 4383
rect 1812 4380 1868 4383
rect 1920 4380 1976 4383
rect 2028 4380 2084 4383
rect 2136 4380 2192 4383
rect 2244 4380 2300 4383
rect 2352 4380 2408 4383
rect 2460 4380 2516 4383
rect 2568 4380 2624 4383
rect 2676 4380 2732 4383
rect 2784 4380 2840 4383
rect 2892 4380 2948 4383
rect 3000 4380 3056 4383
rect 3108 4380 3164 4383
rect 3216 4380 3272 4383
rect 3324 4380 3380 4383
rect 3432 4380 3488 4383
rect 3540 4380 3596 4383
rect 3648 4380 3704 4383
rect 3756 4380 4130 4383
rect 4182 4380 4238 4383
rect 4290 4380 4346 4383
rect 4398 4380 4454 4383
rect 4506 4380 4562 4383
rect 4614 4380 4670 4383
rect 4722 4380 4778 4383
rect 4830 4380 4886 4383
rect 4938 4380 4994 4383
rect 5046 4380 5102 4383
rect 5154 4380 5210 4383
rect 5262 4380 5318 4383
rect 5370 4380 5426 4383
rect 5478 4380 5534 4383
rect 5586 4380 5642 4383
rect 5694 4380 5750 4383
rect 5802 4380 5858 4383
rect 5910 4380 5966 4383
rect 6018 4380 6074 4383
rect 6126 4380 6836 4383
rect 6888 4380 6944 4383
rect 6996 4380 7052 4383
rect 7104 4380 7160 4383
rect 7212 4380 7268 4383
rect 7320 4380 7376 4383
rect 7428 4380 7484 4383
rect 7536 4380 7592 4383
rect 7644 4380 7700 4383
rect 7752 4380 7808 4383
rect 7860 4380 7916 4383
rect 7968 4380 8024 4383
rect 8076 4380 8132 4383
rect 8184 4380 8240 4383
rect 8292 4380 8348 4383
rect 8400 4380 8456 4383
rect 8508 4380 8564 4383
rect 8616 4380 8672 4383
rect 8724 4380 8780 4383
rect 8832 4380 9206 4383
rect 9258 4380 9314 4383
rect 9366 4380 9422 4383
rect 9474 4380 9530 4383
rect 9582 4380 9638 4383
rect 9690 4380 9746 4383
rect 9798 4380 9854 4383
rect 9906 4380 9962 4383
rect 10014 4380 10070 4383
rect 10122 4380 10178 4383
rect 10230 4380 10286 4383
rect 10338 4380 10394 4383
rect 10446 4380 10502 4383
rect 10554 4380 10610 4383
rect 10662 4380 10718 4383
rect 10770 4380 10826 4383
rect 10878 4380 10934 4383
rect 10986 4380 11042 4383
rect 11094 4380 11150 4383
rect 11202 4380 11481 4383
rect 1481 4334 1494 4380
rect 11468 4334 11481 4380
rect 1481 4331 1760 4334
rect 1812 4331 1868 4334
rect 1920 4331 1976 4334
rect 2028 4331 2084 4334
rect 2136 4331 2192 4334
rect 2244 4331 2300 4334
rect 2352 4331 2408 4334
rect 2460 4331 2516 4334
rect 2568 4331 2624 4334
rect 2676 4331 2732 4334
rect 2784 4331 2840 4334
rect 2892 4331 2948 4334
rect 3000 4331 3056 4334
rect 3108 4331 3164 4334
rect 3216 4331 3272 4334
rect 3324 4331 3380 4334
rect 3432 4331 3488 4334
rect 3540 4331 3596 4334
rect 3648 4331 3704 4334
rect 3756 4331 4130 4334
rect 4182 4331 4238 4334
rect 4290 4331 4346 4334
rect 4398 4331 4454 4334
rect 4506 4331 4562 4334
rect 4614 4331 4670 4334
rect 4722 4331 4778 4334
rect 4830 4331 4886 4334
rect 4938 4331 4994 4334
rect 5046 4331 5102 4334
rect 5154 4331 5210 4334
rect 5262 4331 5318 4334
rect 5370 4331 5426 4334
rect 5478 4331 5534 4334
rect 5586 4331 5642 4334
rect 5694 4331 5750 4334
rect 5802 4331 5858 4334
rect 5910 4331 5966 4334
rect 6018 4331 6074 4334
rect 6126 4331 6836 4334
rect 6888 4331 6944 4334
rect 6996 4331 7052 4334
rect 7104 4331 7160 4334
rect 7212 4331 7268 4334
rect 7320 4331 7376 4334
rect 7428 4331 7484 4334
rect 7536 4331 7592 4334
rect 7644 4331 7700 4334
rect 7752 4331 7808 4334
rect 7860 4331 7916 4334
rect 7968 4331 8024 4334
rect 8076 4331 8132 4334
rect 8184 4331 8240 4334
rect 8292 4331 8348 4334
rect 8400 4331 8456 4334
rect 8508 4331 8564 4334
rect 8616 4331 8672 4334
rect 8724 4331 8780 4334
rect 8832 4331 9206 4334
rect 9258 4331 9314 4334
rect 9366 4331 9422 4334
rect 9474 4331 9530 4334
rect 9582 4331 9638 4334
rect 9690 4331 9746 4334
rect 9798 4331 9854 4334
rect 9906 4331 9962 4334
rect 10014 4331 10070 4334
rect 10122 4331 10178 4334
rect 10230 4331 10286 4334
rect 10338 4331 10394 4334
rect 10446 4331 10502 4334
rect 10554 4331 10610 4334
rect 10662 4331 10718 4334
rect 10770 4331 10826 4334
rect 10878 4331 10934 4334
rect 10986 4331 11042 4334
rect 11094 4331 11150 4334
rect 11202 4331 11481 4334
rect 1481 4319 11481 4331
rect 1481 4139 11481 4151
rect 1481 4087 1493 4139
rect 1545 4136 1601 4139
rect 1653 4136 3863 4139
rect 3915 4136 3971 4139
rect 4023 4136 6239 4139
rect 6291 4136 6347 4139
rect 6399 4136 6455 4139
rect 6507 4136 6563 4139
rect 6615 4136 6671 4139
rect 6723 4136 8939 4139
rect 8991 4136 9047 4139
rect 9099 4136 11309 4139
rect 11361 4136 11417 4139
rect 1545 4087 1601 4090
rect 1653 4087 3863 4090
rect 3915 4087 3971 4090
rect 4023 4087 6239 4090
rect 6291 4087 6347 4090
rect 6399 4087 6455 4090
rect 6507 4087 6563 4090
rect 6615 4087 6671 4090
rect 6723 4087 8939 4090
rect 8991 4087 9047 4090
rect 9099 4087 11309 4090
rect 11361 4087 11417 4090
rect 11469 4087 11481 4139
rect 1481 4075 11481 4087
rect 1481 3895 11481 3907
rect 1481 3892 1760 3895
rect 1812 3892 1868 3895
rect 1920 3892 1976 3895
rect 2028 3892 2084 3895
rect 2136 3892 2192 3895
rect 2244 3892 2300 3895
rect 2352 3892 2408 3895
rect 2460 3892 2516 3895
rect 2568 3892 2624 3895
rect 2676 3892 2732 3895
rect 2784 3892 2840 3895
rect 2892 3892 2948 3895
rect 3000 3892 3056 3895
rect 3108 3892 3164 3895
rect 3216 3892 3272 3895
rect 3324 3892 3380 3895
rect 3432 3892 3488 3895
rect 3540 3892 3596 3895
rect 3648 3892 3704 3895
rect 3756 3892 4130 3895
rect 4182 3892 4238 3895
rect 4290 3892 4346 3895
rect 4398 3892 4454 3895
rect 4506 3892 4562 3895
rect 4614 3892 4670 3895
rect 4722 3892 4778 3895
rect 4830 3892 4886 3895
rect 4938 3892 4994 3895
rect 5046 3892 5102 3895
rect 5154 3892 5210 3895
rect 5262 3892 5318 3895
rect 5370 3892 5426 3895
rect 5478 3892 5534 3895
rect 5586 3892 5642 3895
rect 5694 3892 5750 3895
rect 5802 3892 5858 3895
rect 5910 3892 5966 3895
rect 6018 3892 6074 3895
rect 6126 3892 6836 3895
rect 6888 3892 6944 3895
rect 6996 3892 7052 3895
rect 7104 3892 7160 3895
rect 7212 3892 7268 3895
rect 7320 3892 7376 3895
rect 7428 3892 7484 3895
rect 7536 3892 7592 3895
rect 7644 3892 7700 3895
rect 7752 3892 7808 3895
rect 7860 3892 7916 3895
rect 7968 3892 8024 3895
rect 8076 3892 8132 3895
rect 8184 3892 8240 3895
rect 8292 3892 8348 3895
rect 8400 3892 8456 3895
rect 8508 3892 8564 3895
rect 8616 3892 8672 3895
rect 8724 3892 8780 3895
rect 8832 3892 9206 3895
rect 9258 3892 9314 3895
rect 9366 3892 9422 3895
rect 9474 3892 9530 3895
rect 9582 3892 9638 3895
rect 9690 3892 9746 3895
rect 9798 3892 9854 3895
rect 9906 3892 9962 3895
rect 10014 3892 10070 3895
rect 10122 3892 10178 3895
rect 10230 3892 10286 3895
rect 10338 3892 10394 3895
rect 10446 3892 10502 3895
rect 10554 3892 10610 3895
rect 10662 3892 10718 3895
rect 10770 3892 10826 3895
rect 10878 3892 10934 3895
rect 10986 3892 11042 3895
rect 11094 3892 11150 3895
rect 11202 3892 11481 3895
rect 1481 3846 1494 3892
rect 11468 3846 11481 3892
rect 1481 3843 1760 3846
rect 1812 3843 1868 3846
rect 1920 3843 1976 3846
rect 2028 3843 2084 3846
rect 2136 3843 2192 3846
rect 2244 3843 2300 3846
rect 2352 3843 2408 3846
rect 2460 3843 2516 3846
rect 2568 3843 2624 3846
rect 2676 3843 2732 3846
rect 2784 3843 2840 3846
rect 2892 3843 2948 3846
rect 3000 3843 3056 3846
rect 3108 3843 3164 3846
rect 3216 3843 3272 3846
rect 3324 3843 3380 3846
rect 3432 3843 3488 3846
rect 3540 3843 3596 3846
rect 3648 3843 3704 3846
rect 3756 3843 4130 3846
rect 4182 3843 4238 3846
rect 4290 3843 4346 3846
rect 4398 3843 4454 3846
rect 4506 3843 4562 3846
rect 4614 3843 4670 3846
rect 4722 3843 4778 3846
rect 4830 3843 4886 3846
rect 4938 3843 4994 3846
rect 5046 3843 5102 3846
rect 5154 3843 5210 3846
rect 5262 3843 5318 3846
rect 5370 3843 5426 3846
rect 5478 3843 5534 3846
rect 5586 3843 5642 3846
rect 5694 3843 5750 3846
rect 5802 3843 5858 3846
rect 5910 3843 5966 3846
rect 6018 3843 6074 3846
rect 6126 3843 6836 3846
rect 6888 3843 6944 3846
rect 6996 3843 7052 3846
rect 7104 3843 7160 3846
rect 7212 3843 7268 3846
rect 7320 3843 7376 3846
rect 7428 3843 7484 3846
rect 7536 3843 7592 3846
rect 7644 3843 7700 3846
rect 7752 3843 7808 3846
rect 7860 3843 7916 3846
rect 7968 3843 8024 3846
rect 8076 3843 8132 3846
rect 8184 3843 8240 3846
rect 8292 3843 8348 3846
rect 8400 3843 8456 3846
rect 8508 3843 8564 3846
rect 8616 3843 8672 3846
rect 8724 3843 8780 3846
rect 8832 3843 9206 3846
rect 9258 3843 9314 3846
rect 9366 3843 9422 3846
rect 9474 3843 9530 3846
rect 9582 3843 9638 3846
rect 9690 3843 9746 3846
rect 9798 3843 9854 3846
rect 9906 3843 9962 3846
rect 10014 3843 10070 3846
rect 10122 3843 10178 3846
rect 10230 3843 10286 3846
rect 10338 3843 10394 3846
rect 10446 3843 10502 3846
rect 10554 3843 10610 3846
rect 10662 3843 10718 3846
rect 10770 3843 10826 3846
rect 10878 3843 10934 3846
rect 10986 3843 11042 3846
rect 11094 3843 11150 3846
rect 11202 3843 11481 3846
rect 1481 3831 11481 3843
rect 1481 3651 11481 3663
rect 1481 3599 1493 3651
rect 1545 3648 1601 3651
rect 1653 3648 3863 3651
rect 3915 3648 3971 3651
rect 4023 3648 6239 3651
rect 6291 3648 6347 3651
rect 6399 3648 6455 3651
rect 6507 3648 6563 3651
rect 6615 3648 6671 3651
rect 6723 3648 8939 3651
rect 8991 3648 9047 3651
rect 9099 3648 11309 3651
rect 11361 3648 11417 3651
rect 1545 3599 1601 3602
rect 1653 3599 3863 3602
rect 3915 3599 3971 3602
rect 4023 3599 6239 3602
rect 6291 3599 6347 3602
rect 6399 3599 6455 3602
rect 6507 3599 6563 3602
rect 6615 3599 6671 3602
rect 6723 3599 8939 3602
rect 8991 3599 9047 3602
rect 9099 3599 11309 3602
rect 11361 3599 11417 3602
rect 11469 3599 11481 3651
rect 1481 3587 11481 3599
rect 1481 3407 11481 3419
rect 1481 3404 1760 3407
rect 1812 3404 1868 3407
rect 1920 3404 1976 3407
rect 2028 3404 2084 3407
rect 2136 3404 2192 3407
rect 2244 3404 2300 3407
rect 2352 3404 2408 3407
rect 2460 3404 2516 3407
rect 2568 3404 2624 3407
rect 2676 3404 2732 3407
rect 2784 3404 2840 3407
rect 2892 3404 2948 3407
rect 3000 3404 3056 3407
rect 3108 3404 3164 3407
rect 3216 3404 3272 3407
rect 3324 3404 3380 3407
rect 3432 3404 3488 3407
rect 3540 3404 3596 3407
rect 3648 3404 3704 3407
rect 3756 3404 4130 3407
rect 4182 3404 4238 3407
rect 4290 3404 4346 3407
rect 4398 3404 4454 3407
rect 4506 3404 4562 3407
rect 4614 3404 4670 3407
rect 4722 3404 4778 3407
rect 4830 3404 4886 3407
rect 4938 3404 4994 3407
rect 5046 3404 5102 3407
rect 5154 3404 5210 3407
rect 5262 3404 5318 3407
rect 5370 3404 5426 3407
rect 5478 3404 5534 3407
rect 5586 3404 5642 3407
rect 5694 3404 5750 3407
rect 5802 3404 5858 3407
rect 5910 3404 5966 3407
rect 6018 3404 6074 3407
rect 6126 3404 6836 3407
rect 6888 3404 6944 3407
rect 6996 3404 7052 3407
rect 7104 3404 7160 3407
rect 7212 3404 7268 3407
rect 7320 3404 7376 3407
rect 7428 3404 7484 3407
rect 7536 3404 7592 3407
rect 7644 3404 7700 3407
rect 7752 3404 7808 3407
rect 7860 3404 7916 3407
rect 7968 3404 8024 3407
rect 8076 3404 8132 3407
rect 8184 3404 8240 3407
rect 8292 3404 8348 3407
rect 8400 3404 8456 3407
rect 8508 3404 8564 3407
rect 8616 3404 8672 3407
rect 8724 3404 8780 3407
rect 8832 3404 9206 3407
rect 9258 3404 9314 3407
rect 9366 3404 9422 3407
rect 9474 3404 9530 3407
rect 9582 3404 9638 3407
rect 9690 3404 9746 3407
rect 9798 3404 9854 3407
rect 9906 3404 9962 3407
rect 10014 3404 10070 3407
rect 10122 3404 10178 3407
rect 10230 3404 10286 3407
rect 10338 3404 10394 3407
rect 10446 3404 10502 3407
rect 10554 3404 10610 3407
rect 10662 3404 10718 3407
rect 10770 3404 10826 3407
rect 10878 3404 10934 3407
rect 10986 3404 11042 3407
rect 11094 3404 11150 3407
rect 11202 3404 11481 3407
rect 1481 3358 1494 3404
rect 11468 3358 11481 3404
rect 1481 3355 1760 3358
rect 1812 3355 1868 3358
rect 1920 3355 1976 3358
rect 2028 3355 2084 3358
rect 2136 3355 2192 3358
rect 2244 3355 2300 3358
rect 2352 3355 2408 3358
rect 2460 3355 2516 3358
rect 2568 3355 2624 3358
rect 2676 3355 2732 3358
rect 2784 3355 2840 3358
rect 2892 3355 2948 3358
rect 3000 3355 3056 3358
rect 3108 3355 3164 3358
rect 3216 3355 3272 3358
rect 3324 3355 3380 3358
rect 3432 3355 3488 3358
rect 3540 3355 3596 3358
rect 3648 3355 3704 3358
rect 3756 3355 4130 3358
rect 4182 3355 4238 3358
rect 4290 3355 4346 3358
rect 4398 3355 4454 3358
rect 4506 3355 4562 3358
rect 4614 3355 4670 3358
rect 4722 3355 4778 3358
rect 4830 3355 4886 3358
rect 4938 3355 4994 3358
rect 5046 3355 5102 3358
rect 5154 3355 5210 3358
rect 5262 3355 5318 3358
rect 5370 3355 5426 3358
rect 5478 3355 5534 3358
rect 5586 3355 5642 3358
rect 5694 3355 5750 3358
rect 5802 3355 5858 3358
rect 5910 3355 5966 3358
rect 6018 3355 6074 3358
rect 6126 3355 6836 3358
rect 6888 3355 6944 3358
rect 6996 3355 7052 3358
rect 7104 3355 7160 3358
rect 7212 3355 7268 3358
rect 7320 3355 7376 3358
rect 7428 3355 7484 3358
rect 7536 3355 7592 3358
rect 7644 3355 7700 3358
rect 7752 3355 7808 3358
rect 7860 3355 7916 3358
rect 7968 3355 8024 3358
rect 8076 3355 8132 3358
rect 8184 3355 8240 3358
rect 8292 3355 8348 3358
rect 8400 3355 8456 3358
rect 8508 3355 8564 3358
rect 8616 3355 8672 3358
rect 8724 3355 8780 3358
rect 8832 3355 9206 3358
rect 9258 3355 9314 3358
rect 9366 3355 9422 3358
rect 9474 3355 9530 3358
rect 9582 3355 9638 3358
rect 9690 3355 9746 3358
rect 9798 3355 9854 3358
rect 9906 3355 9962 3358
rect 10014 3355 10070 3358
rect 10122 3355 10178 3358
rect 10230 3355 10286 3358
rect 10338 3355 10394 3358
rect 10446 3355 10502 3358
rect 10554 3355 10610 3358
rect 10662 3355 10718 3358
rect 10770 3355 10826 3358
rect 10878 3355 10934 3358
rect 10986 3355 11042 3358
rect 11094 3355 11150 3358
rect 11202 3355 11481 3358
rect 1481 3343 11481 3355
rect 1481 3163 11481 3175
rect 1481 3111 1493 3163
rect 1545 3160 1601 3163
rect 1653 3160 3863 3163
rect 3915 3160 3971 3163
rect 4023 3160 6239 3163
rect 6291 3160 6347 3163
rect 6399 3160 6455 3163
rect 6507 3160 6563 3163
rect 6615 3160 6671 3163
rect 6723 3160 8939 3163
rect 8991 3160 9047 3163
rect 9099 3160 11309 3163
rect 11361 3160 11417 3163
rect 1545 3111 1601 3114
rect 1653 3111 3863 3114
rect 3915 3111 3971 3114
rect 4023 3111 6239 3114
rect 6291 3111 6347 3114
rect 6399 3111 6455 3114
rect 6507 3111 6563 3114
rect 6615 3111 6671 3114
rect 6723 3111 8939 3114
rect 8991 3111 9047 3114
rect 9099 3111 11309 3114
rect 11361 3111 11417 3114
rect 11469 3111 11481 3163
rect 1481 3099 11481 3111
rect 1481 2919 11481 2931
rect 1481 2916 1760 2919
rect 1812 2916 1868 2919
rect 1920 2916 1976 2919
rect 2028 2916 2084 2919
rect 2136 2916 2192 2919
rect 2244 2916 2300 2919
rect 2352 2916 2408 2919
rect 2460 2916 2516 2919
rect 2568 2916 2624 2919
rect 2676 2916 2732 2919
rect 2784 2916 2840 2919
rect 2892 2916 2948 2919
rect 3000 2916 3056 2919
rect 3108 2916 3164 2919
rect 3216 2916 3272 2919
rect 3324 2916 3380 2919
rect 3432 2916 3488 2919
rect 3540 2916 3596 2919
rect 3648 2916 3704 2919
rect 3756 2916 4130 2919
rect 4182 2916 4238 2919
rect 4290 2916 4346 2919
rect 4398 2916 4454 2919
rect 4506 2916 4562 2919
rect 4614 2916 4670 2919
rect 4722 2916 4778 2919
rect 4830 2916 4886 2919
rect 4938 2916 4994 2919
rect 5046 2916 5102 2919
rect 5154 2916 5210 2919
rect 5262 2916 5318 2919
rect 5370 2916 5426 2919
rect 5478 2916 5534 2919
rect 5586 2916 5642 2919
rect 5694 2916 5750 2919
rect 5802 2916 5858 2919
rect 5910 2916 5966 2919
rect 6018 2916 6074 2919
rect 6126 2916 6836 2919
rect 6888 2916 6944 2919
rect 6996 2916 7052 2919
rect 7104 2916 7160 2919
rect 7212 2916 7268 2919
rect 7320 2916 7376 2919
rect 7428 2916 7484 2919
rect 7536 2916 7592 2919
rect 7644 2916 7700 2919
rect 7752 2916 7808 2919
rect 7860 2916 7916 2919
rect 7968 2916 8024 2919
rect 8076 2916 8132 2919
rect 8184 2916 8240 2919
rect 8292 2916 8348 2919
rect 8400 2916 8456 2919
rect 8508 2916 8564 2919
rect 8616 2916 8672 2919
rect 8724 2916 8780 2919
rect 8832 2916 9206 2919
rect 9258 2916 9314 2919
rect 9366 2916 9422 2919
rect 9474 2916 9530 2919
rect 9582 2916 9638 2919
rect 9690 2916 9746 2919
rect 9798 2916 9854 2919
rect 9906 2916 9962 2919
rect 10014 2916 10070 2919
rect 10122 2916 10178 2919
rect 10230 2916 10286 2919
rect 10338 2916 10394 2919
rect 10446 2916 10502 2919
rect 10554 2916 10610 2919
rect 10662 2916 10718 2919
rect 10770 2916 10826 2919
rect 10878 2916 10934 2919
rect 10986 2916 11042 2919
rect 11094 2916 11150 2919
rect 11202 2916 11481 2919
rect 1481 2870 1494 2916
rect 11468 2870 11481 2916
rect 1481 2867 1760 2870
rect 1812 2867 1868 2870
rect 1920 2867 1976 2870
rect 2028 2867 2084 2870
rect 2136 2867 2192 2870
rect 2244 2867 2300 2870
rect 2352 2867 2408 2870
rect 2460 2867 2516 2870
rect 2568 2867 2624 2870
rect 2676 2867 2732 2870
rect 2784 2867 2840 2870
rect 2892 2867 2948 2870
rect 3000 2867 3056 2870
rect 3108 2867 3164 2870
rect 3216 2867 3272 2870
rect 3324 2867 3380 2870
rect 3432 2867 3488 2870
rect 3540 2867 3596 2870
rect 3648 2867 3704 2870
rect 3756 2867 4130 2870
rect 4182 2867 4238 2870
rect 4290 2867 4346 2870
rect 4398 2867 4454 2870
rect 4506 2867 4562 2870
rect 4614 2867 4670 2870
rect 4722 2867 4778 2870
rect 4830 2867 4886 2870
rect 4938 2867 4994 2870
rect 5046 2867 5102 2870
rect 5154 2867 5210 2870
rect 5262 2867 5318 2870
rect 5370 2867 5426 2870
rect 5478 2867 5534 2870
rect 5586 2867 5642 2870
rect 5694 2867 5750 2870
rect 5802 2867 5858 2870
rect 5910 2867 5966 2870
rect 6018 2867 6074 2870
rect 6126 2867 6836 2870
rect 6888 2867 6944 2870
rect 6996 2867 7052 2870
rect 7104 2867 7160 2870
rect 7212 2867 7268 2870
rect 7320 2867 7376 2870
rect 7428 2867 7484 2870
rect 7536 2867 7592 2870
rect 7644 2867 7700 2870
rect 7752 2867 7808 2870
rect 7860 2867 7916 2870
rect 7968 2867 8024 2870
rect 8076 2867 8132 2870
rect 8184 2867 8240 2870
rect 8292 2867 8348 2870
rect 8400 2867 8456 2870
rect 8508 2867 8564 2870
rect 8616 2867 8672 2870
rect 8724 2867 8780 2870
rect 8832 2867 9206 2870
rect 9258 2867 9314 2870
rect 9366 2867 9422 2870
rect 9474 2867 9530 2870
rect 9582 2867 9638 2870
rect 9690 2867 9746 2870
rect 9798 2867 9854 2870
rect 9906 2867 9962 2870
rect 10014 2867 10070 2870
rect 10122 2867 10178 2870
rect 10230 2867 10286 2870
rect 10338 2867 10394 2870
rect 10446 2867 10502 2870
rect 10554 2867 10610 2870
rect 10662 2867 10718 2870
rect 10770 2867 10826 2870
rect 10878 2867 10934 2870
rect 10986 2867 11042 2870
rect 11094 2867 11150 2870
rect 11202 2867 11481 2870
rect 1481 2855 11481 2867
rect 1481 2675 11481 2687
rect 1481 2623 1493 2675
rect 1545 2672 1601 2675
rect 1653 2672 3863 2675
rect 3915 2672 3971 2675
rect 4023 2672 6239 2675
rect 6291 2672 6347 2675
rect 6399 2672 6455 2675
rect 6507 2672 6563 2675
rect 6615 2672 6671 2675
rect 6723 2672 8939 2675
rect 8991 2672 9047 2675
rect 9099 2672 11309 2675
rect 11361 2672 11417 2675
rect 1545 2623 1601 2626
rect 1653 2623 3863 2626
rect 3915 2623 3971 2626
rect 4023 2623 6239 2626
rect 6291 2623 6347 2626
rect 6399 2623 6455 2626
rect 6507 2623 6563 2626
rect 6615 2623 6671 2626
rect 6723 2623 8939 2626
rect 8991 2623 9047 2626
rect 9099 2623 11309 2626
rect 11361 2623 11417 2626
rect 11469 2623 11481 2675
rect 1481 2611 11481 2623
rect 1481 2431 11481 2443
rect 1481 2428 1760 2431
rect 1812 2428 1868 2431
rect 1920 2428 1976 2431
rect 2028 2428 2084 2431
rect 2136 2428 2192 2431
rect 2244 2428 2300 2431
rect 2352 2428 2408 2431
rect 2460 2428 2516 2431
rect 2568 2428 2624 2431
rect 2676 2428 2732 2431
rect 2784 2428 2840 2431
rect 2892 2428 2948 2431
rect 3000 2428 3056 2431
rect 3108 2428 3164 2431
rect 3216 2428 3272 2431
rect 3324 2428 3380 2431
rect 3432 2428 3488 2431
rect 3540 2428 3596 2431
rect 3648 2428 3704 2431
rect 3756 2428 4130 2431
rect 4182 2428 4238 2431
rect 4290 2428 4346 2431
rect 4398 2428 4454 2431
rect 4506 2428 4562 2431
rect 4614 2428 4670 2431
rect 4722 2428 4778 2431
rect 4830 2428 4886 2431
rect 4938 2428 4994 2431
rect 5046 2428 5102 2431
rect 5154 2428 5210 2431
rect 5262 2428 5318 2431
rect 5370 2428 5426 2431
rect 5478 2428 5534 2431
rect 5586 2428 5642 2431
rect 5694 2428 5750 2431
rect 5802 2428 5858 2431
rect 5910 2428 5966 2431
rect 6018 2428 6074 2431
rect 6126 2428 6836 2431
rect 6888 2428 6944 2431
rect 6996 2428 7052 2431
rect 7104 2428 7160 2431
rect 7212 2428 7268 2431
rect 7320 2428 7376 2431
rect 7428 2428 7484 2431
rect 7536 2428 7592 2431
rect 7644 2428 7700 2431
rect 7752 2428 7808 2431
rect 7860 2428 7916 2431
rect 7968 2428 8024 2431
rect 8076 2428 8132 2431
rect 8184 2428 8240 2431
rect 8292 2428 8348 2431
rect 8400 2428 8456 2431
rect 8508 2428 8564 2431
rect 8616 2428 8672 2431
rect 8724 2428 8780 2431
rect 8832 2428 9206 2431
rect 9258 2428 9314 2431
rect 9366 2428 9422 2431
rect 9474 2428 9530 2431
rect 9582 2428 9638 2431
rect 9690 2428 9746 2431
rect 9798 2428 9854 2431
rect 9906 2428 9962 2431
rect 10014 2428 10070 2431
rect 10122 2428 10178 2431
rect 10230 2428 10286 2431
rect 10338 2428 10394 2431
rect 10446 2428 10502 2431
rect 10554 2428 10610 2431
rect 10662 2428 10718 2431
rect 10770 2428 10826 2431
rect 10878 2428 10934 2431
rect 10986 2428 11042 2431
rect 11094 2428 11150 2431
rect 11202 2428 11481 2431
rect 1481 2382 1494 2428
rect 11468 2382 11481 2428
rect 1481 2379 1760 2382
rect 1812 2379 1868 2382
rect 1920 2379 1976 2382
rect 2028 2379 2084 2382
rect 2136 2379 2192 2382
rect 2244 2379 2300 2382
rect 2352 2379 2408 2382
rect 2460 2379 2516 2382
rect 2568 2379 2624 2382
rect 2676 2379 2732 2382
rect 2784 2379 2840 2382
rect 2892 2379 2948 2382
rect 3000 2379 3056 2382
rect 3108 2379 3164 2382
rect 3216 2379 3272 2382
rect 3324 2379 3380 2382
rect 3432 2379 3488 2382
rect 3540 2379 3596 2382
rect 3648 2379 3704 2382
rect 3756 2379 4130 2382
rect 4182 2379 4238 2382
rect 4290 2379 4346 2382
rect 4398 2379 4454 2382
rect 4506 2379 4562 2382
rect 4614 2379 4670 2382
rect 4722 2379 4778 2382
rect 4830 2379 4886 2382
rect 4938 2379 4994 2382
rect 5046 2379 5102 2382
rect 5154 2379 5210 2382
rect 5262 2379 5318 2382
rect 5370 2379 5426 2382
rect 5478 2379 5534 2382
rect 5586 2379 5642 2382
rect 5694 2379 5750 2382
rect 5802 2379 5858 2382
rect 5910 2379 5966 2382
rect 6018 2379 6074 2382
rect 6126 2379 6836 2382
rect 6888 2379 6944 2382
rect 6996 2379 7052 2382
rect 7104 2379 7160 2382
rect 7212 2379 7268 2382
rect 7320 2379 7376 2382
rect 7428 2379 7484 2382
rect 7536 2379 7592 2382
rect 7644 2379 7700 2382
rect 7752 2379 7808 2382
rect 7860 2379 7916 2382
rect 7968 2379 8024 2382
rect 8076 2379 8132 2382
rect 8184 2379 8240 2382
rect 8292 2379 8348 2382
rect 8400 2379 8456 2382
rect 8508 2379 8564 2382
rect 8616 2379 8672 2382
rect 8724 2379 8780 2382
rect 8832 2379 9206 2382
rect 9258 2379 9314 2382
rect 9366 2379 9422 2382
rect 9474 2379 9530 2382
rect 9582 2379 9638 2382
rect 9690 2379 9746 2382
rect 9798 2379 9854 2382
rect 9906 2379 9962 2382
rect 10014 2379 10070 2382
rect 10122 2379 10178 2382
rect 10230 2379 10286 2382
rect 10338 2379 10394 2382
rect 10446 2379 10502 2382
rect 10554 2379 10610 2382
rect 10662 2379 10718 2382
rect 10770 2379 10826 2382
rect 10878 2379 10934 2382
rect 10986 2379 11042 2382
rect 11094 2379 11150 2382
rect 11202 2379 11481 2382
rect 1481 2367 11481 2379
rect 1481 2187 11481 2199
rect 1481 2135 1493 2187
rect 1545 2184 1601 2187
rect 1653 2184 3863 2187
rect 3915 2184 3971 2187
rect 4023 2184 6239 2187
rect 6291 2184 6347 2187
rect 6399 2184 6455 2187
rect 6507 2184 6563 2187
rect 6615 2184 6671 2187
rect 6723 2184 8939 2187
rect 8991 2184 9047 2187
rect 9099 2184 11309 2187
rect 11361 2184 11417 2187
rect 1545 2135 1601 2138
rect 1653 2135 3863 2138
rect 3915 2135 3971 2138
rect 4023 2135 6239 2138
rect 6291 2135 6347 2138
rect 6399 2135 6455 2138
rect 6507 2135 6563 2138
rect 6615 2135 6671 2138
rect 6723 2135 8939 2138
rect 8991 2135 9047 2138
rect 9099 2135 11309 2138
rect 11361 2135 11417 2138
rect 11469 2135 11481 2187
rect 1481 2123 11481 2135
rect 1481 1943 11481 1955
rect 1481 1940 1760 1943
rect 1812 1940 1868 1943
rect 1920 1940 1976 1943
rect 2028 1940 2084 1943
rect 2136 1940 2192 1943
rect 2244 1940 2300 1943
rect 2352 1940 2408 1943
rect 2460 1940 2516 1943
rect 2568 1940 2624 1943
rect 2676 1940 2732 1943
rect 2784 1940 2840 1943
rect 2892 1940 2948 1943
rect 3000 1940 3056 1943
rect 3108 1940 3164 1943
rect 3216 1940 3272 1943
rect 3324 1940 3380 1943
rect 3432 1940 3488 1943
rect 3540 1940 3596 1943
rect 3648 1940 3704 1943
rect 3756 1940 4130 1943
rect 4182 1940 4238 1943
rect 4290 1940 4346 1943
rect 4398 1940 4454 1943
rect 4506 1940 4562 1943
rect 4614 1940 4670 1943
rect 4722 1940 4778 1943
rect 4830 1940 4886 1943
rect 4938 1940 4994 1943
rect 5046 1940 5102 1943
rect 5154 1940 5210 1943
rect 5262 1940 5318 1943
rect 5370 1940 5426 1943
rect 5478 1940 5534 1943
rect 5586 1940 5642 1943
rect 5694 1940 5750 1943
rect 5802 1940 5858 1943
rect 5910 1940 5966 1943
rect 6018 1940 6074 1943
rect 6126 1940 6836 1943
rect 6888 1940 6944 1943
rect 6996 1940 7052 1943
rect 7104 1940 7160 1943
rect 7212 1940 7268 1943
rect 7320 1940 7376 1943
rect 7428 1940 7484 1943
rect 7536 1940 7592 1943
rect 7644 1940 7700 1943
rect 7752 1940 7808 1943
rect 7860 1940 7916 1943
rect 7968 1940 8024 1943
rect 8076 1940 8132 1943
rect 8184 1940 8240 1943
rect 8292 1940 8348 1943
rect 8400 1940 8456 1943
rect 8508 1940 8564 1943
rect 8616 1940 8672 1943
rect 8724 1940 8780 1943
rect 8832 1940 9206 1943
rect 9258 1940 9314 1943
rect 9366 1940 9422 1943
rect 9474 1940 9530 1943
rect 9582 1940 9638 1943
rect 9690 1940 9746 1943
rect 9798 1940 9854 1943
rect 9906 1940 9962 1943
rect 10014 1940 10070 1943
rect 10122 1940 10178 1943
rect 10230 1940 10286 1943
rect 10338 1940 10394 1943
rect 10446 1940 10502 1943
rect 10554 1940 10610 1943
rect 10662 1940 10718 1943
rect 10770 1940 10826 1943
rect 10878 1940 10934 1943
rect 10986 1940 11042 1943
rect 11094 1940 11150 1943
rect 11202 1940 11481 1943
rect 1481 1894 1494 1940
rect 11468 1894 11481 1940
rect 1481 1891 1760 1894
rect 1812 1891 1868 1894
rect 1920 1891 1976 1894
rect 2028 1891 2084 1894
rect 2136 1891 2192 1894
rect 2244 1891 2300 1894
rect 2352 1891 2408 1894
rect 2460 1891 2516 1894
rect 2568 1891 2624 1894
rect 2676 1891 2732 1894
rect 2784 1891 2840 1894
rect 2892 1891 2948 1894
rect 3000 1891 3056 1894
rect 3108 1891 3164 1894
rect 3216 1891 3272 1894
rect 3324 1891 3380 1894
rect 3432 1891 3488 1894
rect 3540 1891 3596 1894
rect 3648 1891 3704 1894
rect 3756 1891 4130 1894
rect 4182 1891 4238 1894
rect 4290 1891 4346 1894
rect 4398 1891 4454 1894
rect 4506 1891 4562 1894
rect 4614 1891 4670 1894
rect 4722 1891 4778 1894
rect 4830 1891 4886 1894
rect 4938 1891 4994 1894
rect 5046 1891 5102 1894
rect 5154 1891 5210 1894
rect 5262 1891 5318 1894
rect 5370 1891 5426 1894
rect 5478 1891 5534 1894
rect 5586 1891 5642 1894
rect 5694 1891 5750 1894
rect 5802 1891 5858 1894
rect 5910 1891 5966 1894
rect 6018 1891 6074 1894
rect 6126 1891 6836 1894
rect 6888 1891 6944 1894
rect 6996 1891 7052 1894
rect 7104 1891 7160 1894
rect 7212 1891 7268 1894
rect 7320 1891 7376 1894
rect 7428 1891 7484 1894
rect 7536 1891 7592 1894
rect 7644 1891 7700 1894
rect 7752 1891 7808 1894
rect 7860 1891 7916 1894
rect 7968 1891 8024 1894
rect 8076 1891 8132 1894
rect 8184 1891 8240 1894
rect 8292 1891 8348 1894
rect 8400 1891 8456 1894
rect 8508 1891 8564 1894
rect 8616 1891 8672 1894
rect 8724 1891 8780 1894
rect 8832 1891 9206 1894
rect 9258 1891 9314 1894
rect 9366 1891 9422 1894
rect 9474 1891 9530 1894
rect 9582 1891 9638 1894
rect 9690 1891 9746 1894
rect 9798 1891 9854 1894
rect 9906 1891 9962 1894
rect 10014 1891 10070 1894
rect 10122 1891 10178 1894
rect 10230 1891 10286 1894
rect 10338 1891 10394 1894
rect 10446 1891 10502 1894
rect 10554 1891 10610 1894
rect 10662 1891 10718 1894
rect 10770 1891 10826 1894
rect 10878 1891 10934 1894
rect 10986 1891 11042 1894
rect 11094 1891 11150 1894
rect 11202 1891 11481 1894
rect 1481 1879 11481 1891
rect 1481 1699 11481 1711
rect 1481 1647 1493 1699
rect 1545 1696 1601 1699
rect 1653 1696 3863 1699
rect 3915 1696 3971 1699
rect 4023 1696 6239 1699
rect 6291 1696 6347 1699
rect 6399 1696 6455 1699
rect 6507 1696 6563 1699
rect 6615 1696 6671 1699
rect 6723 1696 8939 1699
rect 8991 1696 9047 1699
rect 9099 1696 11309 1699
rect 11361 1696 11417 1699
rect 1545 1647 1601 1650
rect 1653 1647 3863 1650
rect 3915 1647 3971 1650
rect 4023 1647 6239 1650
rect 6291 1647 6347 1650
rect 6399 1647 6455 1650
rect 6507 1647 6563 1650
rect 6615 1647 6671 1650
rect 6723 1647 8939 1650
rect 8991 1647 9047 1650
rect 9099 1647 11309 1650
rect 11361 1647 11417 1650
rect 11469 1647 11481 1699
rect 1481 1635 11481 1647
rect 1213 1519 1413 1546
rect 1213 1467 1233 1519
rect 1285 1467 1341 1519
rect 1393 1467 1413 1519
rect 11549 1546 11560 6192
rect 11706 6163 11749 6192
rect 11729 6111 11749 6163
rect 11706 6055 11749 6111
rect 11729 6003 11749 6055
rect 11706 5947 11749 6003
rect 11729 5895 11749 5947
rect 11706 5839 11749 5895
rect 11729 5787 11749 5839
rect 11706 5731 11749 5787
rect 11729 5679 11749 5731
rect 11706 5623 11749 5679
rect 11729 5571 11749 5623
rect 11706 5515 11749 5571
rect 11729 5463 11749 5515
rect 11706 5407 11749 5463
rect 11729 5355 11749 5407
rect 11706 5299 11749 5355
rect 11729 5247 11749 5299
rect 11706 5191 11749 5247
rect 11729 5139 11749 5191
rect 11706 5083 11749 5139
rect 11729 5031 11749 5083
rect 11706 4975 11749 5031
rect 11729 4923 11749 4975
rect 11706 4867 11749 4923
rect 11729 4815 11749 4867
rect 11706 4759 11749 4815
rect 11729 4707 11749 4759
rect 11706 4651 11749 4707
rect 11729 4599 11749 4651
rect 11706 4543 11749 4599
rect 11729 4491 11749 4543
rect 11706 4435 11749 4491
rect 11729 4383 11749 4435
rect 11706 4327 11749 4383
rect 11729 4275 11749 4327
rect 11706 4219 11749 4275
rect 11729 4167 11749 4219
rect 11706 4111 11749 4167
rect 11729 4059 11749 4111
rect 11706 4003 11749 4059
rect 11729 3951 11749 4003
rect 11706 3895 11749 3951
rect 11729 3843 11749 3895
rect 11706 3787 11749 3843
rect 11729 3735 11749 3787
rect 11706 3679 11749 3735
rect 11729 3627 11749 3679
rect 11706 3571 11749 3627
rect 11729 3519 11749 3571
rect 11706 3463 11749 3519
rect 11729 3411 11749 3463
rect 11706 3355 11749 3411
rect 11729 3303 11749 3355
rect 11706 3247 11749 3303
rect 11729 3195 11749 3247
rect 11706 3139 11749 3195
rect 11729 3087 11749 3139
rect 11706 3031 11749 3087
rect 11729 2979 11749 3031
rect 11706 2923 11749 2979
rect 11729 2871 11749 2923
rect 11706 2815 11749 2871
rect 11729 2763 11749 2815
rect 11706 2707 11749 2763
rect 11729 2655 11749 2707
rect 11706 2599 11749 2655
rect 11729 2547 11749 2599
rect 11706 2491 11749 2547
rect 11729 2439 11749 2491
rect 11706 2383 11749 2439
rect 11729 2331 11749 2383
rect 11706 2275 11749 2331
rect 11729 2223 11749 2275
rect 11706 2167 11749 2223
rect 11729 2115 11749 2167
rect 11706 2059 11749 2115
rect 11729 2007 11749 2059
rect 11706 1951 11749 2007
rect 11729 1899 11749 1951
rect 11706 1843 11749 1899
rect 11729 1791 11749 1843
rect 11706 1735 11749 1791
rect 11729 1683 11749 1735
rect 11706 1627 11749 1683
rect 11729 1575 11749 1627
rect 11706 1546 11749 1575
rect 11549 1519 11749 1546
rect 11549 1467 11569 1519
rect 11621 1467 11677 1519
rect 11729 1467 11749 1519
rect 1213 1298 1413 1467
rect 1481 1455 11481 1467
rect 1481 1452 1760 1455
rect 1812 1452 1868 1455
rect 1920 1452 1976 1455
rect 2028 1452 2084 1455
rect 2136 1452 2192 1455
rect 2244 1452 2300 1455
rect 2352 1452 2408 1455
rect 2460 1452 2516 1455
rect 2568 1452 2624 1455
rect 2676 1452 2732 1455
rect 2784 1452 2840 1455
rect 2892 1452 2948 1455
rect 3000 1452 3056 1455
rect 3108 1452 3164 1455
rect 3216 1452 3272 1455
rect 3324 1452 3380 1455
rect 3432 1452 3488 1455
rect 3540 1452 3596 1455
rect 3648 1452 3704 1455
rect 3756 1452 4130 1455
rect 4182 1452 4238 1455
rect 4290 1452 4346 1455
rect 4398 1452 4454 1455
rect 4506 1452 4562 1455
rect 4614 1452 4670 1455
rect 4722 1452 4778 1455
rect 4830 1452 4886 1455
rect 4938 1452 4994 1455
rect 5046 1452 5102 1455
rect 5154 1452 5210 1455
rect 5262 1452 5318 1455
rect 5370 1452 5426 1455
rect 5478 1452 5534 1455
rect 5586 1452 5642 1455
rect 5694 1452 5750 1455
rect 5802 1452 5858 1455
rect 5910 1452 5966 1455
rect 6018 1452 6074 1455
rect 6126 1452 6836 1455
rect 6888 1452 6944 1455
rect 6996 1452 7052 1455
rect 7104 1452 7160 1455
rect 7212 1452 7268 1455
rect 7320 1452 7376 1455
rect 7428 1452 7484 1455
rect 7536 1452 7592 1455
rect 7644 1452 7700 1455
rect 7752 1452 7808 1455
rect 7860 1452 7916 1455
rect 7968 1452 8024 1455
rect 8076 1452 8132 1455
rect 8184 1452 8240 1455
rect 8292 1452 8348 1455
rect 8400 1452 8456 1455
rect 8508 1452 8564 1455
rect 8616 1452 8672 1455
rect 8724 1452 8780 1455
rect 8832 1452 9206 1455
rect 9258 1452 9314 1455
rect 9366 1452 9422 1455
rect 9474 1452 9530 1455
rect 9582 1452 9638 1455
rect 9690 1452 9746 1455
rect 9798 1452 9854 1455
rect 9906 1452 9962 1455
rect 10014 1452 10070 1455
rect 10122 1452 10178 1455
rect 10230 1452 10286 1455
rect 10338 1452 10394 1455
rect 10446 1452 10502 1455
rect 10554 1452 10610 1455
rect 10662 1452 10718 1455
rect 10770 1452 10826 1455
rect 10878 1452 10934 1455
rect 10986 1452 11042 1455
rect 11094 1452 11150 1455
rect 11202 1452 11481 1455
rect 1481 1406 1494 1452
rect 11468 1406 11481 1452
rect 1481 1403 1760 1406
rect 1812 1403 1868 1406
rect 1920 1403 1976 1406
rect 2028 1403 2084 1406
rect 2136 1403 2192 1406
rect 2244 1403 2300 1406
rect 2352 1403 2408 1406
rect 2460 1403 2516 1406
rect 2568 1403 2624 1406
rect 2676 1403 2732 1406
rect 2784 1403 2840 1406
rect 2892 1403 2948 1406
rect 3000 1403 3056 1406
rect 3108 1403 3164 1406
rect 3216 1403 3272 1406
rect 3324 1403 3380 1406
rect 3432 1403 3488 1406
rect 3540 1403 3596 1406
rect 3648 1403 3704 1406
rect 3756 1403 4130 1406
rect 4182 1403 4238 1406
rect 4290 1403 4346 1406
rect 4398 1403 4454 1406
rect 4506 1403 4562 1406
rect 4614 1403 4670 1406
rect 4722 1403 4778 1406
rect 4830 1403 4886 1406
rect 4938 1403 4994 1406
rect 5046 1403 5102 1406
rect 5154 1403 5210 1406
rect 5262 1403 5318 1406
rect 5370 1403 5426 1406
rect 5478 1403 5534 1406
rect 5586 1403 5642 1406
rect 5694 1403 5750 1406
rect 5802 1403 5858 1406
rect 5910 1403 5966 1406
rect 6018 1403 6074 1406
rect 6126 1403 6836 1406
rect 6888 1403 6944 1406
rect 6996 1403 7052 1406
rect 7104 1403 7160 1406
rect 7212 1403 7268 1406
rect 7320 1403 7376 1406
rect 7428 1403 7484 1406
rect 7536 1403 7592 1406
rect 7644 1403 7700 1406
rect 7752 1403 7808 1406
rect 7860 1403 7916 1406
rect 7968 1403 8024 1406
rect 8076 1403 8132 1406
rect 8184 1403 8240 1406
rect 8292 1403 8348 1406
rect 8400 1403 8456 1406
rect 8508 1403 8564 1406
rect 8616 1403 8672 1406
rect 8724 1403 8780 1406
rect 8832 1403 9206 1406
rect 9258 1403 9314 1406
rect 9366 1403 9422 1406
rect 9474 1403 9530 1406
rect 9582 1403 9638 1406
rect 9690 1403 9746 1406
rect 9798 1403 9854 1406
rect 9906 1403 9962 1406
rect 10014 1403 10070 1406
rect 10122 1403 10178 1406
rect 10230 1403 10286 1406
rect 10338 1403 10394 1406
rect 10446 1403 10502 1406
rect 10554 1403 10610 1406
rect 10662 1403 10718 1406
rect 10770 1403 10826 1406
rect 10878 1403 10934 1406
rect 10986 1403 11042 1406
rect 11094 1403 11150 1406
rect 11202 1403 11481 1406
rect 1481 1391 11481 1403
rect 11549 1298 11749 1467
rect 1213 1098 11749 1298
rect 12001 1011 12012 6713
rect 950 1000 12012 1011
rect 950 654 1058 1000
rect 11904 654 12012 1000
rect 12358 654 12369 24700
rect 593 643 12369 654
rect 12551 411 12562 24943
rect 400 400 12562 411
rect 400 54 508 400
rect 12454 54 12562 400
rect 12908 54 12919 25300
rect 43 43 12919 54
<< via1 >>
rect 1493 25209 1545 25261
rect 1601 25209 1653 25261
rect 3863 25209 3915 25261
rect 3971 25209 4023 25261
rect 6239 25209 6291 25261
rect 6347 25209 6399 25261
rect 6455 25209 6507 25261
rect 6563 25209 6615 25261
rect 6671 25209 6723 25261
rect 8939 25209 8991 25261
rect 9047 25209 9099 25261
rect 11309 25209 11361 25261
rect 11417 25209 11469 25261
rect 1493 25101 1545 25153
rect 1601 25101 1653 25153
rect 3863 25101 3915 25153
rect 3971 25101 4023 25153
rect 6239 25101 6291 25153
rect 6347 25101 6399 25153
rect 6455 25101 6507 25153
rect 6563 25101 6615 25153
rect 6671 25101 6723 25153
rect 8939 25101 8991 25153
rect 9047 25101 9099 25153
rect 11309 25101 11361 25153
rect 11417 25101 11469 25153
rect 1493 24993 1545 25045
rect 1601 24993 1653 25045
rect 3863 24993 3915 25045
rect 3971 24993 4023 25045
rect 6239 24993 6291 25045
rect 6347 24993 6399 25045
rect 6455 24993 6507 25045
rect 6563 24993 6615 25045
rect 6671 24993 6723 25045
rect 8939 24993 8991 25045
rect 9047 24993 9099 25045
rect 11309 24993 11361 25045
rect 11417 24993 11469 25045
rect 643 24639 695 24691
rect 751 24639 803 24691
rect 859 24639 911 24691
rect 643 24531 695 24583
rect 751 24531 803 24583
rect 859 24531 911 24583
rect 643 24423 695 24475
rect 751 24423 803 24475
rect 859 24423 911 24475
rect 643 24315 695 24367
rect 751 24315 803 24367
rect 859 24315 911 24367
rect 1760 24609 1812 24661
rect 1868 24609 1920 24661
rect 1976 24609 2028 24661
rect 2084 24609 2136 24661
rect 2192 24609 2244 24661
rect 2300 24609 2352 24661
rect 2408 24609 2460 24661
rect 2516 24609 2568 24661
rect 2624 24609 2676 24661
rect 2732 24609 2784 24661
rect 2840 24609 2892 24661
rect 2948 24609 3000 24661
rect 3056 24609 3108 24661
rect 3164 24609 3216 24661
rect 3272 24609 3324 24661
rect 3380 24609 3432 24661
rect 3488 24609 3540 24661
rect 3596 24609 3648 24661
rect 3704 24609 3756 24661
rect 4130 24609 4182 24661
rect 4238 24609 4290 24661
rect 4346 24609 4398 24661
rect 4454 24609 4506 24661
rect 4562 24609 4614 24661
rect 4670 24609 4722 24661
rect 4778 24609 4830 24661
rect 4886 24609 4938 24661
rect 4994 24609 5046 24661
rect 5102 24609 5154 24661
rect 5210 24609 5262 24661
rect 5318 24609 5370 24661
rect 5426 24609 5478 24661
rect 5534 24609 5586 24661
rect 5642 24609 5694 24661
rect 5750 24609 5802 24661
rect 5858 24609 5910 24661
rect 5966 24609 6018 24661
rect 6074 24609 6126 24661
rect 6836 24609 6888 24661
rect 6944 24609 6996 24661
rect 7052 24609 7104 24661
rect 7160 24609 7212 24661
rect 7268 24609 7320 24661
rect 7376 24609 7428 24661
rect 7484 24609 7536 24661
rect 7592 24609 7644 24661
rect 7700 24609 7752 24661
rect 7808 24609 7860 24661
rect 7916 24609 7968 24661
rect 8024 24609 8076 24661
rect 8132 24609 8184 24661
rect 8240 24609 8292 24661
rect 8348 24609 8400 24661
rect 8456 24609 8508 24661
rect 8564 24609 8616 24661
rect 8672 24609 8724 24661
rect 8780 24609 8832 24661
rect 9206 24609 9258 24661
rect 9314 24609 9366 24661
rect 9422 24609 9474 24661
rect 9530 24609 9582 24661
rect 9638 24609 9690 24661
rect 9746 24609 9798 24661
rect 9854 24609 9906 24661
rect 9962 24609 10014 24661
rect 10070 24609 10122 24661
rect 10178 24609 10230 24661
rect 10286 24609 10338 24661
rect 10394 24609 10446 24661
rect 10502 24609 10554 24661
rect 10610 24609 10662 24661
rect 10718 24609 10770 24661
rect 10826 24609 10878 24661
rect 10934 24609 10986 24661
rect 11042 24609 11094 24661
rect 11150 24609 11202 24661
rect 1760 24501 1812 24553
rect 1868 24501 1920 24553
rect 1976 24501 2028 24553
rect 2084 24501 2136 24553
rect 2192 24501 2244 24553
rect 2300 24501 2352 24553
rect 2408 24501 2460 24553
rect 2516 24501 2568 24553
rect 2624 24501 2676 24553
rect 2732 24501 2784 24553
rect 2840 24501 2892 24553
rect 2948 24501 3000 24553
rect 3056 24501 3108 24553
rect 3164 24501 3216 24553
rect 3272 24501 3324 24553
rect 3380 24501 3432 24553
rect 3488 24501 3540 24553
rect 3596 24501 3648 24553
rect 3704 24501 3756 24553
rect 4130 24501 4182 24553
rect 4238 24501 4290 24553
rect 4346 24501 4398 24553
rect 4454 24501 4506 24553
rect 4562 24501 4614 24553
rect 4670 24501 4722 24553
rect 4778 24501 4830 24553
rect 4886 24501 4938 24553
rect 4994 24501 5046 24553
rect 5102 24501 5154 24553
rect 5210 24501 5262 24553
rect 5318 24501 5370 24553
rect 5426 24501 5478 24553
rect 5534 24501 5586 24553
rect 5642 24501 5694 24553
rect 5750 24501 5802 24553
rect 5858 24501 5910 24553
rect 5966 24501 6018 24553
rect 6074 24501 6126 24553
rect 6836 24501 6888 24553
rect 6944 24501 6996 24553
rect 7052 24501 7104 24553
rect 7160 24501 7212 24553
rect 7268 24501 7320 24553
rect 7376 24501 7428 24553
rect 7484 24501 7536 24553
rect 7592 24501 7644 24553
rect 7700 24501 7752 24553
rect 7808 24501 7860 24553
rect 7916 24501 7968 24553
rect 8024 24501 8076 24553
rect 8132 24501 8184 24553
rect 8240 24501 8292 24553
rect 8348 24501 8400 24553
rect 8456 24501 8508 24553
rect 8564 24501 8616 24553
rect 8672 24501 8724 24553
rect 8780 24501 8832 24553
rect 9206 24501 9258 24553
rect 9314 24501 9366 24553
rect 9422 24501 9474 24553
rect 9530 24501 9582 24553
rect 9638 24501 9690 24553
rect 9746 24501 9798 24553
rect 9854 24501 9906 24553
rect 9962 24501 10014 24553
rect 10070 24501 10122 24553
rect 10178 24501 10230 24553
rect 10286 24501 10338 24553
rect 10394 24501 10446 24553
rect 10502 24501 10554 24553
rect 10610 24501 10662 24553
rect 10718 24501 10770 24553
rect 10826 24501 10878 24553
rect 10934 24501 10986 24553
rect 11042 24501 11094 24553
rect 11150 24501 11202 24553
rect 1760 24393 1812 24445
rect 1868 24393 1920 24445
rect 1976 24393 2028 24445
rect 2084 24393 2136 24445
rect 2192 24393 2244 24445
rect 2300 24393 2352 24445
rect 2408 24393 2460 24445
rect 2516 24393 2568 24445
rect 2624 24393 2676 24445
rect 2732 24393 2784 24445
rect 2840 24393 2892 24445
rect 2948 24393 3000 24445
rect 3056 24393 3108 24445
rect 3164 24393 3216 24445
rect 3272 24393 3324 24445
rect 3380 24393 3432 24445
rect 3488 24393 3540 24445
rect 3596 24393 3648 24445
rect 3704 24393 3756 24445
rect 4130 24393 4182 24445
rect 4238 24393 4290 24445
rect 4346 24393 4398 24445
rect 4454 24393 4506 24445
rect 4562 24393 4614 24445
rect 4670 24393 4722 24445
rect 4778 24393 4830 24445
rect 4886 24393 4938 24445
rect 4994 24393 5046 24445
rect 5102 24393 5154 24445
rect 5210 24393 5262 24445
rect 5318 24393 5370 24445
rect 5426 24393 5478 24445
rect 5534 24393 5586 24445
rect 5642 24393 5694 24445
rect 5750 24393 5802 24445
rect 5858 24393 5910 24445
rect 5966 24393 6018 24445
rect 6074 24393 6126 24445
rect 6836 24393 6888 24445
rect 6944 24393 6996 24445
rect 7052 24393 7104 24445
rect 7160 24393 7212 24445
rect 7268 24393 7320 24445
rect 7376 24393 7428 24445
rect 7484 24393 7536 24445
rect 7592 24393 7644 24445
rect 7700 24393 7752 24445
rect 7808 24393 7860 24445
rect 7916 24393 7968 24445
rect 8024 24393 8076 24445
rect 8132 24393 8184 24445
rect 8240 24393 8292 24445
rect 8348 24393 8400 24445
rect 8456 24393 8508 24445
rect 8564 24393 8616 24445
rect 8672 24393 8724 24445
rect 8780 24393 8832 24445
rect 9206 24393 9258 24445
rect 9314 24393 9366 24445
rect 9422 24393 9474 24445
rect 9530 24393 9582 24445
rect 9638 24393 9690 24445
rect 9746 24393 9798 24445
rect 9854 24393 9906 24445
rect 9962 24393 10014 24445
rect 10070 24393 10122 24445
rect 10178 24393 10230 24445
rect 10286 24393 10338 24445
rect 10394 24393 10446 24445
rect 10502 24393 10554 24445
rect 10610 24393 10662 24445
rect 10718 24393 10770 24445
rect 10826 24393 10878 24445
rect 10934 24393 10986 24445
rect 11042 24393 11094 24445
rect 11150 24393 11202 24445
rect 12051 24639 12103 24691
rect 12159 24639 12211 24691
rect 12267 24639 12319 24691
rect 12051 24531 12103 24583
rect 12159 24531 12211 24583
rect 12267 24531 12319 24583
rect 12051 24423 12103 24475
rect 12159 24423 12211 24475
rect 12267 24423 12319 24475
rect 643 24207 695 24259
rect 751 24207 803 24259
rect 859 24207 911 24259
rect 643 24099 695 24151
rect 751 24099 803 24151
rect 859 24099 911 24151
rect 643 23991 695 24043
rect 751 23991 803 24043
rect 859 23991 911 24043
rect 643 23883 695 23935
rect 751 23883 803 23935
rect 859 23883 911 23935
rect 643 23775 695 23827
rect 751 23775 803 23827
rect 859 23775 911 23827
rect 643 23667 695 23719
rect 751 23667 803 23719
rect 859 23667 911 23719
rect 643 23559 695 23611
rect 751 23559 803 23611
rect 859 23559 911 23611
rect 643 23451 695 23503
rect 751 23451 803 23503
rect 859 23451 911 23503
rect 643 23343 695 23395
rect 751 23343 803 23395
rect 859 23343 911 23395
rect 643 23235 695 23287
rect 751 23235 803 23287
rect 859 23235 911 23287
rect 643 23127 695 23179
rect 751 23127 803 23179
rect 859 23127 911 23179
rect 643 23019 695 23071
rect 751 23019 803 23071
rect 859 23019 911 23071
rect 643 22911 695 22963
rect 751 22911 803 22963
rect 859 22911 911 22963
rect 643 22803 695 22855
rect 751 22803 803 22855
rect 859 22803 911 22855
rect 643 22695 695 22747
rect 751 22695 803 22747
rect 859 22695 911 22747
rect 643 22587 695 22639
rect 751 22587 803 22639
rect 859 22587 911 22639
rect 643 22479 695 22531
rect 751 22479 803 22531
rect 859 22479 911 22531
rect 643 22371 695 22423
rect 751 22371 803 22423
rect 859 22371 911 22423
rect 643 22263 695 22315
rect 751 22263 803 22315
rect 859 22263 911 22315
rect 643 22155 695 22207
rect 751 22155 803 22207
rect 859 22155 911 22207
rect 643 22047 695 22099
rect 751 22047 803 22099
rect 859 22047 911 22099
rect 643 21939 695 21991
rect 751 21939 803 21991
rect 859 21939 911 21991
rect 643 21831 695 21883
rect 751 21831 803 21883
rect 859 21831 911 21883
rect 643 21723 695 21775
rect 751 21723 803 21775
rect 859 21723 911 21775
rect 643 21615 695 21667
rect 751 21615 803 21667
rect 859 21615 911 21667
rect 643 21507 695 21559
rect 751 21507 803 21559
rect 859 21507 911 21559
rect 643 21399 695 21451
rect 751 21399 803 21451
rect 859 21399 911 21451
rect 643 21291 695 21343
rect 751 21291 803 21343
rect 859 21291 911 21343
rect 643 21183 695 21235
rect 751 21183 803 21235
rect 859 21183 911 21235
rect 643 21075 695 21127
rect 751 21075 803 21127
rect 859 21075 911 21127
rect 643 20967 695 21019
rect 751 20967 803 21019
rect 859 20967 911 21019
rect 643 20859 695 20911
rect 751 20859 803 20911
rect 859 20859 911 20911
rect 643 20751 695 20803
rect 751 20751 803 20803
rect 859 20751 911 20803
rect 643 20643 695 20695
rect 751 20643 803 20695
rect 859 20643 911 20695
rect 643 20535 695 20587
rect 751 20535 803 20587
rect 859 20535 911 20587
rect 643 20427 695 20479
rect 751 20427 803 20479
rect 859 20427 911 20479
rect 643 20319 695 20371
rect 751 20319 803 20371
rect 859 20319 911 20371
rect 643 20211 695 20263
rect 751 20211 803 20263
rect 859 20211 911 20263
rect 643 20103 695 20155
rect 751 20103 803 20155
rect 859 20103 911 20155
rect 643 19995 695 20047
rect 751 19995 803 20047
rect 859 19995 911 20047
rect 643 19887 695 19939
rect 751 19887 803 19939
rect 859 19887 911 19939
rect 643 19779 695 19831
rect 751 19779 803 19831
rect 859 19779 911 19831
rect 643 19671 695 19723
rect 751 19671 803 19723
rect 859 19671 911 19723
rect 643 19563 695 19615
rect 751 19563 803 19615
rect 859 19563 911 19615
rect 643 19455 695 19507
rect 751 19455 803 19507
rect 859 19455 911 19507
rect 643 19347 695 19399
rect 751 19347 803 19399
rect 859 19347 911 19399
rect 643 19239 695 19291
rect 751 19239 803 19291
rect 859 19239 911 19291
rect 643 19131 695 19183
rect 751 19131 803 19183
rect 859 19131 911 19183
rect 643 19023 695 19075
rect 751 19023 803 19075
rect 859 19023 911 19075
rect 643 18915 695 18967
rect 751 18915 803 18967
rect 859 18915 911 18967
rect 643 18807 695 18859
rect 751 18807 803 18859
rect 859 18807 911 18859
rect 643 18699 695 18751
rect 751 18699 803 18751
rect 859 18699 911 18751
rect 643 18591 695 18643
rect 751 18591 803 18643
rect 859 18591 911 18643
rect 1760 23948 1812 23951
rect 1868 23948 1920 23951
rect 1976 23948 2028 23951
rect 2084 23948 2136 23951
rect 2192 23948 2244 23951
rect 2300 23948 2352 23951
rect 2408 23948 2460 23951
rect 2516 23948 2568 23951
rect 2624 23948 2676 23951
rect 2732 23948 2784 23951
rect 2840 23948 2892 23951
rect 2948 23948 3000 23951
rect 3056 23948 3108 23951
rect 3164 23948 3216 23951
rect 3272 23948 3324 23951
rect 3380 23948 3432 23951
rect 3488 23948 3540 23951
rect 3596 23948 3648 23951
rect 3704 23948 3756 23951
rect 4130 23948 4182 23951
rect 4238 23948 4290 23951
rect 4346 23948 4398 23951
rect 4454 23948 4506 23951
rect 4562 23948 4614 23951
rect 4670 23948 4722 23951
rect 4778 23948 4830 23951
rect 4886 23948 4938 23951
rect 4994 23948 5046 23951
rect 5102 23948 5154 23951
rect 5210 23948 5262 23951
rect 5318 23948 5370 23951
rect 5426 23948 5478 23951
rect 5534 23948 5586 23951
rect 5642 23948 5694 23951
rect 5750 23948 5802 23951
rect 5858 23948 5910 23951
rect 5966 23948 6018 23951
rect 6074 23948 6126 23951
rect 6836 23948 6888 23951
rect 6944 23948 6996 23951
rect 7052 23948 7104 23951
rect 7160 23948 7212 23951
rect 7268 23948 7320 23951
rect 7376 23948 7428 23951
rect 7484 23948 7536 23951
rect 7592 23948 7644 23951
rect 7700 23948 7752 23951
rect 7808 23948 7860 23951
rect 7916 23948 7968 23951
rect 8024 23948 8076 23951
rect 8132 23948 8184 23951
rect 8240 23948 8292 23951
rect 8348 23948 8400 23951
rect 8456 23948 8508 23951
rect 8564 23948 8616 23951
rect 8672 23948 8724 23951
rect 8780 23948 8832 23951
rect 9206 23948 9258 23951
rect 9314 23948 9366 23951
rect 9422 23948 9474 23951
rect 9530 23948 9582 23951
rect 9638 23948 9690 23951
rect 9746 23948 9798 23951
rect 9854 23948 9906 23951
rect 9962 23948 10014 23951
rect 10070 23948 10122 23951
rect 10178 23948 10230 23951
rect 10286 23948 10338 23951
rect 10394 23948 10446 23951
rect 10502 23948 10554 23951
rect 10610 23948 10662 23951
rect 10718 23948 10770 23951
rect 10826 23948 10878 23951
rect 10934 23948 10986 23951
rect 11042 23948 11094 23951
rect 11150 23948 11202 23951
rect 1760 23902 1812 23948
rect 1868 23902 1920 23948
rect 1976 23902 2028 23948
rect 2084 23902 2136 23948
rect 2192 23902 2244 23948
rect 2300 23902 2352 23948
rect 2408 23902 2460 23948
rect 2516 23902 2568 23948
rect 2624 23902 2676 23948
rect 2732 23902 2784 23948
rect 2840 23902 2892 23948
rect 2948 23902 3000 23948
rect 3056 23902 3108 23948
rect 3164 23902 3216 23948
rect 3272 23902 3324 23948
rect 3380 23902 3432 23948
rect 3488 23902 3540 23948
rect 3596 23902 3648 23948
rect 3704 23902 3756 23948
rect 4130 23902 4182 23948
rect 4238 23902 4290 23948
rect 4346 23902 4398 23948
rect 4454 23902 4506 23948
rect 4562 23902 4614 23948
rect 4670 23902 4722 23948
rect 4778 23902 4830 23948
rect 4886 23902 4938 23948
rect 4994 23902 5046 23948
rect 5102 23902 5154 23948
rect 5210 23902 5262 23948
rect 5318 23902 5370 23948
rect 5426 23902 5478 23948
rect 5534 23902 5586 23948
rect 5642 23902 5694 23948
rect 5750 23902 5802 23948
rect 5858 23902 5910 23948
rect 5966 23902 6018 23948
rect 6074 23902 6126 23948
rect 6836 23902 6888 23948
rect 6944 23902 6996 23948
rect 7052 23902 7104 23948
rect 7160 23902 7212 23948
rect 7268 23902 7320 23948
rect 7376 23902 7428 23948
rect 7484 23902 7536 23948
rect 7592 23902 7644 23948
rect 7700 23902 7752 23948
rect 7808 23902 7860 23948
rect 7916 23902 7968 23948
rect 8024 23902 8076 23948
rect 8132 23902 8184 23948
rect 8240 23902 8292 23948
rect 8348 23902 8400 23948
rect 8456 23902 8508 23948
rect 8564 23902 8616 23948
rect 8672 23902 8724 23948
rect 8780 23902 8832 23948
rect 9206 23902 9258 23948
rect 9314 23902 9366 23948
rect 9422 23902 9474 23948
rect 9530 23902 9582 23948
rect 9638 23902 9690 23948
rect 9746 23902 9798 23948
rect 9854 23902 9906 23948
rect 9962 23902 10014 23948
rect 10070 23902 10122 23948
rect 10178 23902 10230 23948
rect 10286 23902 10338 23948
rect 10394 23902 10446 23948
rect 10502 23902 10554 23948
rect 10610 23902 10662 23948
rect 10718 23902 10770 23948
rect 10826 23902 10878 23948
rect 10934 23902 10986 23948
rect 11042 23902 11094 23948
rect 11150 23902 11202 23948
rect 1760 23899 1812 23902
rect 1868 23899 1920 23902
rect 1976 23899 2028 23902
rect 2084 23899 2136 23902
rect 2192 23899 2244 23902
rect 2300 23899 2352 23902
rect 2408 23899 2460 23902
rect 2516 23899 2568 23902
rect 2624 23899 2676 23902
rect 2732 23899 2784 23902
rect 2840 23899 2892 23902
rect 2948 23899 3000 23902
rect 3056 23899 3108 23902
rect 3164 23899 3216 23902
rect 3272 23899 3324 23902
rect 3380 23899 3432 23902
rect 3488 23899 3540 23902
rect 3596 23899 3648 23902
rect 3704 23899 3756 23902
rect 4130 23899 4182 23902
rect 4238 23899 4290 23902
rect 4346 23899 4398 23902
rect 4454 23899 4506 23902
rect 4562 23899 4614 23902
rect 4670 23899 4722 23902
rect 4778 23899 4830 23902
rect 4886 23899 4938 23902
rect 4994 23899 5046 23902
rect 5102 23899 5154 23902
rect 5210 23899 5262 23902
rect 5318 23899 5370 23902
rect 5426 23899 5478 23902
rect 5534 23899 5586 23902
rect 5642 23899 5694 23902
rect 5750 23899 5802 23902
rect 5858 23899 5910 23902
rect 5966 23899 6018 23902
rect 6074 23899 6126 23902
rect 6836 23899 6888 23902
rect 6944 23899 6996 23902
rect 7052 23899 7104 23902
rect 7160 23899 7212 23902
rect 7268 23899 7320 23902
rect 7376 23899 7428 23902
rect 7484 23899 7536 23902
rect 7592 23899 7644 23902
rect 7700 23899 7752 23902
rect 7808 23899 7860 23902
rect 7916 23899 7968 23902
rect 8024 23899 8076 23902
rect 8132 23899 8184 23902
rect 8240 23899 8292 23902
rect 8348 23899 8400 23902
rect 8456 23899 8508 23902
rect 8564 23899 8616 23902
rect 8672 23899 8724 23902
rect 8780 23899 8832 23902
rect 9206 23899 9258 23902
rect 9314 23899 9366 23902
rect 9422 23899 9474 23902
rect 9530 23899 9582 23902
rect 9638 23899 9690 23902
rect 9746 23899 9798 23902
rect 9854 23899 9906 23902
rect 9962 23899 10014 23902
rect 10070 23899 10122 23902
rect 10178 23899 10230 23902
rect 10286 23899 10338 23902
rect 10394 23899 10446 23902
rect 10502 23899 10554 23902
rect 10610 23899 10662 23902
rect 10718 23899 10770 23902
rect 10826 23899 10878 23902
rect 10934 23899 10986 23902
rect 11042 23899 11094 23902
rect 11150 23899 11202 23902
rect 1233 23835 1285 23887
rect 1341 23835 1393 23887
rect 1233 23727 1256 23779
rect 1256 23727 1285 23779
rect 1341 23727 1393 23779
rect 1233 23619 1256 23671
rect 1256 23619 1285 23671
rect 1341 23619 1393 23671
rect 1233 23511 1256 23563
rect 1256 23511 1285 23563
rect 1341 23511 1393 23563
rect 1233 23403 1256 23455
rect 1256 23403 1285 23455
rect 1341 23403 1393 23455
rect 1233 23295 1256 23347
rect 1256 23295 1285 23347
rect 1341 23295 1393 23347
rect 1233 23187 1256 23239
rect 1256 23187 1285 23239
rect 1341 23187 1393 23239
rect 1233 23079 1256 23131
rect 1256 23079 1285 23131
rect 1341 23079 1393 23131
rect 1233 22971 1256 23023
rect 1256 22971 1285 23023
rect 1341 22971 1393 23023
rect 1233 22863 1256 22915
rect 1256 22863 1285 22915
rect 1341 22863 1393 22915
rect 1233 22755 1256 22807
rect 1256 22755 1285 22807
rect 1341 22755 1393 22807
rect 1233 22647 1256 22699
rect 1256 22647 1285 22699
rect 1341 22647 1393 22699
rect 1233 22539 1256 22591
rect 1256 22539 1285 22591
rect 1341 22539 1393 22591
rect 1233 22431 1256 22483
rect 1256 22431 1285 22483
rect 1341 22431 1393 22483
rect 1233 22323 1256 22375
rect 1256 22323 1285 22375
rect 1341 22323 1393 22375
rect 1233 22215 1256 22267
rect 1256 22215 1285 22267
rect 1341 22215 1393 22267
rect 1233 22107 1256 22159
rect 1256 22107 1285 22159
rect 1341 22107 1393 22159
rect 1233 21999 1256 22051
rect 1256 21999 1285 22051
rect 1341 21999 1393 22051
rect 1233 21891 1256 21943
rect 1256 21891 1285 21943
rect 1341 21891 1393 21943
rect 1233 21783 1256 21835
rect 1256 21783 1285 21835
rect 1341 21783 1393 21835
rect 1233 21675 1256 21727
rect 1256 21675 1285 21727
rect 1341 21675 1393 21727
rect 1233 21567 1256 21619
rect 1256 21567 1285 21619
rect 1341 21567 1393 21619
rect 1233 21459 1256 21511
rect 1256 21459 1285 21511
rect 1341 21459 1393 21511
rect 1233 21351 1256 21403
rect 1256 21351 1285 21403
rect 1341 21351 1393 21403
rect 1233 21243 1256 21295
rect 1256 21243 1285 21295
rect 1341 21243 1393 21295
rect 1233 21135 1256 21187
rect 1256 21135 1285 21187
rect 1341 21135 1393 21187
rect 1233 21027 1256 21079
rect 1256 21027 1285 21079
rect 1341 21027 1393 21079
rect 1233 20919 1256 20971
rect 1256 20919 1285 20971
rect 1341 20919 1393 20971
rect 1233 20811 1256 20863
rect 1256 20811 1285 20863
rect 1341 20811 1393 20863
rect 1233 20703 1256 20755
rect 1256 20703 1285 20755
rect 1341 20703 1393 20755
rect 1233 20595 1256 20647
rect 1256 20595 1285 20647
rect 1341 20595 1393 20647
rect 1233 20487 1256 20539
rect 1256 20487 1285 20539
rect 1341 20487 1393 20539
rect 1233 20379 1256 20431
rect 1256 20379 1285 20431
rect 1341 20379 1393 20431
rect 1233 20271 1256 20323
rect 1256 20271 1285 20323
rect 1341 20271 1393 20323
rect 1233 20163 1256 20215
rect 1256 20163 1285 20215
rect 1341 20163 1393 20215
rect 1233 20055 1256 20107
rect 1256 20055 1285 20107
rect 1341 20055 1393 20107
rect 1233 19947 1256 19999
rect 1256 19947 1285 19999
rect 1341 19947 1393 19999
rect 1233 19839 1256 19891
rect 1256 19839 1285 19891
rect 1341 19839 1393 19891
rect 1233 19731 1256 19783
rect 1256 19731 1285 19783
rect 1341 19731 1393 19783
rect 1233 19623 1256 19675
rect 1256 19623 1285 19675
rect 1341 19623 1393 19675
rect 1233 19515 1256 19567
rect 1256 19515 1285 19567
rect 1341 19515 1393 19567
rect 1233 19407 1256 19459
rect 1256 19407 1285 19459
rect 1341 19407 1393 19459
rect 1233 19299 1256 19351
rect 1256 19299 1285 19351
rect 1341 19299 1393 19351
rect 1233 19191 1256 19243
rect 1256 19191 1285 19243
rect 1341 19191 1393 19243
rect 11569 23835 11621 23887
rect 11677 23835 11729 23887
rect 1493 23704 1545 23707
rect 1601 23704 1653 23707
rect 3863 23704 3915 23707
rect 3971 23704 4023 23707
rect 6239 23704 6291 23707
rect 6347 23704 6399 23707
rect 6455 23704 6507 23707
rect 6563 23704 6615 23707
rect 6671 23704 6723 23707
rect 8939 23704 8991 23707
rect 9047 23704 9099 23707
rect 11309 23704 11361 23707
rect 11417 23704 11469 23707
rect 1493 23658 1494 23704
rect 1494 23658 1545 23704
rect 1601 23658 1653 23704
rect 3863 23658 3915 23704
rect 3971 23658 4023 23704
rect 6239 23658 6291 23704
rect 6347 23658 6399 23704
rect 6455 23658 6507 23704
rect 6563 23658 6615 23704
rect 6671 23658 6723 23704
rect 8939 23658 8991 23704
rect 9047 23658 9099 23704
rect 11309 23658 11361 23704
rect 11417 23658 11468 23704
rect 11468 23658 11469 23704
rect 1493 23655 1545 23658
rect 1601 23655 1653 23658
rect 3863 23655 3915 23658
rect 3971 23655 4023 23658
rect 6239 23655 6291 23658
rect 6347 23655 6399 23658
rect 6455 23655 6507 23658
rect 6563 23655 6615 23658
rect 6671 23655 6723 23658
rect 8939 23655 8991 23658
rect 9047 23655 9099 23658
rect 11309 23655 11361 23658
rect 11417 23655 11469 23658
rect 1760 23460 1812 23463
rect 1868 23460 1920 23463
rect 1976 23460 2028 23463
rect 2084 23460 2136 23463
rect 2192 23460 2244 23463
rect 2300 23460 2352 23463
rect 2408 23460 2460 23463
rect 2516 23460 2568 23463
rect 2624 23460 2676 23463
rect 2732 23460 2784 23463
rect 2840 23460 2892 23463
rect 2948 23460 3000 23463
rect 3056 23460 3108 23463
rect 3164 23460 3216 23463
rect 3272 23460 3324 23463
rect 3380 23460 3432 23463
rect 3488 23460 3540 23463
rect 3596 23460 3648 23463
rect 3704 23460 3756 23463
rect 4130 23460 4182 23463
rect 4238 23460 4290 23463
rect 4346 23460 4398 23463
rect 4454 23460 4506 23463
rect 4562 23460 4614 23463
rect 4670 23460 4722 23463
rect 4778 23460 4830 23463
rect 4886 23460 4938 23463
rect 4994 23460 5046 23463
rect 5102 23460 5154 23463
rect 5210 23460 5262 23463
rect 5318 23460 5370 23463
rect 5426 23460 5478 23463
rect 5534 23460 5586 23463
rect 5642 23460 5694 23463
rect 5750 23460 5802 23463
rect 5858 23460 5910 23463
rect 5966 23460 6018 23463
rect 6074 23460 6126 23463
rect 6836 23460 6888 23463
rect 6944 23460 6996 23463
rect 7052 23460 7104 23463
rect 7160 23460 7212 23463
rect 7268 23460 7320 23463
rect 7376 23460 7428 23463
rect 7484 23460 7536 23463
rect 7592 23460 7644 23463
rect 7700 23460 7752 23463
rect 7808 23460 7860 23463
rect 7916 23460 7968 23463
rect 8024 23460 8076 23463
rect 8132 23460 8184 23463
rect 8240 23460 8292 23463
rect 8348 23460 8400 23463
rect 8456 23460 8508 23463
rect 8564 23460 8616 23463
rect 8672 23460 8724 23463
rect 8780 23460 8832 23463
rect 9206 23460 9258 23463
rect 9314 23460 9366 23463
rect 9422 23460 9474 23463
rect 9530 23460 9582 23463
rect 9638 23460 9690 23463
rect 9746 23460 9798 23463
rect 9854 23460 9906 23463
rect 9962 23460 10014 23463
rect 10070 23460 10122 23463
rect 10178 23460 10230 23463
rect 10286 23460 10338 23463
rect 10394 23460 10446 23463
rect 10502 23460 10554 23463
rect 10610 23460 10662 23463
rect 10718 23460 10770 23463
rect 10826 23460 10878 23463
rect 10934 23460 10986 23463
rect 11042 23460 11094 23463
rect 11150 23460 11202 23463
rect 1760 23414 1812 23460
rect 1868 23414 1920 23460
rect 1976 23414 2028 23460
rect 2084 23414 2136 23460
rect 2192 23414 2244 23460
rect 2300 23414 2352 23460
rect 2408 23414 2460 23460
rect 2516 23414 2568 23460
rect 2624 23414 2676 23460
rect 2732 23414 2784 23460
rect 2840 23414 2892 23460
rect 2948 23414 3000 23460
rect 3056 23414 3108 23460
rect 3164 23414 3216 23460
rect 3272 23414 3324 23460
rect 3380 23414 3432 23460
rect 3488 23414 3540 23460
rect 3596 23414 3648 23460
rect 3704 23414 3756 23460
rect 4130 23414 4182 23460
rect 4238 23414 4290 23460
rect 4346 23414 4398 23460
rect 4454 23414 4506 23460
rect 4562 23414 4614 23460
rect 4670 23414 4722 23460
rect 4778 23414 4830 23460
rect 4886 23414 4938 23460
rect 4994 23414 5046 23460
rect 5102 23414 5154 23460
rect 5210 23414 5262 23460
rect 5318 23414 5370 23460
rect 5426 23414 5478 23460
rect 5534 23414 5586 23460
rect 5642 23414 5694 23460
rect 5750 23414 5802 23460
rect 5858 23414 5910 23460
rect 5966 23414 6018 23460
rect 6074 23414 6126 23460
rect 6836 23414 6888 23460
rect 6944 23414 6996 23460
rect 7052 23414 7104 23460
rect 7160 23414 7212 23460
rect 7268 23414 7320 23460
rect 7376 23414 7428 23460
rect 7484 23414 7536 23460
rect 7592 23414 7644 23460
rect 7700 23414 7752 23460
rect 7808 23414 7860 23460
rect 7916 23414 7968 23460
rect 8024 23414 8076 23460
rect 8132 23414 8184 23460
rect 8240 23414 8292 23460
rect 8348 23414 8400 23460
rect 8456 23414 8508 23460
rect 8564 23414 8616 23460
rect 8672 23414 8724 23460
rect 8780 23414 8832 23460
rect 9206 23414 9258 23460
rect 9314 23414 9366 23460
rect 9422 23414 9474 23460
rect 9530 23414 9582 23460
rect 9638 23414 9690 23460
rect 9746 23414 9798 23460
rect 9854 23414 9906 23460
rect 9962 23414 10014 23460
rect 10070 23414 10122 23460
rect 10178 23414 10230 23460
rect 10286 23414 10338 23460
rect 10394 23414 10446 23460
rect 10502 23414 10554 23460
rect 10610 23414 10662 23460
rect 10718 23414 10770 23460
rect 10826 23414 10878 23460
rect 10934 23414 10986 23460
rect 11042 23414 11094 23460
rect 11150 23414 11202 23460
rect 1760 23411 1812 23414
rect 1868 23411 1920 23414
rect 1976 23411 2028 23414
rect 2084 23411 2136 23414
rect 2192 23411 2244 23414
rect 2300 23411 2352 23414
rect 2408 23411 2460 23414
rect 2516 23411 2568 23414
rect 2624 23411 2676 23414
rect 2732 23411 2784 23414
rect 2840 23411 2892 23414
rect 2948 23411 3000 23414
rect 3056 23411 3108 23414
rect 3164 23411 3216 23414
rect 3272 23411 3324 23414
rect 3380 23411 3432 23414
rect 3488 23411 3540 23414
rect 3596 23411 3648 23414
rect 3704 23411 3756 23414
rect 4130 23411 4182 23414
rect 4238 23411 4290 23414
rect 4346 23411 4398 23414
rect 4454 23411 4506 23414
rect 4562 23411 4614 23414
rect 4670 23411 4722 23414
rect 4778 23411 4830 23414
rect 4886 23411 4938 23414
rect 4994 23411 5046 23414
rect 5102 23411 5154 23414
rect 5210 23411 5262 23414
rect 5318 23411 5370 23414
rect 5426 23411 5478 23414
rect 5534 23411 5586 23414
rect 5642 23411 5694 23414
rect 5750 23411 5802 23414
rect 5858 23411 5910 23414
rect 5966 23411 6018 23414
rect 6074 23411 6126 23414
rect 6836 23411 6888 23414
rect 6944 23411 6996 23414
rect 7052 23411 7104 23414
rect 7160 23411 7212 23414
rect 7268 23411 7320 23414
rect 7376 23411 7428 23414
rect 7484 23411 7536 23414
rect 7592 23411 7644 23414
rect 7700 23411 7752 23414
rect 7808 23411 7860 23414
rect 7916 23411 7968 23414
rect 8024 23411 8076 23414
rect 8132 23411 8184 23414
rect 8240 23411 8292 23414
rect 8348 23411 8400 23414
rect 8456 23411 8508 23414
rect 8564 23411 8616 23414
rect 8672 23411 8724 23414
rect 8780 23411 8832 23414
rect 9206 23411 9258 23414
rect 9314 23411 9366 23414
rect 9422 23411 9474 23414
rect 9530 23411 9582 23414
rect 9638 23411 9690 23414
rect 9746 23411 9798 23414
rect 9854 23411 9906 23414
rect 9962 23411 10014 23414
rect 10070 23411 10122 23414
rect 10178 23411 10230 23414
rect 10286 23411 10338 23414
rect 10394 23411 10446 23414
rect 10502 23411 10554 23414
rect 10610 23411 10662 23414
rect 10718 23411 10770 23414
rect 10826 23411 10878 23414
rect 10934 23411 10986 23414
rect 11042 23411 11094 23414
rect 11150 23411 11202 23414
rect 1493 23216 1545 23219
rect 1601 23216 1653 23219
rect 3863 23216 3915 23219
rect 3971 23216 4023 23219
rect 6239 23216 6291 23219
rect 6347 23216 6399 23219
rect 6455 23216 6507 23219
rect 6563 23216 6615 23219
rect 6671 23216 6723 23219
rect 8939 23216 8991 23219
rect 9047 23216 9099 23219
rect 11309 23216 11361 23219
rect 11417 23216 11469 23219
rect 1493 23170 1494 23216
rect 1494 23170 1545 23216
rect 1601 23170 1653 23216
rect 3863 23170 3915 23216
rect 3971 23170 4023 23216
rect 6239 23170 6291 23216
rect 6347 23170 6399 23216
rect 6455 23170 6507 23216
rect 6563 23170 6615 23216
rect 6671 23170 6723 23216
rect 8939 23170 8991 23216
rect 9047 23170 9099 23216
rect 11309 23170 11361 23216
rect 11417 23170 11468 23216
rect 11468 23170 11469 23216
rect 1493 23167 1545 23170
rect 1601 23167 1653 23170
rect 3863 23167 3915 23170
rect 3971 23167 4023 23170
rect 6239 23167 6291 23170
rect 6347 23167 6399 23170
rect 6455 23167 6507 23170
rect 6563 23167 6615 23170
rect 6671 23167 6723 23170
rect 8939 23167 8991 23170
rect 9047 23167 9099 23170
rect 11309 23167 11361 23170
rect 11417 23167 11469 23170
rect 1760 22972 1812 22975
rect 1868 22972 1920 22975
rect 1976 22972 2028 22975
rect 2084 22972 2136 22975
rect 2192 22972 2244 22975
rect 2300 22972 2352 22975
rect 2408 22972 2460 22975
rect 2516 22972 2568 22975
rect 2624 22972 2676 22975
rect 2732 22972 2784 22975
rect 2840 22972 2892 22975
rect 2948 22972 3000 22975
rect 3056 22972 3108 22975
rect 3164 22972 3216 22975
rect 3272 22972 3324 22975
rect 3380 22972 3432 22975
rect 3488 22972 3540 22975
rect 3596 22972 3648 22975
rect 3704 22972 3756 22975
rect 4130 22972 4182 22975
rect 4238 22972 4290 22975
rect 4346 22972 4398 22975
rect 4454 22972 4506 22975
rect 4562 22972 4614 22975
rect 4670 22972 4722 22975
rect 4778 22972 4830 22975
rect 4886 22972 4938 22975
rect 4994 22972 5046 22975
rect 5102 22972 5154 22975
rect 5210 22972 5262 22975
rect 5318 22972 5370 22975
rect 5426 22972 5478 22975
rect 5534 22972 5586 22975
rect 5642 22972 5694 22975
rect 5750 22972 5802 22975
rect 5858 22972 5910 22975
rect 5966 22972 6018 22975
rect 6074 22972 6126 22975
rect 6836 22972 6888 22975
rect 6944 22972 6996 22975
rect 7052 22972 7104 22975
rect 7160 22972 7212 22975
rect 7268 22972 7320 22975
rect 7376 22972 7428 22975
rect 7484 22972 7536 22975
rect 7592 22972 7644 22975
rect 7700 22972 7752 22975
rect 7808 22972 7860 22975
rect 7916 22972 7968 22975
rect 8024 22972 8076 22975
rect 8132 22972 8184 22975
rect 8240 22972 8292 22975
rect 8348 22972 8400 22975
rect 8456 22972 8508 22975
rect 8564 22972 8616 22975
rect 8672 22972 8724 22975
rect 8780 22972 8832 22975
rect 9206 22972 9258 22975
rect 9314 22972 9366 22975
rect 9422 22972 9474 22975
rect 9530 22972 9582 22975
rect 9638 22972 9690 22975
rect 9746 22972 9798 22975
rect 9854 22972 9906 22975
rect 9962 22972 10014 22975
rect 10070 22972 10122 22975
rect 10178 22972 10230 22975
rect 10286 22972 10338 22975
rect 10394 22972 10446 22975
rect 10502 22972 10554 22975
rect 10610 22972 10662 22975
rect 10718 22972 10770 22975
rect 10826 22972 10878 22975
rect 10934 22972 10986 22975
rect 11042 22972 11094 22975
rect 11150 22972 11202 22975
rect 1760 22926 1812 22972
rect 1868 22926 1920 22972
rect 1976 22926 2028 22972
rect 2084 22926 2136 22972
rect 2192 22926 2244 22972
rect 2300 22926 2352 22972
rect 2408 22926 2460 22972
rect 2516 22926 2568 22972
rect 2624 22926 2676 22972
rect 2732 22926 2784 22972
rect 2840 22926 2892 22972
rect 2948 22926 3000 22972
rect 3056 22926 3108 22972
rect 3164 22926 3216 22972
rect 3272 22926 3324 22972
rect 3380 22926 3432 22972
rect 3488 22926 3540 22972
rect 3596 22926 3648 22972
rect 3704 22926 3756 22972
rect 4130 22926 4182 22972
rect 4238 22926 4290 22972
rect 4346 22926 4398 22972
rect 4454 22926 4506 22972
rect 4562 22926 4614 22972
rect 4670 22926 4722 22972
rect 4778 22926 4830 22972
rect 4886 22926 4938 22972
rect 4994 22926 5046 22972
rect 5102 22926 5154 22972
rect 5210 22926 5262 22972
rect 5318 22926 5370 22972
rect 5426 22926 5478 22972
rect 5534 22926 5586 22972
rect 5642 22926 5694 22972
rect 5750 22926 5802 22972
rect 5858 22926 5910 22972
rect 5966 22926 6018 22972
rect 6074 22926 6126 22972
rect 6836 22926 6888 22972
rect 6944 22926 6996 22972
rect 7052 22926 7104 22972
rect 7160 22926 7212 22972
rect 7268 22926 7320 22972
rect 7376 22926 7428 22972
rect 7484 22926 7536 22972
rect 7592 22926 7644 22972
rect 7700 22926 7752 22972
rect 7808 22926 7860 22972
rect 7916 22926 7968 22972
rect 8024 22926 8076 22972
rect 8132 22926 8184 22972
rect 8240 22926 8292 22972
rect 8348 22926 8400 22972
rect 8456 22926 8508 22972
rect 8564 22926 8616 22972
rect 8672 22926 8724 22972
rect 8780 22926 8832 22972
rect 9206 22926 9258 22972
rect 9314 22926 9366 22972
rect 9422 22926 9474 22972
rect 9530 22926 9582 22972
rect 9638 22926 9690 22972
rect 9746 22926 9798 22972
rect 9854 22926 9906 22972
rect 9962 22926 10014 22972
rect 10070 22926 10122 22972
rect 10178 22926 10230 22972
rect 10286 22926 10338 22972
rect 10394 22926 10446 22972
rect 10502 22926 10554 22972
rect 10610 22926 10662 22972
rect 10718 22926 10770 22972
rect 10826 22926 10878 22972
rect 10934 22926 10986 22972
rect 11042 22926 11094 22972
rect 11150 22926 11202 22972
rect 1760 22923 1812 22926
rect 1868 22923 1920 22926
rect 1976 22923 2028 22926
rect 2084 22923 2136 22926
rect 2192 22923 2244 22926
rect 2300 22923 2352 22926
rect 2408 22923 2460 22926
rect 2516 22923 2568 22926
rect 2624 22923 2676 22926
rect 2732 22923 2784 22926
rect 2840 22923 2892 22926
rect 2948 22923 3000 22926
rect 3056 22923 3108 22926
rect 3164 22923 3216 22926
rect 3272 22923 3324 22926
rect 3380 22923 3432 22926
rect 3488 22923 3540 22926
rect 3596 22923 3648 22926
rect 3704 22923 3756 22926
rect 4130 22923 4182 22926
rect 4238 22923 4290 22926
rect 4346 22923 4398 22926
rect 4454 22923 4506 22926
rect 4562 22923 4614 22926
rect 4670 22923 4722 22926
rect 4778 22923 4830 22926
rect 4886 22923 4938 22926
rect 4994 22923 5046 22926
rect 5102 22923 5154 22926
rect 5210 22923 5262 22926
rect 5318 22923 5370 22926
rect 5426 22923 5478 22926
rect 5534 22923 5586 22926
rect 5642 22923 5694 22926
rect 5750 22923 5802 22926
rect 5858 22923 5910 22926
rect 5966 22923 6018 22926
rect 6074 22923 6126 22926
rect 6836 22923 6888 22926
rect 6944 22923 6996 22926
rect 7052 22923 7104 22926
rect 7160 22923 7212 22926
rect 7268 22923 7320 22926
rect 7376 22923 7428 22926
rect 7484 22923 7536 22926
rect 7592 22923 7644 22926
rect 7700 22923 7752 22926
rect 7808 22923 7860 22926
rect 7916 22923 7968 22926
rect 8024 22923 8076 22926
rect 8132 22923 8184 22926
rect 8240 22923 8292 22926
rect 8348 22923 8400 22926
rect 8456 22923 8508 22926
rect 8564 22923 8616 22926
rect 8672 22923 8724 22926
rect 8780 22923 8832 22926
rect 9206 22923 9258 22926
rect 9314 22923 9366 22926
rect 9422 22923 9474 22926
rect 9530 22923 9582 22926
rect 9638 22923 9690 22926
rect 9746 22923 9798 22926
rect 9854 22923 9906 22926
rect 9962 22923 10014 22926
rect 10070 22923 10122 22926
rect 10178 22923 10230 22926
rect 10286 22923 10338 22926
rect 10394 22923 10446 22926
rect 10502 22923 10554 22926
rect 10610 22923 10662 22926
rect 10718 22923 10770 22926
rect 10826 22923 10878 22926
rect 10934 22923 10986 22926
rect 11042 22923 11094 22926
rect 11150 22923 11202 22926
rect 1493 22728 1545 22731
rect 1601 22728 1653 22731
rect 3863 22728 3915 22731
rect 3971 22728 4023 22731
rect 6239 22728 6291 22731
rect 6347 22728 6399 22731
rect 6455 22728 6507 22731
rect 6563 22728 6615 22731
rect 6671 22728 6723 22731
rect 8939 22728 8991 22731
rect 9047 22728 9099 22731
rect 11309 22728 11361 22731
rect 11417 22728 11469 22731
rect 1493 22682 1494 22728
rect 1494 22682 1545 22728
rect 1601 22682 1653 22728
rect 3863 22682 3915 22728
rect 3971 22682 4023 22728
rect 6239 22682 6291 22728
rect 6347 22682 6399 22728
rect 6455 22682 6507 22728
rect 6563 22682 6615 22728
rect 6671 22682 6723 22728
rect 8939 22682 8991 22728
rect 9047 22682 9099 22728
rect 11309 22682 11361 22728
rect 11417 22682 11468 22728
rect 11468 22682 11469 22728
rect 1493 22679 1545 22682
rect 1601 22679 1653 22682
rect 3863 22679 3915 22682
rect 3971 22679 4023 22682
rect 6239 22679 6291 22682
rect 6347 22679 6399 22682
rect 6455 22679 6507 22682
rect 6563 22679 6615 22682
rect 6671 22679 6723 22682
rect 8939 22679 8991 22682
rect 9047 22679 9099 22682
rect 11309 22679 11361 22682
rect 11417 22679 11469 22682
rect 1760 22484 1812 22487
rect 1868 22484 1920 22487
rect 1976 22484 2028 22487
rect 2084 22484 2136 22487
rect 2192 22484 2244 22487
rect 2300 22484 2352 22487
rect 2408 22484 2460 22487
rect 2516 22484 2568 22487
rect 2624 22484 2676 22487
rect 2732 22484 2784 22487
rect 2840 22484 2892 22487
rect 2948 22484 3000 22487
rect 3056 22484 3108 22487
rect 3164 22484 3216 22487
rect 3272 22484 3324 22487
rect 3380 22484 3432 22487
rect 3488 22484 3540 22487
rect 3596 22484 3648 22487
rect 3704 22484 3756 22487
rect 4130 22484 4182 22487
rect 4238 22484 4290 22487
rect 4346 22484 4398 22487
rect 4454 22484 4506 22487
rect 4562 22484 4614 22487
rect 4670 22484 4722 22487
rect 4778 22484 4830 22487
rect 4886 22484 4938 22487
rect 4994 22484 5046 22487
rect 5102 22484 5154 22487
rect 5210 22484 5262 22487
rect 5318 22484 5370 22487
rect 5426 22484 5478 22487
rect 5534 22484 5586 22487
rect 5642 22484 5694 22487
rect 5750 22484 5802 22487
rect 5858 22484 5910 22487
rect 5966 22484 6018 22487
rect 6074 22484 6126 22487
rect 6836 22484 6888 22487
rect 6944 22484 6996 22487
rect 7052 22484 7104 22487
rect 7160 22484 7212 22487
rect 7268 22484 7320 22487
rect 7376 22484 7428 22487
rect 7484 22484 7536 22487
rect 7592 22484 7644 22487
rect 7700 22484 7752 22487
rect 7808 22484 7860 22487
rect 7916 22484 7968 22487
rect 8024 22484 8076 22487
rect 8132 22484 8184 22487
rect 8240 22484 8292 22487
rect 8348 22484 8400 22487
rect 8456 22484 8508 22487
rect 8564 22484 8616 22487
rect 8672 22484 8724 22487
rect 8780 22484 8832 22487
rect 9206 22484 9258 22487
rect 9314 22484 9366 22487
rect 9422 22484 9474 22487
rect 9530 22484 9582 22487
rect 9638 22484 9690 22487
rect 9746 22484 9798 22487
rect 9854 22484 9906 22487
rect 9962 22484 10014 22487
rect 10070 22484 10122 22487
rect 10178 22484 10230 22487
rect 10286 22484 10338 22487
rect 10394 22484 10446 22487
rect 10502 22484 10554 22487
rect 10610 22484 10662 22487
rect 10718 22484 10770 22487
rect 10826 22484 10878 22487
rect 10934 22484 10986 22487
rect 11042 22484 11094 22487
rect 11150 22484 11202 22487
rect 1760 22438 1812 22484
rect 1868 22438 1920 22484
rect 1976 22438 2028 22484
rect 2084 22438 2136 22484
rect 2192 22438 2244 22484
rect 2300 22438 2352 22484
rect 2408 22438 2460 22484
rect 2516 22438 2568 22484
rect 2624 22438 2676 22484
rect 2732 22438 2784 22484
rect 2840 22438 2892 22484
rect 2948 22438 3000 22484
rect 3056 22438 3108 22484
rect 3164 22438 3216 22484
rect 3272 22438 3324 22484
rect 3380 22438 3432 22484
rect 3488 22438 3540 22484
rect 3596 22438 3648 22484
rect 3704 22438 3756 22484
rect 4130 22438 4182 22484
rect 4238 22438 4290 22484
rect 4346 22438 4398 22484
rect 4454 22438 4506 22484
rect 4562 22438 4614 22484
rect 4670 22438 4722 22484
rect 4778 22438 4830 22484
rect 4886 22438 4938 22484
rect 4994 22438 5046 22484
rect 5102 22438 5154 22484
rect 5210 22438 5262 22484
rect 5318 22438 5370 22484
rect 5426 22438 5478 22484
rect 5534 22438 5586 22484
rect 5642 22438 5694 22484
rect 5750 22438 5802 22484
rect 5858 22438 5910 22484
rect 5966 22438 6018 22484
rect 6074 22438 6126 22484
rect 6836 22438 6888 22484
rect 6944 22438 6996 22484
rect 7052 22438 7104 22484
rect 7160 22438 7212 22484
rect 7268 22438 7320 22484
rect 7376 22438 7428 22484
rect 7484 22438 7536 22484
rect 7592 22438 7644 22484
rect 7700 22438 7752 22484
rect 7808 22438 7860 22484
rect 7916 22438 7968 22484
rect 8024 22438 8076 22484
rect 8132 22438 8184 22484
rect 8240 22438 8292 22484
rect 8348 22438 8400 22484
rect 8456 22438 8508 22484
rect 8564 22438 8616 22484
rect 8672 22438 8724 22484
rect 8780 22438 8832 22484
rect 9206 22438 9258 22484
rect 9314 22438 9366 22484
rect 9422 22438 9474 22484
rect 9530 22438 9582 22484
rect 9638 22438 9690 22484
rect 9746 22438 9798 22484
rect 9854 22438 9906 22484
rect 9962 22438 10014 22484
rect 10070 22438 10122 22484
rect 10178 22438 10230 22484
rect 10286 22438 10338 22484
rect 10394 22438 10446 22484
rect 10502 22438 10554 22484
rect 10610 22438 10662 22484
rect 10718 22438 10770 22484
rect 10826 22438 10878 22484
rect 10934 22438 10986 22484
rect 11042 22438 11094 22484
rect 11150 22438 11202 22484
rect 1760 22435 1812 22438
rect 1868 22435 1920 22438
rect 1976 22435 2028 22438
rect 2084 22435 2136 22438
rect 2192 22435 2244 22438
rect 2300 22435 2352 22438
rect 2408 22435 2460 22438
rect 2516 22435 2568 22438
rect 2624 22435 2676 22438
rect 2732 22435 2784 22438
rect 2840 22435 2892 22438
rect 2948 22435 3000 22438
rect 3056 22435 3108 22438
rect 3164 22435 3216 22438
rect 3272 22435 3324 22438
rect 3380 22435 3432 22438
rect 3488 22435 3540 22438
rect 3596 22435 3648 22438
rect 3704 22435 3756 22438
rect 4130 22435 4182 22438
rect 4238 22435 4290 22438
rect 4346 22435 4398 22438
rect 4454 22435 4506 22438
rect 4562 22435 4614 22438
rect 4670 22435 4722 22438
rect 4778 22435 4830 22438
rect 4886 22435 4938 22438
rect 4994 22435 5046 22438
rect 5102 22435 5154 22438
rect 5210 22435 5262 22438
rect 5318 22435 5370 22438
rect 5426 22435 5478 22438
rect 5534 22435 5586 22438
rect 5642 22435 5694 22438
rect 5750 22435 5802 22438
rect 5858 22435 5910 22438
rect 5966 22435 6018 22438
rect 6074 22435 6126 22438
rect 6836 22435 6888 22438
rect 6944 22435 6996 22438
rect 7052 22435 7104 22438
rect 7160 22435 7212 22438
rect 7268 22435 7320 22438
rect 7376 22435 7428 22438
rect 7484 22435 7536 22438
rect 7592 22435 7644 22438
rect 7700 22435 7752 22438
rect 7808 22435 7860 22438
rect 7916 22435 7968 22438
rect 8024 22435 8076 22438
rect 8132 22435 8184 22438
rect 8240 22435 8292 22438
rect 8348 22435 8400 22438
rect 8456 22435 8508 22438
rect 8564 22435 8616 22438
rect 8672 22435 8724 22438
rect 8780 22435 8832 22438
rect 9206 22435 9258 22438
rect 9314 22435 9366 22438
rect 9422 22435 9474 22438
rect 9530 22435 9582 22438
rect 9638 22435 9690 22438
rect 9746 22435 9798 22438
rect 9854 22435 9906 22438
rect 9962 22435 10014 22438
rect 10070 22435 10122 22438
rect 10178 22435 10230 22438
rect 10286 22435 10338 22438
rect 10394 22435 10446 22438
rect 10502 22435 10554 22438
rect 10610 22435 10662 22438
rect 10718 22435 10770 22438
rect 10826 22435 10878 22438
rect 10934 22435 10986 22438
rect 11042 22435 11094 22438
rect 11150 22435 11202 22438
rect 1493 22240 1545 22243
rect 1601 22240 1653 22243
rect 3863 22240 3915 22243
rect 3971 22240 4023 22243
rect 6239 22240 6291 22243
rect 6347 22240 6399 22243
rect 6455 22240 6507 22243
rect 6563 22240 6615 22243
rect 6671 22240 6723 22243
rect 8939 22240 8991 22243
rect 9047 22240 9099 22243
rect 11309 22240 11361 22243
rect 11417 22240 11469 22243
rect 1493 22194 1494 22240
rect 1494 22194 1545 22240
rect 1601 22194 1653 22240
rect 3863 22194 3915 22240
rect 3971 22194 4023 22240
rect 6239 22194 6291 22240
rect 6347 22194 6399 22240
rect 6455 22194 6507 22240
rect 6563 22194 6615 22240
rect 6671 22194 6723 22240
rect 8939 22194 8991 22240
rect 9047 22194 9099 22240
rect 11309 22194 11361 22240
rect 11417 22194 11468 22240
rect 11468 22194 11469 22240
rect 1493 22191 1545 22194
rect 1601 22191 1653 22194
rect 3863 22191 3915 22194
rect 3971 22191 4023 22194
rect 6239 22191 6291 22194
rect 6347 22191 6399 22194
rect 6455 22191 6507 22194
rect 6563 22191 6615 22194
rect 6671 22191 6723 22194
rect 8939 22191 8991 22194
rect 9047 22191 9099 22194
rect 11309 22191 11361 22194
rect 11417 22191 11469 22194
rect 1760 21996 1812 21999
rect 1868 21996 1920 21999
rect 1976 21996 2028 21999
rect 2084 21996 2136 21999
rect 2192 21996 2244 21999
rect 2300 21996 2352 21999
rect 2408 21996 2460 21999
rect 2516 21996 2568 21999
rect 2624 21996 2676 21999
rect 2732 21996 2784 21999
rect 2840 21996 2892 21999
rect 2948 21996 3000 21999
rect 3056 21996 3108 21999
rect 3164 21996 3216 21999
rect 3272 21996 3324 21999
rect 3380 21996 3432 21999
rect 3488 21996 3540 21999
rect 3596 21996 3648 21999
rect 3704 21996 3756 21999
rect 4130 21996 4182 21999
rect 4238 21996 4290 21999
rect 4346 21996 4398 21999
rect 4454 21996 4506 21999
rect 4562 21996 4614 21999
rect 4670 21996 4722 21999
rect 4778 21996 4830 21999
rect 4886 21996 4938 21999
rect 4994 21996 5046 21999
rect 5102 21996 5154 21999
rect 5210 21996 5262 21999
rect 5318 21996 5370 21999
rect 5426 21996 5478 21999
rect 5534 21996 5586 21999
rect 5642 21996 5694 21999
rect 5750 21996 5802 21999
rect 5858 21996 5910 21999
rect 5966 21996 6018 21999
rect 6074 21996 6126 21999
rect 6836 21996 6888 21999
rect 6944 21996 6996 21999
rect 7052 21996 7104 21999
rect 7160 21996 7212 21999
rect 7268 21996 7320 21999
rect 7376 21996 7428 21999
rect 7484 21996 7536 21999
rect 7592 21996 7644 21999
rect 7700 21996 7752 21999
rect 7808 21996 7860 21999
rect 7916 21996 7968 21999
rect 8024 21996 8076 21999
rect 8132 21996 8184 21999
rect 8240 21996 8292 21999
rect 8348 21996 8400 21999
rect 8456 21996 8508 21999
rect 8564 21996 8616 21999
rect 8672 21996 8724 21999
rect 8780 21996 8832 21999
rect 9206 21996 9258 21999
rect 9314 21996 9366 21999
rect 9422 21996 9474 21999
rect 9530 21996 9582 21999
rect 9638 21996 9690 21999
rect 9746 21996 9798 21999
rect 9854 21996 9906 21999
rect 9962 21996 10014 21999
rect 10070 21996 10122 21999
rect 10178 21996 10230 21999
rect 10286 21996 10338 21999
rect 10394 21996 10446 21999
rect 10502 21996 10554 21999
rect 10610 21996 10662 21999
rect 10718 21996 10770 21999
rect 10826 21996 10878 21999
rect 10934 21996 10986 21999
rect 11042 21996 11094 21999
rect 11150 21996 11202 21999
rect 1760 21950 1812 21996
rect 1868 21950 1920 21996
rect 1976 21950 2028 21996
rect 2084 21950 2136 21996
rect 2192 21950 2244 21996
rect 2300 21950 2352 21996
rect 2408 21950 2460 21996
rect 2516 21950 2568 21996
rect 2624 21950 2676 21996
rect 2732 21950 2784 21996
rect 2840 21950 2892 21996
rect 2948 21950 3000 21996
rect 3056 21950 3108 21996
rect 3164 21950 3216 21996
rect 3272 21950 3324 21996
rect 3380 21950 3432 21996
rect 3488 21950 3540 21996
rect 3596 21950 3648 21996
rect 3704 21950 3756 21996
rect 4130 21950 4182 21996
rect 4238 21950 4290 21996
rect 4346 21950 4398 21996
rect 4454 21950 4506 21996
rect 4562 21950 4614 21996
rect 4670 21950 4722 21996
rect 4778 21950 4830 21996
rect 4886 21950 4938 21996
rect 4994 21950 5046 21996
rect 5102 21950 5154 21996
rect 5210 21950 5262 21996
rect 5318 21950 5370 21996
rect 5426 21950 5478 21996
rect 5534 21950 5586 21996
rect 5642 21950 5694 21996
rect 5750 21950 5802 21996
rect 5858 21950 5910 21996
rect 5966 21950 6018 21996
rect 6074 21950 6126 21996
rect 6836 21950 6888 21996
rect 6944 21950 6996 21996
rect 7052 21950 7104 21996
rect 7160 21950 7212 21996
rect 7268 21950 7320 21996
rect 7376 21950 7428 21996
rect 7484 21950 7536 21996
rect 7592 21950 7644 21996
rect 7700 21950 7752 21996
rect 7808 21950 7860 21996
rect 7916 21950 7968 21996
rect 8024 21950 8076 21996
rect 8132 21950 8184 21996
rect 8240 21950 8292 21996
rect 8348 21950 8400 21996
rect 8456 21950 8508 21996
rect 8564 21950 8616 21996
rect 8672 21950 8724 21996
rect 8780 21950 8832 21996
rect 9206 21950 9258 21996
rect 9314 21950 9366 21996
rect 9422 21950 9474 21996
rect 9530 21950 9582 21996
rect 9638 21950 9690 21996
rect 9746 21950 9798 21996
rect 9854 21950 9906 21996
rect 9962 21950 10014 21996
rect 10070 21950 10122 21996
rect 10178 21950 10230 21996
rect 10286 21950 10338 21996
rect 10394 21950 10446 21996
rect 10502 21950 10554 21996
rect 10610 21950 10662 21996
rect 10718 21950 10770 21996
rect 10826 21950 10878 21996
rect 10934 21950 10986 21996
rect 11042 21950 11094 21996
rect 11150 21950 11202 21996
rect 1760 21947 1812 21950
rect 1868 21947 1920 21950
rect 1976 21947 2028 21950
rect 2084 21947 2136 21950
rect 2192 21947 2244 21950
rect 2300 21947 2352 21950
rect 2408 21947 2460 21950
rect 2516 21947 2568 21950
rect 2624 21947 2676 21950
rect 2732 21947 2784 21950
rect 2840 21947 2892 21950
rect 2948 21947 3000 21950
rect 3056 21947 3108 21950
rect 3164 21947 3216 21950
rect 3272 21947 3324 21950
rect 3380 21947 3432 21950
rect 3488 21947 3540 21950
rect 3596 21947 3648 21950
rect 3704 21947 3756 21950
rect 4130 21947 4182 21950
rect 4238 21947 4290 21950
rect 4346 21947 4398 21950
rect 4454 21947 4506 21950
rect 4562 21947 4614 21950
rect 4670 21947 4722 21950
rect 4778 21947 4830 21950
rect 4886 21947 4938 21950
rect 4994 21947 5046 21950
rect 5102 21947 5154 21950
rect 5210 21947 5262 21950
rect 5318 21947 5370 21950
rect 5426 21947 5478 21950
rect 5534 21947 5586 21950
rect 5642 21947 5694 21950
rect 5750 21947 5802 21950
rect 5858 21947 5910 21950
rect 5966 21947 6018 21950
rect 6074 21947 6126 21950
rect 6836 21947 6888 21950
rect 6944 21947 6996 21950
rect 7052 21947 7104 21950
rect 7160 21947 7212 21950
rect 7268 21947 7320 21950
rect 7376 21947 7428 21950
rect 7484 21947 7536 21950
rect 7592 21947 7644 21950
rect 7700 21947 7752 21950
rect 7808 21947 7860 21950
rect 7916 21947 7968 21950
rect 8024 21947 8076 21950
rect 8132 21947 8184 21950
rect 8240 21947 8292 21950
rect 8348 21947 8400 21950
rect 8456 21947 8508 21950
rect 8564 21947 8616 21950
rect 8672 21947 8724 21950
rect 8780 21947 8832 21950
rect 9206 21947 9258 21950
rect 9314 21947 9366 21950
rect 9422 21947 9474 21950
rect 9530 21947 9582 21950
rect 9638 21947 9690 21950
rect 9746 21947 9798 21950
rect 9854 21947 9906 21950
rect 9962 21947 10014 21950
rect 10070 21947 10122 21950
rect 10178 21947 10230 21950
rect 10286 21947 10338 21950
rect 10394 21947 10446 21950
rect 10502 21947 10554 21950
rect 10610 21947 10662 21950
rect 10718 21947 10770 21950
rect 10826 21947 10878 21950
rect 10934 21947 10986 21950
rect 11042 21947 11094 21950
rect 11150 21947 11202 21950
rect 1493 21752 1545 21755
rect 1601 21752 1653 21755
rect 3863 21752 3915 21755
rect 3971 21752 4023 21755
rect 6239 21752 6291 21755
rect 6347 21752 6399 21755
rect 6455 21752 6507 21755
rect 6563 21752 6615 21755
rect 6671 21752 6723 21755
rect 8939 21752 8991 21755
rect 9047 21752 9099 21755
rect 11309 21752 11361 21755
rect 11417 21752 11469 21755
rect 1493 21706 1494 21752
rect 1494 21706 1545 21752
rect 1601 21706 1653 21752
rect 3863 21706 3915 21752
rect 3971 21706 4023 21752
rect 6239 21706 6291 21752
rect 6347 21706 6399 21752
rect 6455 21706 6507 21752
rect 6563 21706 6615 21752
rect 6671 21706 6723 21752
rect 8939 21706 8991 21752
rect 9047 21706 9099 21752
rect 11309 21706 11361 21752
rect 11417 21706 11468 21752
rect 11468 21706 11469 21752
rect 1493 21703 1545 21706
rect 1601 21703 1653 21706
rect 3863 21703 3915 21706
rect 3971 21703 4023 21706
rect 6239 21703 6291 21706
rect 6347 21703 6399 21706
rect 6455 21703 6507 21706
rect 6563 21703 6615 21706
rect 6671 21703 6723 21706
rect 8939 21703 8991 21706
rect 9047 21703 9099 21706
rect 11309 21703 11361 21706
rect 11417 21703 11469 21706
rect 1760 21508 1812 21511
rect 1868 21508 1920 21511
rect 1976 21508 2028 21511
rect 2084 21508 2136 21511
rect 2192 21508 2244 21511
rect 2300 21508 2352 21511
rect 2408 21508 2460 21511
rect 2516 21508 2568 21511
rect 2624 21508 2676 21511
rect 2732 21508 2784 21511
rect 2840 21508 2892 21511
rect 2948 21508 3000 21511
rect 3056 21508 3108 21511
rect 3164 21508 3216 21511
rect 3272 21508 3324 21511
rect 3380 21508 3432 21511
rect 3488 21508 3540 21511
rect 3596 21508 3648 21511
rect 3704 21508 3756 21511
rect 4130 21508 4182 21511
rect 4238 21508 4290 21511
rect 4346 21508 4398 21511
rect 4454 21508 4506 21511
rect 4562 21508 4614 21511
rect 4670 21508 4722 21511
rect 4778 21508 4830 21511
rect 4886 21508 4938 21511
rect 4994 21508 5046 21511
rect 5102 21508 5154 21511
rect 5210 21508 5262 21511
rect 5318 21508 5370 21511
rect 5426 21508 5478 21511
rect 5534 21508 5586 21511
rect 5642 21508 5694 21511
rect 5750 21508 5802 21511
rect 5858 21508 5910 21511
rect 5966 21508 6018 21511
rect 6074 21508 6126 21511
rect 6836 21508 6888 21511
rect 6944 21508 6996 21511
rect 7052 21508 7104 21511
rect 7160 21508 7212 21511
rect 7268 21508 7320 21511
rect 7376 21508 7428 21511
rect 7484 21508 7536 21511
rect 7592 21508 7644 21511
rect 7700 21508 7752 21511
rect 7808 21508 7860 21511
rect 7916 21508 7968 21511
rect 8024 21508 8076 21511
rect 8132 21508 8184 21511
rect 8240 21508 8292 21511
rect 8348 21508 8400 21511
rect 8456 21508 8508 21511
rect 8564 21508 8616 21511
rect 8672 21508 8724 21511
rect 8780 21508 8832 21511
rect 9206 21508 9258 21511
rect 9314 21508 9366 21511
rect 9422 21508 9474 21511
rect 9530 21508 9582 21511
rect 9638 21508 9690 21511
rect 9746 21508 9798 21511
rect 9854 21508 9906 21511
rect 9962 21508 10014 21511
rect 10070 21508 10122 21511
rect 10178 21508 10230 21511
rect 10286 21508 10338 21511
rect 10394 21508 10446 21511
rect 10502 21508 10554 21511
rect 10610 21508 10662 21511
rect 10718 21508 10770 21511
rect 10826 21508 10878 21511
rect 10934 21508 10986 21511
rect 11042 21508 11094 21511
rect 11150 21508 11202 21511
rect 1760 21462 1812 21508
rect 1868 21462 1920 21508
rect 1976 21462 2028 21508
rect 2084 21462 2136 21508
rect 2192 21462 2244 21508
rect 2300 21462 2352 21508
rect 2408 21462 2460 21508
rect 2516 21462 2568 21508
rect 2624 21462 2676 21508
rect 2732 21462 2784 21508
rect 2840 21462 2892 21508
rect 2948 21462 3000 21508
rect 3056 21462 3108 21508
rect 3164 21462 3216 21508
rect 3272 21462 3324 21508
rect 3380 21462 3432 21508
rect 3488 21462 3540 21508
rect 3596 21462 3648 21508
rect 3704 21462 3756 21508
rect 4130 21462 4182 21508
rect 4238 21462 4290 21508
rect 4346 21462 4398 21508
rect 4454 21462 4506 21508
rect 4562 21462 4614 21508
rect 4670 21462 4722 21508
rect 4778 21462 4830 21508
rect 4886 21462 4938 21508
rect 4994 21462 5046 21508
rect 5102 21462 5154 21508
rect 5210 21462 5262 21508
rect 5318 21462 5370 21508
rect 5426 21462 5478 21508
rect 5534 21462 5586 21508
rect 5642 21462 5694 21508
rect 5750 21462 5802 21508
rect 5858 21462 5910 21508
rect 5966 21462 6018 21508
rect 6074 21462 6126 21508
rect 6836 21462 6888 21508
rect 6944 21462 6996 21508
rect 7052 21462 7104 21508
rect 7160 21462 7212 21508
rect 7268 21462 7320 21508
rect 7376 21462 7428 21508
rect 7484 21462 7536 21508
rect 7592 21462 7644 21508
rect 7700 21462 7752 21508
rect 7808 21462 7860 21508
rect 7916 21462 7968 21508
rect 8024 21462 8076 21508
rect 8132 21462 8184 21508
rect 8240 21462 8292 21508
rect 8348 21462 8400 21508
rect 8456 21462 8508 21508
rect 8564 21462 8616 21508
rect 8672 21462 8724 21508
rect 8780 21462 8832 21508
rect 9206 21462 9258 21508
rect 9314 21462 9366 21508
rect 9422 21462 9474 21508
rect 9530 21462 9582 21508
rect 9638 21462 9690 21508
rect 9746 21462 9798 21508
rect 9854 21462 9906 21508
rect 9962 21462 10014 21508
rect 10070 21462 10122 21508
rect 10178 21462 10230 21508
rect 10286 21462 10338 21508
rect 10394 21462 10446 21508
rect 10502 21462 10554 21508
rect 10610 21462 10662 21508
rect 10718 21462 10770 21508
rect 10826 21462 10878 21508
rect 10934 21462 10986 21508
rect 11042 21462 11094 21508
rect 11150 21462 11202 21508
rect 1760 21459 1812 21462
rect 1868 21459 1920 21462
rect 1976 21459 2028 21462
rect 2084 21459 2136 21462
rect 2192 21459 2244 21462
rect 2300 21459 2352 21462
rect 2408 21459 2460 21462
rect 2516 21459 2568 21462
rect 2624 21459 2676 21462
rect 2732 21459 2784 21462
rect 2840 21459 2892 21462
rect 2948 21459 3000 21462
rect 3056 21459 3108 21462
rect 3164 21459 3216 21462
rect 3272 21459 3324 21462
rect 3380 21459 3432 21462
rect 3488 21459 3540 21462
rect 3596 21459 3648 21462
rect 3704 21459 3756 21462
rect 4130 21459 4182 21462
rect 4238 21459 4290 21462
rect 4346 21459 4398 21462
rect 4454 21459 4506 21462
rect 4562 21459 4614 21462
rect 4670 21459 4722 21462
rect 4778 21459 4830 21462
rect 4886 21459 4938 21462
rect 4994 21459 5046 21462
rect 5102 21459 5154 21462
rect 5210 21459 5262 21462
rect 5318 21459 5370 21462
rect 5426 21459 5478 21462
rect 5534 21459 5586 21462
rect 5642 21459 5694 21462
rect 5750 21459 5802 21462
rect 5858 21459 5910 21462
rect 5966 21459 6018 21462
rect 6074 21459 6126 21462
rect 6836 21459 6888 21462
rect 6944 21459 6996 21462
rect 7052 21459 7104 21462
rect 7160 21459 7212 21462
rect 7268 21459 7320 21462
rect 7376 21459 7428 21462
rect 7484 21459 7536 21462
rect 7592 21459 7644 21462
rect 7700 21459 7752 21462
rect 7808 21459 7860 21462
rect 7916 21459 7968 21462
rect 8024 21459 8076 21462
rect 8132 21459 8184 21462
rect 8240 21459 8292 21462
rect 8348 21459 8400 21462
rect 8456 21459 8508 21462
rect 8564 21459 8616 21462
rect 8672 21459 8724 21462
rect 8780 21459 8832 21462
rect 9206 21459 9258 21462
rect 9314 21459 9366 21462
rect 9422 21459 9474 21462
rect 9530 21459 9582 21462
rect 9638 21459 9690 21462
rect 9746 21459 9798 21462
rect 9854 21459 9906 21462
rect 9962 21459 10014 21462
rect 10070 21459 10122 21462
rect 10178 21459 10230 21462
rect 10286 21459 10338 21462
rect 10394 21459 10446 21462
rect 10502 21459 10554 21462
rect 10610 21459 10662 21462
rect 10718 21459 10770 21462
rect 10826 21459 10878 21462
rect 10934 21459 10986 21462
rect 11042 21459 11094 21462
rect 11150 21459 11202 21462
rect 1493 21264 1545 21267
rect 1601 21264 1653 21267
rect 3863 21264 3915 21267
rect 3971 21264 4023 21267
rect 6239 21264 6291 21267
rect 6347 21264 6399 21267
rect 6455 21264 6507 21267
rect 6563 21264 6615 21267
rect 6671 21264 6723 21267
rect 8939 21264 8991 21267
rect 9047 21264 9099 21267
rect 11309 21264 11361 21267
rect 11417 21264 11469 21267
rect 1493 21218 1494 21264
rect 1494 21218 1545 21264
rect 1601 21218 1653 21264
rect 3863 21218 3915 21264
rect 3971 21218 4023 21264
rect 6239 21218 6291 21264
rect 6347 21218 6399 21264
rect 6455 21218 6507 21264
rect 6563 21218 6615 21264
rect 6671 21218 6723 21264
rect 8939 21218 8991 21264
rect 9047 21218 9099 21264
rect 11309 21218 11361 21264
rect 11417 21218 11468 21264
rect 11468 21218 11469 21264
rect 1493 21215 1545 21218
rect 1601 21215 1653 21218
rect 3863 21215 3915 21218
rect 3971 21215 4023 21218
rect 6239 21215 6291 21218
rect 6347 21215 6399 21218
rect 6455 21215 6507 21218
rect 6563 21215 6615 21218
rect 6671 21215 6723 21218
rect 8939 21215 8991 21218
rect 9047 21215 9099 21218
rect 11309 21215 11361 21218
rect 11417 21215 11469 21218
rect 1760 21020 1812 21023
rect 1868 21020 1920 21023
rect 1976 21020 2028 21023
rect 2084 21020 2136 21023
rect 2192 21020 2244 21023
rect 2300 21020 2352 21023
rect 2408 21020 2460 21023
rect 2516 21020 2568 21023
rect 2624 21020 2676 21023
rect 2732 21020 2784 21023
rect 2840 21020 2892 21023
rect 2948 21020 3000 21023
rect 3056 21020 3108 21023
rect 3164 21020 3216 21023
rect 3272 21020 3324 21023
rect 3380 21020 3432 21023
rect 3488 21020 3540 21023
rect 3596 21020 3648 21023
rect 3704 21020 3756 21023
rect 4130 21020 4182 21023
rect 4238 21020 4290 21023
rect 4346 21020 4398 21023
rect 4454 21020 4506 21023
rect 4562 21020 4614 21023
rect 4670 21020 4722 21023
rect 4778 21020 4830 21023
rect 4886 21020 4938 21023
rect 4994 21020 5046 21023
rect 5102 21020 5154 21023
rect 5210 21020 5262 21023
rect 5318 21020 5370 21023
rect 5426 21020 5478 21023
rect 5534 21020 5586 21023
rect 5642 21020 5694 21023
rect 5750 21020 5802 21023
rect 5858 21020 5910 21023
rect 5966 21020 6018 21023
rect 6074 21020 6126 21023
rect 6836 21020 6888 21023
rect 6944 21020 6996 21023
rect 7052 21020 7104 21023
rect 7160 21020 7212 21023
rect 7268 21020 7320 21023
rect 7376 21020 7428 21023
rect 7484 21020 7536 21023
rect 7592 21020 7644 21023
rect 7700 21020 7752 21023
rect 7808 21020 7860 21023
rect 7916 21020 7968 21023
rect 8024 21020 8076 21023
rect 8132 21020 8184 21023
rect 8240 21020 8292 21023
rect 8348 21020 8400 21023
rect 8456 21020 8508 21023
rect 8564 21020 8616 21023
rect 8672 21020 8724 21023
rect 8780 21020 8832 21023
rect 9206 21020 9258 21023
rect 9314 21020 9366 21023
rect 9422 21020 9474 21023
rect 9530 21020 9582 21023
rect 9638 21020 9690 21023
rect 9746 21020 9798 21023
rect 9854 21020 9906 21023
rect 9962 21020 10014 21023
rect 10070 21020 10122 21023
rect 10178 21020 10230 21023
rect 10286 21020 10338 21023
rect 10394 21020 10446 21023
rect 10502 21020 10554 21023
rect 10610 21020 10662 21023
rect 10718 21020 10770 21023
rect 10826 21020 10878 21023
rect 10934 21020 10986 21023
rect 11042 21020 11094 21023
rect 11150 21020 11202 21023
rect 1760 20974 1812 21020
rect 1868 20974 1920 21020
rect 1976 20974 2028 21020
rect 2084 20974 2136 21020
rect 2192 20974 2244 21020
rect 2300 20974 2352 21020
rect 2408 20974 2460 21020
rect 2516 20974 2568 21020
rect 2624 20974 2676 21020
rect 2732 20974 2784 21020
rect 2840 20974 2892 21020
rect 2948 20974 3000 21020
rect 3056 20974 3108 21020
rect 3164 20974 3216 21020
rect 3272 20974 3324 21020
rect 3380 20974 3432 21020
rect 3488 20974 3540 21020
rect 3596 20974 3648 21020
rect 3704 20974 3756 21020
rect 4130 20974 4182 21020
rect 4238 20974 4290 21020
rect 4346 20974 4398 21020
rect 4454 20974 4506 21020
rect 4562 20974 4614 21020
rect 4670 20974 4722 21020
rect 4778 20974 4830 21020
rect 4886 20974 4938 21020
rect 4994 20974 5046 21020
rect 5102 20974 5154 21020
rect 5210 20974 5262 21020
rect 5318 20974 5370 21020
rect 5426 20974 5478 21020
rect 5534 20974 5586 21020
rect 5642 20974 5694 21020
rect 5750 20974 5802 21020
rect 5858 20974 5910 21020
rect 5966 20974 6018 21020
rect 6074 20974 6126 21020
rect 6836 20974 6888 21020
rect 6944 20974 6996 21020
rect 7052 20974 7104 21020
rect 7160 20974 7212 21020
rect 7268 20974 7320 21020
rect 7376 20974 7428 21020
rect 7484 20974 7536 21020
rect 7592 20974 7644 21020
rect 7700 20974 7752 21020
rect 7808 20974 7860 21020
rect 7916 20974 7968 21020
rect 8024 20974 8076 21020
rect 8132 20974 8184 21020
rect 8240 20974 8292 21020
rect 8348 20974 8400 21020
rect 8456 20974 8508 21020
rect 8564 20974 8616 21020
rect 8672 20974 8724 21020
rect 8780 20974 8832 21020
rect 9206 20974 9258 21020
rect 9314 20974 9366 21020
rect 9422 20974 9474 21020
rect 9530 20974 9582 21020
rect 9638 20974 9690 21020
rect 9746 20974 9798 21020
rect 9854 20974 9906 21020
rect 9962 20974 10014 21020
rect 10070 20974 10122 21020
rect 10178 20974 10230 21020
rect 10286 20974 10338 21020
rect 10394 20974 10446 21020
rect 10502 20974 10554 21020
rect 10610 20974 10662 21020
rect 10718 20974 10770 21020
rect 10826 20974 10878 21020
rect 10934 20974 10986 21020
rect 11042 20974 11094 21020
rect 11150 20974 11202 21020
rect 1760 20971 1812 20974
rect 1868 20971 1920 20974
rect 1976 20971 2028 20974
rect 2084 20971 2136 20974
rect 2192 20971 2244 20974
rect 2300 20971 2352 20974
rect 2408 20971 2460 20974
rect 2516 20971 2568 20974
rect 2624 20971 2676 20974
rect 2732 20971 2784 20974
rect 2840 20971 2892 20974
rect 2948 20971 3000 20974
rect 3056 20971 3108 20974
rect 3164 20971 3216 20974
rect 3272 20971 3324 20974
rect 3380 20971 3432 20974
rect 3488 20971 3540 20974
rect 3596 20971 3648 20974
rect 3704 20971 3756 20974
rect 4130 20971 4182 20974
rect 4238 20971 4290 20974
rect 4346 20971 4398 20974
rect 4454 20971 4506 20974
rect 4562 20971 4614 20974
rect 4670 20971 4722 20974
rect 4778 20971 4830 20974
rect 4886 20971 4938 20974
rect 4994 20971 5046 20974
rect 5102 20971 5154 20974
rect 5210 20971 5262 20974
rect 5318 20971 5370 20974
rect 5426 20971 5478 20974
rect 5534 20971 5586 20974
rect 5642 20971 5694 20974
rect 5750 20971 5802 20974
rect 5858 20971 5910 20974
rect 5966 20971 6018 20974
rect 6074 20971 6126 20974
rect 6836 20971 6888 20974
rect 6944 20971 6996 20974
rect 7052 20971 7104 20974
rect 7160 20971 7212 20974
rect 7268 20971 7320 20974
rect 7376 20971 7428 20974
rect 7484 20971 7536 20974
rect 7592 20971 7644 20974
rect 7700 20971 7752 20974
rect 7808 20971 7860 20974
rect 7916 20971 7968 20974
rect 8024 20971 8076 20974
rect 8132 20971 8184 20974
rect 8240 20971 8292 20974
rect 8348 20971 8400 20974
rect 8456 20971 8508 20974
rect 8564 20971 8616 20974
rect 8672 20971 8724 20974
rect 8780 20971 8832 20974
rect 9206 20971 9258 20974
rect 9314 20971 9366 20974
rect 9422 20971 9474 20974
rect 9530 20971 9582 20974
rect 9638 20971 9690 20974
rect 9746 20971 9798 20974
rect 9854 20971 9906 20974
rect 9962 20971 10014 20974
rect 10070 20971 10122 20974
rect 10178 20971 10230 20974
rect 10286 20971 10338 20974
rect 10394 20971 10446 20974
rect 10502 20971 10554 20974
rect 10610 20971 10662 20974
rect 10718 20971 10770 20974
rect 10826 20971 10878 20974
rect 10934 20971 10986 20974
rect 11042 20971 11094 20974
rect 11150 20971 11202 20974
rect 1493 20776 1545 20779
rect 1601 20776 1653 20779
rect 3863 20776 3915 20779
rect 3971 20776 4023 20779
rect 6239 20776 6291 20779
rect 6347 20776 6399 20779
rect 6455 20776 6507 20779
rect 6563 20776 6615 20779
rect 6671 20776 6723 20779
rect 8939 20776 8991 20779
rect 9047 20776 9099 20779
rect 11309 20776 11361 20779
rect 11417 20776 11469 20779
rect 1493 20730 1494 20776
rect 1494 20730 1545 20776
rect 1601 20730 1653 20776
rect 3863 20730 3915 20776
rect 3971 20730 4023 20776
rect 6239 20730 6291 20776
rect 6347 20730 6399 20776
rect 6455 20730 6507 20776
rect 6563 20730 6615 20776
rect 6671 20730 6723 20776
rect 8939 20730 8991 20776
rect 9047 20730 9099 20776
rect 11309 20730 11361 20776
rect 11417 20730 11468 20776
rect 11468 20730 11469 20776
rect 1493 20727 1545 20730
rect 1601 20727 1653 20730
rect 3863 20727 3915 20730
rect 3971 20727 4023 20730
rect 6239 20727 6291 20730
rect 6347 20727 6399 20730
rect 6455 20727 6507 20730
rect 6563 20727 6615 20730
rect 6671 20727 6723 20730
rect 8939 20727 8991 20730
rect 9047 20727 9099 20730
rect 11309 20727 11361 20730
rect 11417 20727 11469 20730
rect 1760 20532 1812 20535
rect 1868 20532 1920 20535
rect 1976 20532 2028 20535
rect 2084 20532 2136 20535
rect 2192 20532 2244 20535
rect 2300 20532 2352 20535
rect 2408 20532 2460 20535
rect 2516 20532 2568 20535
rect 2624 20532 2676 20535
rect 2732 20532 2784 20535
rect 2840 20532 2892 20535
rect 2948 20532 3000 20535
rect 3056 20532 3108 20535
rect 3164 20532 3216 20535
rect 3272 20532 3324 20535
rect 3380 20532 3432 20535
rect 3488 20532 3540 20535
rect 3596 20532 3648 20535
rect 3704 20532 3756 20535
rect 4130 20532 4182 20535
rect 4238 20532 4290 20535
rect 4346 20532 4398 20535
rect 4454 20532 4506 20535
rect 4562 20532 4614 20535
rect 4670 20532 4722 20535
rect 4778 20532 4830 20535
rect 4886 20532 4938 20535
rect 4994 20532 5046 20535
rect 5102 20532 5154 20535
rect 5210 20532 5262 20535
rect 5318 20532 5370 20535
rect 5426 20532 5478 20535
rect 5534 20532 5586 20535
rect 5642 20532 5694 20535
rect 5750 20532 5802 20535
rect 5858 20532 5910 20535
rect 5966 20532 6018 20535
rect 6074 20532 6126 20535
rect 6836 20532 6888 20535
rect 6944 20532 6996 20535
rect 7052 20532 7104 20535
rect 7160 20532 7212 20535
rect 7268 20532 7320 20535
rect 7376 20532 7428 20535
rect 7484 20532 7536 20535
rect 7592 20532 7644 20535
rect 7700 20532 7752 20535
rect 7808 20532 7860 20535
rect 7916 20532 7968 20535
rect 8024 20532 8076 20535
rect 8132 20532 8184 20535
rect 8240 20532 8292 20535
rect 8348 20532 8400 20535
rect 8456 20532 8508 20535
rect 8564 20532 8616 20535
rect 8672 20532 8724 20535
rect 8780 20532 8832 20535
rect 9206 20532 9258 20535
rect 9314 20532 9366 20535
rect 9422 20532 9474 20535
rect 9530 20532 9582 20535
rect 9638 20532 9690 20535
rect 9746 20532 9798 20535
rect 9854 20532 9906 20535
rect 9962 20532 10014 20535
rect 10070 20532 10122 20535
rect 10178 20532 10230 20535
rect 10286 20532 10338 20535
rect 10394 20532 10446 20535
rect 10502 20532 10554 20535
rect 10610 20532 10662 20535
rect 10718 20532 10770 20535
rect 10826 20532 10878 20535
rect 10934 20532 10986 20535
rect 11042 20532 11094 20535
rect 11150 20532 11202 20535
rect 1760 20486 1812 20532
rect 1868 20486 1920 20532
rect 1976 20486 2028 20532
rect 2084 20486 2136 20532
rect 2192 20486 2244 20532
rect 2300 20486 2352 20532
rect 2408 20486 2460 20532
rect 2516 20486 2568 20532
rect 2624 20486 2676 20532
rect 2732 20486 2784 20532
rect 2840 20486 2892 20532
rect 2948 20486 3000 20532
rect 3056 20486 3108 20532
rect 3164 20486 3216 20532
rect 3272 20486 3324 20532
rect 3380 20486 3432 20532
rect 3488 20486 3540 20532
rect 3596 20486 3648 20532
rect 3704 20486 3756 20532
rect 4130 20486 4182 20532
rect 4238 20486 4290 20532
rect 4346 20486 4398 20532
rect 4454 20486 4506 20532
rect 4562 20486 4614 20532
rect 4670 20486 4722 20532
rect 4778 20486 4830 20532
rect 4886 20486 4938 20532
rect 4994 20486 5046 20532
rect 5102 20486 5154 20532
rect 5210 20486 5262 20532
rect 5318 20486 5370 20532
rect 5426 20486 5478 20532
rect 5534 20486 5586 20532
rect 5642 20486 5694 20532
rect 5750 20486 5802 20532
rect 5858 20486 5910 20532
rect 5966 20486 6018 20532
rect 6074 20486 6126 20532
rect 6836 20486 6888 20532
rect 6944 20486 6996 20532
rect 7052 20486 7104 20532
rect 7160 20486 7212 20532
rect 7268 20486 7320 20532
rect 7376 20486 7428 20532
rect 7484 20486 7536 20532
rect 7592 20486 7644 20532
rect 7700 20486 7752 20532
rect 7808 20486 7860 20532
rect 7916 20486 7968 20532
rect 8024 20486 8076 20532
rect 8132 20486 8184 20532
rect 8240 20486 8292 20532
rect 8348 20486 8400 20532
rect 8456 20486 8508 20532
rect 8564 20486 8616 20532
rect 8672 20486 8724 20532
rect 8780 20486 8832 20532
rect 9206 20486 9258 20532
rect 9314 20486 9366 20532
rect 9422 20486 9474 20532
rect 9530 20486 9582 20532
rect 9638 20486 9690 20532
rect 9746 20486 9798 20532
rect 9854 20486 9906 20532
rect 9962 20486 10014 20532
rect 10070 20486 10122 20532
rect 10178 20486 10230 20532
rect 10286 20486 10338 20532
rect 10394 20486 10446 20532
rect 10502 20486 10554 20532
rect 10610 20486 10662 20532
rect 10718 20486 10770 20532
rect 10826 20486 10878 20532
rect 10934 20486 10986 20532
rect 11042 20486 11094 20532
rect 11150 20486 11202 20532
rect 1760 20483 1812 20486
rect 1868 20483 1920 20486
rect 1976 20483 2028 20486
rect 2084 20483 2136 20486
rect 2192 20483 2244 20486
rect 2300 20483 2352 20486
rect 2408 20483 2460 20486
rect 2516 20483 2568 20486
rect 2624 20483 2676 20486
rect 2732 20483 2784 20486
rect 2840 20483 2892 20486
rect 2948 20483 3000 20486
rect 3056 20483 3108 20486
rect 3164 20483 3216 20486
rect 3272 20483 3324 20486
rect 3380 20483 3432 20486
rect 3488 20483 3540 20486
rect 3596 20483 3648 20486
rect 3704 20483 3756 20486
rect 4130 20483 4182 20486
rect 4238 20483 4290 20486
rect 4346 20483 4398 20486
rect 4454 20483 4506 20486
rect 4562 20483 4614 20486
rect 4670 20483 4722 20486
rect 4778 20483 4830 20486
rect 4886 20483 4938 20486
rect 4994 20483 5046 20486
rect 5102 20483 5154 20486
rect 5210 20483 5262 20486
rect 5318 20483 5370 20486
rect 5426 20483 5478 20486
rect 5534 20483 5586 20486
rect 5642 20483 5694 20486
rect 5750 20483 5802 20486
rect 5858 20483 5910 20486
rect 5966 20483 6018 20486
rect 6074 20483 6126 20486
rect 6836 20483 6888 20486
rect 6944 20483 6996 20486
rect 7052 20483 7104 20486
rect 7160 20483 7212 20486
rect 7268 20483 7320 20486
rect 7376 20483 7428 20486
rect 7484 20483 7536 20486
rect 7592 20483 7644 20486
rect 7700 20483 7752 20486
rect 7808 20483 7860 20486
rect 7916 20483 7968 20486
rect 8024 20483 8076 20486
rect 8132 20483 8184 20486
rect 8240 20483 8292 20486
rect 8348 20483 8400 20486
rect 8456 20483 8508 20486
rect 8564 20483 8616 20486
rect 8672 20483 8724 20486
rect 8780 20483 8832 20486
rect 9206 20483 9258 20486
rect 9314 20483 9366 20486
rect 9422 20483 9474 20486
rect 9530 20483 9582 20486
rect 9638 20483 9690 20486
rect 9746 20483 9798 20486
rect 9854 20483 9906 20486
rect 9962 20483 10014 20486
rect 10070 20483 10122 20486
rect 10178 20483 10230 20486
rect 10286 20483 10338 20486
rect 10394 20483 10446 20486
rect 10502 20483 10554 20486
rect 10610 20483 10662 20486
rect 10718 20483 10770 20486
rect 10826 20483 10878 20486
rect 10934 20483 10986 20486
rect 11042 20483 11094 20486
rect 11150 20483 11202 20486
rect 1493 20288 1545 20291
rect 1601 20288 1653 20291
rect 3863 20288 3915 20291
rect 3971 20288 4023 20291
rect 6239 20288 6291 20291
rect 6347 20288 6399 20291
rect 6455 20288 6507 20291
rect 6563 20288 6615 20291
rect 6671 20288 6723 20291
rect 8939 20288 8991 20291
rect 9047 20288 9099 20291
rect 11309 20288 11361 20291
rect 11417 20288 11469 20291
rect 1493 20242 1494 20288
rect 1494 20242 1545 20288
rect 1601 20242 1653 20288
rect 3863 20242 3915 20288
rect 3971 20242 4023 20288
rect 6239 20242 6291 20288
rect 6347 20242 6399 20288
rect 6455 20242 6507 20288
rect 6563 20242 6615 20288
rect 6671 20242 6723 20288
rect 8939 20242 8991 20288
rect 9047 20242 9099 20288
rect 11309 20242 11361 20288
rect 11417 20242 11468 20288
rect 11468 20242 11469 20288
rect 1493 20239 1545 20242
rect 1601 20239 1653 20242
rect 3863 20239 3915 20242
rect 3971 20239 4023 20242
rect 6239 20239 6291 20242
rect 6347 20239 6399 20242
rect 6455 20239 6507 20242
rect 6563 20239 6615 20242
rect 6671 20239 6723 20242
rect 8939 20239 8991 20242
rect 9047 20239 9099 20242
rect 11309 20239 11361 20242
rect 11417 20239 11469 20242
rect 1760 20044 1812 20047
rect 1868 20044 1920 20047
rect 1976 20044 2028 20047
rect 2084 20044 2136 20047
rect 2192 20044 2244 20047
rect 2300 20044 2352 20047
rect 2408 20044 2460 20047
rect 2516 20044 2568 20047
rect 2624 20044 2676 20047
rect 2732 20044 2784 20047
rect 2840 20044 2892 20047
rect 2948 20044 3000 20047
rect 3056 20044 3108 20047
rect 3164 20044 3216 20047
rect 3272 20044 3324 20047
rect 3380 20044 3432 20047
rect 3488 20044 3540 20047
rect 3596 20044 3648 20047
rect 3704 20044 3756 20047
rect 4130 20044 4182 20047
rect 4238 20044 4290 20047
rect 4346 20044 4398 20047
rect 4454 20044 4506 20047
rect 4562 20044 4614 20047
rect 4670 20044 4722 20047
rect 4778 20044 4830 20047
rect 4886 20044 4938 20047
rect 4994 20044 5046 20047
rect 5102 20044 5154 20047
rect 5210 20044 5262 20047
rect 5318 20044 5370 20047
rect 5426 20044 5478 20047
rect 5534 20044 5586 20047
rect 5642 20044 5694 20047
rect 5750 20044 5802 20047
rect 5858 20044 5910 20047
rect 5966 20044 6018 20047
rect 6074 20044 6126 20047
rect 6836 20044 6888 20047
rect 6944 20044 6996 20047
rect 7052 20044 7104 20047
rect 7160 20044 7212 20047
rect 7268 20044 7320 20047
rect 7376 20044 7428 20047
rect 7484 20044 7536 20047
rect 7592 20044 7644 20047
rect 7700 20044 7752 20047
rect 7808 20044 7860 20047
rect 7916 20044 7968 20047
rect 8024 20044 8076 20047
rect 8132 20044 8184 20047
rect 8240 20044 8292 20047
rect 8348 20044 8400 20047
rect 8456 20044 8508 20047
rect 8564 20044 8616 20047
rect 8672 20044 8724 20047
rect 8780 20044 8832 20047
rect 9206 20044 9258 20047
rect 9314 20044 9366 20047
rect 9422 20044 9474 20047
rect 9530 20044 9582 20047
rect 9638 20044 9690 20047
rect 9746 20044 9798 20047
rect 9854 20044 9906 20047
rect 9962 20044 10014 20047
rect 10070 20044 10122 20047
rect 10178 20044 10230 20047
rect 10286 20044 10338 20047
rect 10394 20044 10446 20047
rect 10502 20044 10554 20047
rect 10610 20044 10662 20047
rect 10718 20044 10770 20047
rect 10826 20044 10878 20047
rect 10934 20044 10986 20047
rect 11042 20044 11094 20047
rect 11150 20044 11202 20047
rect 1760 19998 1812 20044
rect 1868 19998 1920 20044
rect 1976 19998 2028 20044
rect 2084 19998 2136 20044
rect 2192 19998 2244 20044
rect 2300 19998 2352 20044
rect 2408 19998 2460 20044
rect 2516 19998 2568 20044
rect 2624 19998 2676 20044
rect 2732 19998 2784 20044
rect 2840 19998 2892 20044
rect 2948 19998 3000 20044
rect 3056 19998 3108 20044
rect 3164 19998 3216 20044
rect 3272 19998 3324 20044
rect 3380 19998 3432 20044
rect 3488 19998 3540 20044
rect 3596 19998 3648 20044
rect 3704 19998 3756 20044
rect 4130 19998 4182 20044
rect 4238 19998 4290 20044
rect 4346 19998 4398 20044
rect 4454 19998 4506 20044
rect 4562 19998 4614 20044
rect 4670 19998 4722 20044
rect 4778 19998 4830 20044
rect 4886 19998 4938 20044
rect 4994 19998 5046 20044
rect 5102 19998 5154 20044
rect 5210 19998 5262 20044
rect 5318 19998 5370 20044
rect 5426 19998 5478 20044
rect 5534 19998 5586 20044
rect 5642 19998 5694 20044
rect 5750 19998 5802 20044
rect 5858 19998 5910 20044
rect 5966 19998 6018 20044
rect 6074 19998 6126 20044
rect 6836 19998 6888 20044
rect 6944 19998 6996 20044
rect 7052 19998 7104 20044
rect 7160 19998 7212 20044
rect 7268 19998 7320 20044
rect 7376 19998 7428 20044
rect 7484 19998 7536 20044
rect 7592 19998 7644 20044
rect 7700 19998 7752 20044
rect 7808 19998 7860 20044
rect 7916 19998 7968 20044
rect 8024 19998 8076 20044
rect 8132 19998 8184 20044
rect 8240 19998 8292 20044
rect 8348 19998 8400 20044
rect 8456 19998 8508 20044
rect 8564 19998 8616 20044
rect 8672 19998 8724 20044
rect 8780 19998 8832 20044
rect 9206 19998 9258 20044
rect 9314 19998 9366 20044
rect 9422 19998 9474 20044
rect 9530 19998 9582 20044
rect 9638 19998 9690 20044
rect 9746 19998 9798 20044
rect 9854 19998 9906 20044
rect 9962 19998 10014 20044
rect 10070 19998 10122 20044
rect 10178 19998 10230 20044
rect 10286 19998 10338 20044
rect 10394 19998 10446 20044
rect 10502 19998 10554 20044
rect 10610 19998 10662 20044
rect 10718 19998 10770 20044
rect 10826 19998 10878 20044
rect 10934 19998 10986 20044
rect 11042 19998 11094 20044
rect 11150 19998 11202 20044
rect 1760 19995 1812 19998
rect 1868 19995 1920 19998
rect 1976 19995 2028 19998
rect 2084 19995 2136 19998
rect 2192 19995 2244 19998
rect 2300 19995 2352 19998
rect 2408 19995 2460 19998
rect 2516 19995 2568 19998
rect 2624 19995 2676 19998
rect 2732 19995 2784 19998
rect 2840 19995 2892 19998
rect 2948 19995 3000 19998
rect 3056 19995 3108 19998
rect 3164 19995 3216 19998
rect 3272 19995 3324 19998
rect 3380 19995 3432 19998
rect 3488 19995 3540 19998
rect 3596 19995 3648 19998
rect 3704 19995 3756 19998
rect 4130 19995 4182 19998
rect 4238 19995 4290 19998
rect 4346 19995 4398 19998
rect 4454 19995 4506 19998
rect 4562 19995 4614 19998
rect 4670 19995 4722 19998
rect 4778 19995 4830 19998
rect 4886 19995 4938 19998
rect 4994 19995 5046 19998
rect 5102 19995 5154 19998
rect 5210 19995 5262 19998
rect 5318 19995 5370 19998
rect 5426 19995 5478 19998
rect 5534 19995 5586 19998
rect 5642 19995 5694 19998
rect 5750 19995 5802 19998
rect 5858 19995 5910 19998
rect 5966 19995 6018 19998
rect 6074 19995 6126 19998
rect 6836 19995 6888 19998
rect 6944 19995 6996 19998
rect 7052 19995 7104 19998
rect 7160 19995 7212 19998
rect 7268 19995 7320 19998
rect 7376 19995 7428 19998
rect 7484 19995 7536 19998
rect 7592 19995 7644 19998
rect 7700 19995 7752 19998
rect 7808 19995 7860 19998
rect 7916 19995 7968 19998
rect 8024 19995 8076 19998
rect 8132 19995 8184 19998
rect 8240 19995 8292 19998
rect 8348 19995 8400 19998
rect 8456 19995 8508 19998
rect 8564 19995 8616 19998
rect 8672 19995 8724 19998
rect 8780 19995 8832 19998
rect 9206 19995 9258 19998
rect 9314 19995 9366 19998
rect 9422 19995 9474 19998
rect 9530 19995 9582 19998
rect 9638 19995 9690 19998
rect 9746 19995 9798 19998
rect 9854 19995 9906 19998
rect 9962 19995 10014 19998
rect 10070 19995 10122 19998
rect 10178 19995 10230 19998
rect 10286 19995 10338 19998
rect 10394 19995 10446 19998
rect 10502 19995 10554 19998
rect 10610 19995 10662 19998
rect 10718 19995 10770 19998
rect 10826 19995 10878 19998
rect 10934 19995 10986 19998
rect 11042 19995 11094 19998
rect 11150 19995 11202 19998
rect 1493 19800 1545 19803
rect 1601 19800 1653 19803
rect 3863 19800 3915 19803
rect 3971 19800 4023 19803
rect 6239 19800 6291 19803
rect 6347 19800 6399 19803
rect 6455 19800 6507 19803
rect 6563 19800 6615 19803
rect 6671 19800 6723 19803
rect 8939 19800 8991 19803
rect 9047 19800 9099 19803
rect 11309 19800 11361 19803
rect 11417 19800 11469 19803
rect 1493 19754 1494 19800
rect 1494 19754 1545 19800
rect 1601 19754 1653 19800
rect 3863 19754 3915 19800
rect 3971 19754 4023 19800
rect 6239 19754 6291 19800
rect 6347 19754 6399 19800
rect 6455 19754 6507 19800
rect 6563 19754 6615 19800
rect 6671 19754 6723 19800
rect 8939 19754 8991 19800
rect 9047 19754 9099 19800
rect 11309 19754 11361 19800
rect 11417 19754 11468 19800
rect 11468 19754 11469 19800
rect 1493 19751 1545 19754
rect 1601 19751 1653 19754
rect 3863 19751 3915 19754
rect 3971 19751 4023 19754
rect 6239 19751 6291 19754
rect 6347 19751 6399 19754
rect 6455 19751 6507 19754
rect 6563 19751 6615 19754
rect 6671 19751 6723 19754
rect 8939 19751 8991 19754
rect 9047 19751 9099 19754
rect 11309 19751 11361 19754
rect 11417 19751 11469 19754
rect 1760 19556 1812 19559
rect 1868 19556 1920 19559
rect 1976 19556 2028 19559
rect 2084 19556 2136 19559
rect 2192 19556 2244 19559
rect 2300 19556 2352 19559
rect 2408 19556 2460 19559
rect 2516 19556 2568 19559
rect 2624 19556 2676 19559
rect 2732 19556 2784 19559
rect 2840 19556 2892 19559
rect 2948 19556 3000 19559
rect 3056 19556 3108 19559
rect 3164 19556 3216 19559
rect 3272 19556 3324 19559
rect 3380 19556 3432 19559
rect 3488 19556 3540 19559
rect 3596 19556 3648 19559
rect 3704 19556 3756 19559
rect 4130 19556 4182 19559
rect 4238 19556 4290 19559
rect 4346 19556 4398 19559
rect 4454 19556 4506 19559
rect 4562 19556 4614 19559
rect 4670 19556 4722 19559
rect 4778 19556 4830 19559
rect 4886 19556 4938 19559
rect 4994 19556 5046 19559
rect 5102 19556 5154 19559
rect 5210 19556 5262 19559
rect 5318 19556 5370 19559
rect 5426 19556 5478 19559
rect 5534 19556 5586 19559
rect 5642 19556 5694 19559
rect 5750 19556 5802 19559
rect 5858 19556 5910 19559
rect 5966 19556 6018 19559
rect 6074 19556 6126 19559
rect 6836 19556 6888 19559
rect 6944 19556 6996 19559
rect 7052 19556 7104 19559
rect 7160 19556 7212 19559
rect 7268 19556 7320 19559
rect 7376 19556 7428 19559
rect 7484 19556 7536 19559
rect 7592 19556 7644 19559
rect 7700 19556 7752 19559
rect 7808 19556 7860 19559
rect 7916 19556 7968 19559
rect 8024 19556 8076 19559
rect 8132 19556 8184 19559
rect 8240 19556 8292 19559
rect 8348 19556 8400 19559
rect 8456 19556 8508 19559
rect 8564 19556 8616 19559
rect 8672 19556 8724 19559
rect 8780 19556 8832 19559
rect 9206 19556 9258 19559
rect 9314 19556 9366 19559
rect 9422 19556 9474 19559
rect 9530 19556 9582 19559
rect 9638 19556 9690 19559
rect 9746 19556 9798 19559
rect 9854 19556 9906 19559
rect 9962 19556 10014 19559
rect 10070 19556 10122 19559
rect 10178 19556 10230 19559
rect 10286 19556 10338 19559
rect 10394 19556 10446 19559
rect 10502 19556 10554 19559
rect 10610 19556 10662 19559
rect 10718 19556 10770 19559
rect 10826 19556 10878 19559
rect 10934 19556 10986 19559
rect 11042 19556 11094 19559
rect 11150 19556 11202 19559
rect 1760 19510 1812 19556
rect 1868 19510 1920 19556
rect 1976 19510 2028 19556
rect 2084 19510 2136 19556
rect 2192 19510 2244 19556
rect 2300 19510 2352 19556
rect 2408 19510 2460 19556
rect 2516 19510 2568 19556
rect 2624 19510 2676 19556
rect 2732 19510 2784 19556
rect 2840 19510 2892 19556
rect 2948 19510 3000 19556
rect 3056 19510 3108 19556
rect 3164 19510 3216 19556
rect 3272 19510 3324 19556
rect 3380 19510 3432 19556
rect 3488 19510 3540 19556
rect 3596 19510 3648 19556
rect 3704 19510 3756 19556
rect 4130 19510 4182 19556
rect 4238 19510 4290 19556
rect 4346 19510 4398 19556
rect 4454 19510 4506 19556
rect 4562 19510 4614 19556
rect 4670 19510 4722 19556
rect 4778 19510 4830 19556
rect 4886 19510 4938 19556
rect 4994 19510 5046 19556
rect 5102 19510 5154 19556
rect 5210 19510 5262 19556
rect 5318 19510 5370 19556
rect 5426 19510 5478 19556
rect 5534 19510 5586 19556
rect 5642 19510 5694 19556
rect 5750 19510 5802 19556
rect 5858 19510 5910 19556
rect 5966 19510 6018 19556
rect 6074 19510 6126 19556
rect 6836 19510 6888 19556
rect 6944 19510 6996 19556
rect 7052 19510 7104 19556
rect 7160 19510 7212 19556
rect 7268 19510 7320 19556
rect 7376 19510 7428 19556
rect 7484 19510 7536 19556
rect 7592 19510 7644 19556
rect 7700 19510 7752 19556
rect 7808 19510 7860 19556
rect 7916 19510 7968 19556
rect 8024 19510 8076 19556
rect 8132 19510 8184 19556
rect 8240 19510 8292 19556
rect 8348 19510 8400 19556
rect 8456 19510 8508 19556
rect 8564 19510 8616 19556
rect 8672 19510 8724 19556
rect 8780 19510 8832 19556
rect 9206 19510 9258 19556
rect 9314 19510 9366 19556
rect 9422 19510 9474 19556
rect 9530 19510 9582 19556
rect 9638 19510 9690 19556
rect 9746 19510 9798 19556
rect 9854 19510 9906 19556
rect 9962 19510 10014 19556
rect 10070 19510 10122 19556
rect 10178 19510 10230 19556
rect 10286 19510 10338 19556
rect 10394 19510 10446 19556
rect 10502 19510 10554 19556
rect 10610 19510 10662 19556
rect 10718 19510 10770 19556
rect 10826 19510 10878 19556
rect 10934 19510 10986 19556
rect 11042 19510 11094 19556
rect 11150 19510 11202 19556
rect 1760 19507 1812 19510
rect 1868 19507 1920 19510
rect 1976 19507 2028 19510
rect 2084 19507 2136 19510
rect 2192 19507 2244 19510
rect 2300 19507 2352 19510
rect 2408 19507 2460 19510
rect 2516 19507 2568 19510
rect 2624 19507 2676 19510
rect 2732 19507 2784 19510
rect 2840 19507 2892 19510
rect 2948 19507 3000 19510
rect 3056 19507 3108 19510
rect 3164 19507 3216 19510
rect 3272 19507 3324 19510
rect 3380 19507 3432 19510
rect 3488 19507 3540 19510
rect 3596 19507 3648 19510
rect 3704 19507 3756 19510
rect 4130 19507 4182 19510
rect 4238 19507 4290 19510
rect 4346 19507 4398 19510
rect 4454 19507 4506 19510
rect 4562 19507 4614 19510
rect 4670 19507 4722 19510
rect 4778 19507 4830 19510
rect 4886 19507 4938 19510
rect 4994 19507 5046 19510
rect 5102 19507 5154 19510
rect 5210 19507 5262 19510
rect 5318 19507 5370 19510
rect 5426 19507 5478 19510
rect 5534 19507 5586 19510
rect 5642 19507 5694 19510
rect 5750 19507 5802 19510
rect 5858 19507 5910 19510
rect 5966 19507 6018 19510
rect 6074 19507 6126 19510
rect 6836 19507 6888 19510
rect 6944 19507 6996 19510
rect 7052 19507 7104 19510
rect 7160 19507 7212 19510
rect 7268 19507 7320 19510
rect 7376 19507 7428 19510
rect 7484 19507 7536 19510
rect 7592 19507 7644 19510
rect 7700 19507 7752 19510
rect 7808 19507 7860 19510
rect 7916 19507 7968 19510
rect 8024 19507 8076 19510
rect 8132 19507 8184 19510
rect 8240 19507 8292 19510
rect 8348 19507 8400 19510
rect 8456 19507 8508 19510
rect 8564 19507 8616 19510
rect 8672 19507 8724 19510
rect 8780 19507 8832 19510
rect 9206 19507 9258 19510
rect 9314 19507 9366 19510
rect 9422 19507 9474 19510
rect 9530 19507 9582 19510
rect 9638 19507 9690 19510
rect 9746 19507 9798 19510
rect 9854 19507 9906 19510
rect 9962 19507 10014 19510
rect 10070 19507 10122 19510
rect 10178 19507 10230 19510
rect 10286 19507 10338 19510
rect 10394 19507 10446 19510
rect 10502 19507 10554 19510
rect 10610 19507 10662 19510
rect 10718 19507 10770 19510
rect 10826 19507 10878 19510
rect 10934 19507 10986 19510
rect 11042 19507 11094 19510
rect 11150 19507 11202 19510
rect 1493 19312 1545 19315
rect 1601 19312 1653 19315
rect 3863 19312 3915 19315
rect 3971 19312 4023 19315
rect 6239 19312 6291 19315
rect 6347 19312 6399 19315
rect 6455 19312 6507 19315
rect 6563 19312 6615 19315
rect 6671 19312 6723 19315
rect 8939 19312 8991 19315
rect 9047 19312 9099 19315
rect 11309 19312 11361 19315
rect 11417 19312 11469 19315
rect 1493 19266 1494 19312
rect 1494 19266 1545 19312
rect 1601 19266 1653 19312
rect 3863 19266 3915 19312
rect 3971 19266 4023 19312
rect 6239 19266 6291 19312
rect 6347 19266 6399 19312
rect 6455 19266 6507 19312
rect 6563 19266 6615 19312
rect 6671 19266 6723 19312
rect 8939 19266 8991 19312
rect 9047 19266 9099 19312
rect 11309 19266 11361 19312
rect 11417 19266 11468 19312
rect 11468 19266 11469 19312
rect 1493 19263 1545 19266
rect 1601 19263 1653 19266
rect 3863 19263 3915 19266
rect 3971 19263 4023 19266
rect 6239 19263 6291 19266
rect 6347 19263 6399 19266
rect 6455 19263 6507 19266
rect 6563 19263 6615 19266
rect 6671 19263 6723 19266
rect 8939 19263 8991 19266
rect 9047 19263 9099 19266
rect 11309 19263 11361 19266
rect 11417 19263 11469 19266
rect 1233 19083 1285 19135
rect 1341 19083 1393 19135
rect 11569 23727 11621 23779
rect 11677 23727 11706 23779
rect 11706 23727 11729 23779
rect 11569 23619 11621 23671
rect 11677 23619 11706 23671
rect 11706 23619 11729 23671
rect 11569 23511 11621 23563
rect 11677 23511 11706 23563
rect 11706 23511 11729 23563
rect 11569 23403 11621 23455
rect 11677 23403 11706 23455
rect 11706 23403 11729 23455
rect 11569 23295 11621 23347
rect 11677 23295 11706 23347
rect 11706 23295 11729 23347
rect 11569 23187 11621 23239
rect 11677 23187 11706 23239
rect 11706 23187 11729 23239
rect 11569 23079 11621 23131
rect 11677 23079 11706 23131
rect 11706 23079 11729 23131
rect 11569 22971 11621 23023
rect 11677 22971 11706 23023
rect 11706 22971 11729 23023
rect 11569 22863 11621 22915
rect 11677 22863 11706 22915
rect 11706 22863 11729 22915
rect 11569 22755 11621 22807
rect 11677 22755 11706 22807
rect 11706 22755 11729 22807
rect 11569 22647 11621 22699
rect 11677 22647 11706 22699
rect 11706 22647 11729 22699
rect 11569 22539 11621 22591
rect 11677 22539 11706 22591
rect 11706 22539 11729 22591
rect 11569 22431 11621 22483
rect 11677 22431 11706 22483
rect 11706 22431 11729 22483
rect 11569 22323 11621 22375
rect 11677 22323 11706 22375
rect 11706 22323 11729 22375
rect 11569 22215 11621 22267
rect 11677 22215 11706 22267
rect 11706 22215 11729 22267
rect 11569 22107 11621 22159
rect 11677 22107 11706 22159
rect 11706 22107 11729 22159
rect 11569 21999 11621 22051
rect 11677 21999 11706 22051
rect 11706 21999 11729 22051
rect 11569 21891 11621 21943
rect 11677 21891 11706 21943
rect 11706 21891 11729 21943
rect 11569 21783 11621 21835
rect 11677 21783 11706 21835
rect 11706 21783 11729 21835
rect 11569 21675 11621 21727
rect 11677 21675 11706 21727
rect 11706 21675 11729 21727
rect 11569 21567 11621 21619
rect 11677 21567 11706 21619
rect 11706 21567 11729 21619
rect 11569 21459 11621 21511
rect 11677 21459 11706 21511
rect 11706 21459 11729 21511
rect 11569 21351 11621 21403
rect 11677 21351 11706 21403
rect 11706 21351 11729 21403
rect 11569 21243 11621 21295
rect 11677 21243 11706 21295
rect 11706 21243 11729 21295
rect 11569 21135 11621 21187
rect 11677 21135 11706 21187
rect 11706 21135 11729 21187
rect 11569 21027 11621 21079
rect 11677 21027 11706 21079
rect 11706 21027 11729 21079
rect 11569 20919 11621 20971
rect 11677 20919 11706 20971
rect 11706 20919 11729 20971
rect 11569 20811 11621 20863
rect 11677 20811 11706 20863
rect 11706 20811 11729 20863
rect 11569 20703 11621 20755
rect 11677 20703 11706 20755
rect 11706 20703 11729 20755
rect 11569 20595 11621 20647
rect 11677 20595 11706 20647
rect 11706 20595 11729 20647
rect 11569 20487 11621 20539
rect 11677 20487 11706 20539
rect 11706 20487 11729 20539
rect 11569 20379 11621 20431
rect 11677 20379 11706 20431
rect 11706 20379 11729 20431
rect 11569 20271 11621 20323
rect 11677 20271 11706 20323
rect 11706 20271 11729 20323
rect 11569 20163 11621 20215
rect 11677 20163 11706 20215
rect 11706 20163 11729 20215
rect 11569 20055 11621 20107
rect 11677 20055 11706 20107
rect 11706 20055 11729 20107
rect 11569 19947 11621 19999
rect 11677 19947 11706 19999
rect 11706 19947 11729 19999
rect 11569 19839 11621 19891
rect 11677 19839 11706 19891
rect 11706 19839 11729 19891
rect 11569 19731 11621 19783
rect 11677 19731 11706 19783
rect 11706 19731 11729 19783
rect 11569 19623 11621 19675
rect 11677 19623 11706 19675
rect 11706 19623 11729 19675
rect 11569 19515 11621 19567
rect 11677 19515 11706 19567
rect 11706 19515 11729 19567
rect 11569 19407 11621 19459
rect 11677 19407 11706 19459
rect 11706 19407 11729 19459
rect 11569 19299 11621 19351
rect 11677 19299 11706 19351
rect 11706 19299 11729 19351
rect 11569 19191 11621 19243
rect 11677 19191 11706 19243
rect 11706 19191 11729 19243
rect 11569 19083 11621 19135
rect 11677 19083 11729 19135
rect 1760 19068 1812 19071
rect 1868 19068 1920 19071
rect 1976 19068 2028 19071
rect 2084 19068 2136 19071
rect 2192 19068 2244 19071
rect 2300 19068 2352 19071
rect 2408 19068 2460 19071
rect 2516 19068 2568 19071
rect 2624 19068 2676 19071
rect 2732 19068 2784 19071
rect 2840 19068 2892 19071
rect 2948 19068 3000 19071
rect 3056 19068 3108 19071
rect 3164 19068 3216 19071
rect 3272 19068 3324 19071
rect 3380 19068 3432 19071
rect 3488 19068 3540 19071
rect 3596 19068 3648 19071
rect 3704 19068 3756 19071
rect 4130 19068 4182 19071
rect 4238 19068 4290 19071
rect 4346 19068 4398 19071
rect 4454 19068 4506 19071
rect 4562 19068 4614 19071
rect 4670 19068 4722 19071
rect 4778 19068 4830 19071
rect 4886 19068 4938 19071
rect 4994 19068 5046 19071
rect 5102 19068 5154 19071
rect 5210 19068 5262 19071
rect 5318 19068 5370 19071
rect 5426 19068 5478 19071
rect 5534 19068 5586 19071
rect 5642 19068 5694 19071
rect 5750 19068 5802 19071
rect 5858 19068 5910 19071
rect 5966 19068 6018 19071
rect 6074 19068 6126 19071
rect 6836 19068 6888 19071
rect 6944 19068 6996 19071
rect 7052 19068 7104 19071
rect 7160 19068 7212 19071
rect 7268 19068 7320 19071
rect 7376 19068 7428 19071
rect 7484 19068 7536 19071
rect 7592 19068 7644 19071
rect 7700 19068 7752 19071
rect 7808 19068 7860 19071
rect 7916 19068 7968 19071
rect 8024 19068 8076 19071
rect 8132 19068 8184 19071
rect 8240 19068 8292 19071
rect 8348 19068 8400 19071
rect 8456 19068 8508 19071
rect 8564 19068 8616 19071
rect 8672 19068 8724 19071
rect 8780 19068 8832 19071
rect 9206 19068 9258 19071
rect 9314 19068 9366 19071
rect 9422 19068 9474 19071
rect 9530 19068 9582 19071
rect 9638 19068 9690 19071
rect 9746 19068 9798 19071
rect 9854 19068 9906 19071
rect 9962 19068 10014 19071
rect 10070 19068 10122 19071
rect 10178 19068 10230 19071
rect 10286 19068 10338 19071
rect 10394 19068 10446 19071
rect 10502 19068 10554 19071
rect 10610 19068 10662 19071
rect 10718 19068 10770 19071
rect 10826 19068 10878 19071
rect 10934 19068 10986 19071
rect 11042 19068 11094 19071
rect 11150 19068 11202 19071
rect 1760 19022 1812 19068
rect 1868 19022 1920 19068
rect 1976 19022 2028 19068
rect 2084 19022 2136 19068
rect 2192 19022 2244 19068
rect 2300 19022 2352 19068
rect 2408 19022 2460 19068
rect 2516 19022 2568 19068
rect 2624 19022 2676 19068
rect 2732 19022 2784 19068
rect 2840 19022 2892 19068
rect 2948 19022 3000 19068
rect 3056 19022 3108 19068
rect 3164 19022 3216 19068
rect 3272 19022 3324 19068
rect 3380 19022 3432 19068
rect 3488 19022 3540 19068
rect 3596 19022 3648 19068
rect 3704 19022 3756 19068
rect 4130 19022 4182 19068
rect 4238 19022 4290 19068
rect 4346 19022 4398 19068
rect 4454 19022 4506 19068
rect 4562 19022 4614 19068
rect 4670 19022 4722 19068
rect 4778 19022 4830 19068
rect 4886 19022 4938 19068
rect 4994 19022 5046 19068
rect 5102 19022 5154 19068
rect 5210 19022 5262 19068
rect 5318 19022 5370 19068
rect 5426 19022 5478 19068
rect 5534 19022 5586 19068
rect 5642 19022 5694 19068
rect 5750 19022 5802 19068
rect 5858 19022 5910 19068
rect 5966 19022 6018 19068
rect 6074 19022 6126 19068
rect 6836 19022 6888 19068
rect 6944 19022 6996 19068
rect 7052 19022 7104 19068
rect 7160 19022 7212 19068
rect 7268 19022 7320 19068
rect 7376 19022 7428 19068
rect 7484 19022 7536 19068
rect 7592 19022 7644 19068
rect 7700 19022 7752 19068
rect 7808 19022 7860 19068
rect 7916 19022 7968 19068
rect 8024 19022 8076 19068
rect 8132 19022 8184 19068
rect 8240 19022 8292 19068
rect 8348 19022 8400 19068
rect 8456 19022 8508 19068
rect 8564 19022 8616 19068
rect 8672 19022 8724 19068
rect 8780 19022 8832 19068
rect 9206 19022 9258 19068
rect 9314 19022 9366 19068
rect 9422 19022 9474 19068
rect 9530 19022 9582 19068
rect 9638 19022 9690 19068
rect 9746 19022 9798 19068
rect 9854 19022 9906 19068
rect 9962 19022 10014 19068
rect 10070 19022 10122 19068
rect 10178 19022 10230 19068
rect 10286 19022 10338 19068
rect 10394 19022 10446 19068
rect 10502 19022 10554 19068
rect 10610 19022 10662 19068
rect 10718 19022 10770 19068
rect 10826 19022 10878 19068
rect 10934 19022 10986 19068
rect 11042 19022 11094 19068
rect 11150 19022 11202 19068
rect 1760 19019 1812 19022
rect 1868 19019 1920 19022
rect 1976 19019 2028 19022
rect 2084 19019 2136 19022
rect 2192 19019 2244 19022
rect 2300 19019 2352 19022
rect 2408 19019 2460 19022
rect 2516 19019 2568 19022
rect 2624 19019 2676 19022
rect 2732 19019 2784 19022
rect 2840 19019 2892 19022
rect 2948 19019 3000 19022
rect 3056 19019 3108 19022
rect 3164 19019 3216 19022
rect 3272 19019 3324 19022
rect 3380 19019 3432 19022
rect 3488 19019 3540 19022
rect 3596 19019 3648 19022
rect 3704 19019 3756 19022
rect 4130 19019 4182 19022
rect 4238 19019 4290 19022
rect 4346 19019 4398 19022
rect 4454 19019 4506 19022
rect 4562 19019 4614 19022
rect 4670 19019 4722 19022
rect 4778 19019 4830 19022
rect 4886 19019 4938 19022
rect 4994 19019 5046 19022
rect 5102 19019 5154 19022
rect 5210 19019 5262 19022
rect 5318 19019 5370 19022
rect 5426 19019 5478 19022
rect 5534 19019 5586 19022
rect 5642 19019 5694 19022
rect 5750 19019 5802 19022
rect 5858 19019 5910 19022
rect 5966 19019 6018 19022
rect 6074 19019 6126 19022
rect 6836 19019 6888 19022
rect 6944 19019 6996 19022
rect 7052 19019 7104 19022
rect 7160 19019 7212 19022
rect 7268 19019 7320 19022
rect 7376 19019 7428 19022
rect 7484 19019 7536 19022
rect 7592 19019 7644 19022
rect 7700 19019 7752 19022
rect 7808 19019 7860 19022
rect 7916 19019 7968 19022
rect 8024 19019 8076 19022
rect 8132 19019 8184 19022
rect 8240 19019 8292 19022
rect 8348 19019 8400 19022
rect 8456 19019 8508 19022
rect 8564 19019 8616 19022
rect 8672 19019 8724 19022
rect 8780 19019 8832 19022
rect 9206 19019 9258 19022
rect 9314 19019 9366 19022
rect 9422 19019 9474 19022
rect 9530 19019 9582 19022
rect 9638 19019 9690 19022
rect 9746 19019 9798 19022
rect 9854 19019 9906 19022
rect 9962 19019 10014 19022
rect 10070 19019 10122 19022
rect 10178 19019 10230 19022
rect 10286 19019 10338 19022
rect 10394 19019 10446 19022
rect 10502 19019 10554 19022
rect 10610 19019 10662 19022
rect 10718 19019 10770 19022
rect 10826 19019 10878 19022
rect 10934 19019 10986 19022
rect 11042 19019 11094 19022
rect 11150 19019 11202 19022
rect 12051 24315 12103 24367
rect 12159 24315 12211 24367
rect 12267 24315 12319 24367
rect 12051 24207 12103 24259
rect 12159 24207 12211 24259
rect 12267 24207 12319 24259
rect 12051 24099 12103 24151
rect 12159 24099 12211 24151
rect 12267 24099 12319 24151
rect 12051 23991 12103 24043
rect 12159 23991 12211 24043
rect 12267 23991 12319 24043
rect 12051 23883 12103 23935
rect 12159 23883 12211 23935
rect 12267 23883 12319 23935
rect 12051 23775 12103 23827
rect 12159 23775 12211 23827
rect 12267 23775 12319 23827
rect 12051 23667 12103 23719
rect 12159 23667 12211 23719
rect 12267 23667 12319 23719
rect 12051 23559 12103 23611
rect 12159 23559 12211 23611
rect 12267 23559 12319 23611
rect 12051 23451 12103 23503
rect 12159 23451 12211 23503
rect 12267 23451 12319 23503
rect 12051 23343 12103 23395
rect 12159 23343 12211 23395
rect 12267 23343 12319 23395
rect 12051 23235 12103 23287
rect 12159 23235 12211 23287
rect 12267 23235 12319 23287
rect 12051 23127 12103 23179
rect 12159 23127 12211 23179
rect 12267 23127 12319 23179
rect 12051 23019 12103 23071
rect 12159 23019 12211 23071
rect 12267 23019 12319 23071
rect 12051 22911 12103 22963
rect 12159 22911 12211 22963
rect 12267 22911 12319 22963
rect 12051 22803 12103 22855
rect 12159 22803 12211 22855
rect 12267 22803 12319 22855
rect 12051 22695 12103 22747
rect 12159 22695 12211 22747
rect 12267 22695 12319 22747
rect 12051 22587 12103 22639
rect 12159 22587 12211 22639
rect 12267 22587 12319 22639
rect 12051 22479 12103 22531
rect 12159 22479 12211 22531
rect 12267 22479 12319 22531
rect 12051 22371 12103 22423
rect 12159 22371 12211 22423
rect 12267 22371 12319 22423
rect 12051 22263 12103 22315
rect 12159 22263 12211 22315
rect 12267 22263 12319 22315
rect 12051 22155 12103 22207
rect 12159 22155 12211 22207
rect 12267 22155 12319 22207
rect 12051 22047 12103 22099
rect 12159 22047 12211 22099
rect 12267 22047 12319 22099
rect 12051 21939 12103 21991
rect 12159 21939 12211 21991
rect 12267 21939 12319 21991
rect 12051 21831 12103 21883
rect 12159 21831 12211 21883
rect 12267 21831 12319 21883
rect 12051 21723 12103 21775
rect 12159 21723 12211 21775
rect 12267 21723 12319 21775
rect 12051 21615 12103 21667
rect 12159 21615 12211 21667
rect 12267 21615 12319 21667
rect 12051 21507 12103 21559
rect 12159 21507 12211 21559
rect 12267 21507 12319 21559
rect 12051 21399 12103 21451
rect 12159 21399 12211 21451
rect 12267 21399 12319 21451
rect 12051 21291 12103 21343
rect 12159 21291 12211 21343
rect 12267 21291 12319 21343
rect 12051 21183 12103 21235
rect 12159 21183 12211 21235
rect 12267 21183 12319 21235
rect 12051 21075 12103 21127
rect 12159 21075 12211 21127
rect 12267 21075 12319 21127
rect 12051 20967 12103 21019
rect 12159 20967 12211 21019
rect 12267 20967 12319 21019
rect 12051 20859 12103 20911
rect 12159 20859 12211 20911
rect 12267 20859 12319 20911
rect 12051 20751 12103 20803
rect 12159 20751 12211 20803
rect 12267 20751 12319 20803
rect 12051 20643 12103 20695
rect 12159 20643 12211 20695
rect 12267 20643 12319 20695
rect 12051 20535 12103 20587
rect 12159 20535 12211 20587
rect 12267 20535 12319 20587
rect 12051 20427 12103 20479
rect 12159 20427 12211 20479
rect 12267 20427 12319 20479
rect 12051 20319 12103 20371
rect 12159 20319 12211 20371
rect 12267 20319 12319 20371
rect 12051 20211 12103 20263
rect 12159 20211 12211 20263
rect 12267 20211 12319 20263
rect 12051 20103 12103 20155
rect 12159 20103 12211 20155
rect 12267 20103 12319 20155
rect 12051 19995 12103 20047
rect 12159 19995 12211 20047
rect 12267 19995 12319 20047
rect 12051 19887 12103 19939
rect 12159 19887 12211 19939
rect 12267 19887 12319 19939
rect 12051 19779 12103 19831
rect 12159 19779 12211 19831
rect 12267 19779 12319 19831
rect 12051 19671 12103 19723
rect 12159 19671 12211 19723
rect 12267 19671 12319 19723
rect 12051 19563 12103 19615
rect 12159 19563 12211 19615
rect 12267 19563 12319 19615
rect 12051 19455 12103 19507
rect 12159 19455 12211 19507
rect 12267 19455 12319 19507
rect 12051 19347 12103 19399
rect 12159 19347 12211 19399
rect 12267 19347 12319 19399
rect 12051 19239 12103 19291
rect 12159 19239 12211 19291
rect 12267 19239 12319 19291
rect 12051 19131 12103 19183
rect 12159 19131 12211 19183
rect 12267 19131 12319 19183
rect 12051 19023 12103 19075
rect 12159 19023 12211 19075
rect 12267 19023 12319 19075
rect 12051 18915 12103 18967
rect 12159 18915 12211 18967
rect 12267 18915 12319 18967
rect 12051 18807 12103 18859
rect 12159 18807 12211 18859
rect 12267 18807 12319 18859
rect 12051 18699 12103 18751
rect 12159 18699 12211 18751
rect 12267 18699 12319 18751
rect 1760 18622 1812 18629
rect 1868 18622 1920 18629
rect 1976 18622 2028 18629
rect 2084 18622 2136 18629
rect 2192 18622 2244 18629
rect 2300 18622 2352 18629
rect 2408 18622 2460 18629
rect 2516 18622 2568 18629
rect 2624 18622 2676 18629
rect 2732 18622 2784 18629
rect 2840 18622 2892 18629
rect 2948 18622 3000 18629
rect 3056 18622 3108 18629
rect 3164 18622 3216 18629
rect 3272 18622 3324 18629
rect 3380 18622 3432 18629
rect 3488 18622 3540 18629
rect 3596 18622 3648 18629
rect 3704 18622 3756 18629
rect 4130 18622 4182 18629
rect 4238 18622 4290 18629
rect 4346 18622 4398 18629
rect 4454 18622 4506 18629
rect 4562 18622 4614 18629
rect 4670 18622 4722 18629
rect 4778 18622 4830 18629
rect 4886 18622 4938 18629
rect 4994 18622 5046 18629
rect 5102 18622 5154 18629
rect 5210 18622 5262 18629
rect 5318 18622 5370 18629
rect 5426 18622 5478 18629
rect 5534 18622 5586 18629
rect 5642 18622 5694 18629
rect 5750 18622 5802 18629
rect 5858 18622 5910 18629
rect 5966 18622 6018 18629
rect 6074 18622 6126 18629
rect 6836 18622 6888 18629
rect 6944 18622 6996 18629
rect 7052 18622 7104 18629
rect 7160 18622 7212 18629
rect 7268 18622 7320 18629
rect 7376 18622 7428 18629
rect 7484 18622 7536 18629
rect 7592 18622 7644 18629
rect 7700 18622 7752 18629
rect 7808 18622 7860 18629
rect 7916 18622 7968 18629
rect 8024 18622 8076 18629
rect 8132 18622 8184 18629
rect 8240 18622 8292 18629
rect 8348 18622 8400 18629
rect 8456 18622 8508 18629
rect 8564 18622 8616 18629
rect 8672 18622 8724 18629
rect 8780 18622 8832 18629
rect 9206 18622 9258 18629
rect 9314 18622 9366 18629
rect 9422 18622 9474 18629
rect 9530 18622 9582 18629
rect 9638 18622 9690 18629
rect 9746 18622 9798 18629
rect 9854 18622 9906 18629
rect 9962 18622 10014 18629
rect 10070 18622 10122 18629
rect 10178 18622 10230 18629
rect 10286 18622 10338 18629
rect 10394 18622 10446 18629
rect 10502 18622 10554 18629
rect 10610 18622 10662 18629
rect 10718 18622 10770 18629
rect 10826 18622 10878 18629
rect 10934 18622 10986 18629
rect 11042 18622 11094 18629
rect 11150 18622 11202 18629
rect 643 18483 695 18535
rect 751 18483 803 18535
rect 859 18483 911 18535
rect 1760 18577 1812 18622
rect 1868 18577 1920 18622
rect 1976 18577 2028 18622
rect 2084 18577 2136 18622
rect 2192 18577 2244 18622
rect 2300 18577 2352 18622
rect 2408 18577 2460 18622
rect 2516 18577 2568 18622
rect 2624 18577 2676 18622
rect 2732 18577 2784 18622
rect 2840 18577 2892 18622
rect 2948 18577 3000 18622
rect 3056 18577 3108 18622
rect 3164 18577 3216 18622
rect 3272 18577 3324 18622
rect 3380 18577 3432 18622
rect 3488 18577 3540 18622
rect 3596 18577 3648 18622
rect 3704 18577 3756 18622
rect 4130 18577 4182 18622
rect 4238 18577 4290 18622
rect 4346 18577 4398 18622
rect 4454 18577 4506 18622
rect 4562 18577 4614 18622
rect 4670 18577 4722 18622
rect 4778 18577 4830 18622
rect 4886 18577 4938 18622
rect 4994 18577 5046 18622
rect 5102 18577 5154 18622
rect 5210 18577 5262 18622
rect 5318 18577 5370 18622
rect 5426 18577 5478 18622
rect 5534 18577 5586 18622
rect 5642 18577 5694 18622
rect 5750 18577 5802 18622
rect 5858 18577 5910 18622
rect 5966 18577 6018 18622
rect 6074 18577 6126 18622
rect 6836 18577 6888 18622
rect 6944 18577 6996 18622
rect 7052 18577 7104 18622
rect 7160 18577 7212 18622
rect 7268 18577 7320 18622
rect 7376 18577 7428 18622
rect 7484 18577 7536 18622
rect 7592 18577 7644 18622
rect 7700 18577 7752 18622
rect 7808 18577 7860 18622
rect 7916 18577 7968 18622
rect 8024 18577 8076 18622
rect 8132 18577 8184 18622
rect 8240 18577 8292 18622
rect 8348 18577 8400 18622
rect 8456 18577 8508 18622
rect 8564 18577 8616 18622
rect 8672 18577 8724 18622
rect 8780 18577 8832 18622
rect 9206 18577 9258 18622
rect 9314 18577 9366 18622
rect 9422 18577 9474 18622
rect 9530 18577 9582 18622
rect 9638 18577 9690 18622
rect 9746 18577 9798 18622
rect 9854 18577 9906 18622
rect 9962 18577 10014 18622
rect 10070 18577 10122 18622
rect 10178 18577 10230 18622
rect 10286 18577 10338 18622
rect 10394 18577 10446 18622
rect 10502 18577 10554 18622
rect 10610 18577 10662 18622
rect 10718 18577 10770 18622
rect 10826 18577 10878 18622
rect 10934 18577 10986 18622
rect 11042 18577 11094 18622
rect 11150 18577 11202 18622
rect 1760 18476 1812 18521
rect 1868 18476 1920 18521
rect 1976 18476 2028 18521
rect 2084 18476 2136 18521
rect 2192 18476 2244 18521
rect 2300 18476 2352 18521
rect 2408 18476 2460 18521
rect 2516 18476 2568 18521
rect 2624 18476 2676 18521
rect 2732 18476 2784 18521
rect 2840 18476 2892 18521
rect 2948 18476 3000 18521
rect 3056 18476 3108 18521
rect 3164 18476 3216 18521
rect 3272 18476 3324 18521
rect 3380 18476 3432 18521
rect 3488 18476 3540 18521
rect 3596 18476 3648 18521
rect 3704 18476 3756 18521
rect 4130 18476 4182 18521
rect 4238 18476 4290 18521
rect 4346 18476 4398 18521
rect 4454 18476 4506 18521
rect 4562 18476 4614 18521
rect 4670 18476 4722 18521
rect 4778 18476 4830 18521
rect 4886 18476 4938 18521
rect 4994 18476 5046 18521
rect 5102 18476 5154 18521
rect 5210 18476 5262 18521
rect 5318 18476 5370 18521
rect 5426 18476 5478 18521
rect 5534 18476 5586 18521
rect 5642 18476 5694 18521
rect 5750 18476 5802 18521
rect 5858 18476 5910 18521
rect 5966 18476 6018 18521
rect 6074 18476 6126 18521
rect 6836 18476 6888 18521
rect 6944 18476 6996 18521
rect 7052 18476 7104 18521
rect 7160 18476 7212 18521
rect 7268 18476 7320 18521
rect 7376 18476 7428 18521
rect 7484 18476 7536 18521
rect 7592 18476 7644 18521
rect 7700 18476 7752 18521
rect 7808 18476 7860 18521
rect 7916 18476 7968 18521
rect 8024 18476 8076 18521
rect 8132 18476 8184 18521
rect 8240 18476 8292 18521
rect 8348 18476 8400 18521
rect 8456 18476 8508 18521
rect 8564 18476 8616 18521
rect 8672 18476 8724 18521
rect 8780 18476 8832 18521
rect 9206 18476 9258 18521
rect 9314 18476 9366 18521
rect 9422 18476 9474 18521
rect 9530 18476 9582 18521
rect 9638 18476 9690 18521
rect 9746 18476 9798 18521
rect 9854 18476 9906 18521
rect 9962 18476 10014 18521
rect 10070 18476 10122 18521
rect 10178 18476 10230 18521
rect 10286 18476 10338 18521
rect 10394 18476 10446 18521
rect 10502 18476 10554 18521
rect 10610 18476 10662 18521
rect 10718 18476 10770 18521
rect 10826 18476 10878 18521
rect 10934 18476 10986 18521
rect 11042 18476 11094 18521
rect 11150 18476 11202 18521
rect 12051 18591 12103 18643
rect 12159 18591 12211 18643
rect 12267 18591 12319 18643
rect 12051 18483 12103 18535
rect 12159 18483 12211 18535
rect 12267 18483 12319 18535
rect 1760 18469 1812 18476
rect 1868 18469 1920 18476
rect 1976 18469 2028 18476
rect 2084 18469 2136 18476
rect 2192 18469 2244 18476
rect 2300 18469 2352 18476
rect 2408 18469 2460 18476
rect 2516 18469 2568 18476
rect 2624 18469 2676 18476
rect 2732 18469 2784 18476
rect 2840 18469 2892 18476
rect 2948 18469 3000 18476
rect 3056 18469 3108 18476
rect 3164 18469 3216 18476
rect 3272 18469 3324 18476
rect 3380 18469 3432 18476
rect 3488 18469 3540 18476
rect 3596 18469 3648 18476
rect 3704 18469 3756 18476
rect 4130 18469 4182 18476
rect 4238 18469 4290 18476
rect 4346 18469 4398 18476
rect 4454 18469 4506 18476
rect 4562 18469 4614 18476
rect 4670 18469 4722 18476
rect 4778 18469 4830 18476
rect 4886 18469 4938 18476
rect 4994 18469 5046 18476
rect 5102 18469 5154 18476
rect 5210 18469 5262 18476
rect 5318 18469 5370 18476
rect 5426 18469 5478 18476
rect 5534 18469 5586 18476
rect 5642 18469 5694 18476
rect 5750 18469 5802 18476
rect 5858 18469 5910 18476
rect 5966 18469 6018 18476
rect 6074 18469 6126 18476
rect 6836 18469 6888 18476
rect 6944 18469 6996 18476
rect 7052 18469 7104 18476
rect 7160 18469 7212 18476
rect 7268 18469 7320 18476
rect 7376 18469 7428 18476
rect 7484 18469 7536 18476
rect 7592 18469 7644 18476
rect 7700 18469 7752 18476
rect 7808 18469 7860 18476
rect 7916 18469 7968 18476
rect 8024 18469 8076 18476
rect 8132 18469 8184 18476
rect 8240 18469 8292 18476
rect 8348 18469 8400 18476
rect 8456 18469 8508 18476
rect 8564 18469 8616 18476
rect 8672 18469 8724 18476
rect 8780 18469 8832 18476
rect 9206 18469 9258 18476
rect 9314 18469 9366 18476
rect 9422 18469 9474 18476
rect 9530 18469 9582 18476
rect 9638 18469 9690 18476
rect 9746 18469 9798 18476
rect 9854 18469 9906 18476
rect 9962 18469 10014 18476
rect 10070 18469 10122 18476
rect 10178 18469 10230 18476
rect 10286 18469 10338 18476
rect 10394 18469 10446 18476
rect 10502 18469 10554 18476
rect 10610 18469 10662 18476
rect 10718 18469 10770 18476
rect 10826 18469 10878 18476
rect 10934 18469 10986 18476
rect 11042 18469 11094 18476
rect 11150 18469 11202 18476
rect 643 18375 695 18427
rect 751 18375 803 18427
rect 859 18375 911 18427
rect 643 18267 695 18319
rect 751 18267 803 18319
rect 859 18267 911 18319
rect 643 18159 695 18211
rect 751 18159 803 18211
rect 859 18159 911 18211
rect 643 18051 695 18103
rect 751 18051 803 18103
rect 859 18051 911 18103
rect 643 17943 695 17995
rect 751 17943 803 17995
rect 859 17943 911 17995
rect 643 17835 695 17887
rect 751 17835 803 17887
rect 859 17835 911 17887
rect 643 17727 695 17779
rect 751 17727 803 17779
rect 859 17727 911 17779
rect 643 17619 695 17671
rect 751 17619 803 17671
rect 859 17619 911 17671
rect 643 17511 695 17563
rect 751 17511 803 17563
rect 859 17511 911 17563
rect 643 17403 695 17455
rect 751 17403 803 17455
rect 859 17403 911 17455
rect 643 17295 695 17347
rect 751 17295 803 17347
rect 859 17295 911 17347
rect 643 17187 695 17239
rect 751 17187 803 17239
rect 859 17187 911 17239
rect 643 17079 695 17131
rect 751 17079 803 17131
rect 859 17079 911 17131
rect 643 16971 695 17023
rect 751 16971 803 17023
rect 859 16971 911 17023
rect 643 16863 695 16915
rect 751 16863 803 16915
rect 859 16863 911 16915
rect 643 16755 695 16807
rect 751 16755 803 16807
rect 859 16755 911 16807
rect 643 16647 695 16699
rect 751 16647 803 16699
rect 859 16647 911 16699
rect 643 16539 695 16591
rect 751 16539 803 16591
rect 859 16539 911 16591
rect 643 16431 695 16483
rect 751 16431 803 16483
rect 859 16431 911 16483
rect 643 16323 695 16375
rect 751 16323 803 16375
rect 859 16323 911 16375
rect 643 16215 695 16267
rect 751 16215 803 16267
rect 859 16215 911 16267
rect 643 16107 695 16159
rect 751 16107 803 16159
rect 859 16107 911 16159
rect 643 15999 695 16051
rect 751 15999 803 16051
rect 859 15999 911 16051
rect 643 15891 695 15943
rect 751 15891 803 15943
rect 859 15891 911 15943
rect 643 15783 695 15835
rect 751 15783 803 15835
rect 859 15783 911 15835
rect 643 15675 695 15727
rect 751 15675 803 15727
rect 859 15675 911 15727
rect 643 15567 695 15619
rect 751 15567 803 15619
rect 859 15567 911 15619
rect 643 15459 695 15511
rect 751 15459 803 15511
rect 859 15459 911 15511
rect 643 15351 695 15403
rect 751 15351 803 15403
rect 859 15351 911 15403
rect 643 15243 695 15295
rect 751 15243 803 15295
rect 859 15243 911 15295
rect 643 15135 695 15187
rect 751 15135 803 15187
rect 859 15135 911 15187
rect 643 15027 695 15079
rect 751 15027 803 15079
rect 859 15027 911 15079
rect 643 14919 695 14971
rect 751 14919 803 14971
rect 859 14919 911 14971
rect 643 14811 695 14863
rect 751 14811 803 14863
rect 859 14811 911 14863
rect 643 14703 695 14755
rect 751 14703 803 14755
rect 859 14703 911 14755
rect 643 14595 695 14647
rect 751 14595 803 14647
rect 859 14595 911 14647
rect 643 14487 695 14539
rect 751 14487 803 14539
rect 859 14487 911 14539
rect 643 14379 695 14431
rect 751 14379 803 14431
rect 859 14379 911 14431
rect 643 14271 695 14323
rect 751 14271 803 14323
rect 859 14271 911 14323
rect 643 14163 695 14215
rect 751 14163 803 14215
rect 859 14163 911 14215
rect 643 14055 695 14107
rect 751 14055 803 14107
rect 859 14055 911 14107
rect 643 13947 695 13999
rect 751 13947 803 13999
rect 859 13947 911 13999
rect 643 13839 695 13891
rect 751 13839 803 13891
rect 859 13839 911 13891
rect 643 13731 695 13783
rect 751 13731 803 13783
rect 859 13731 911 13783
rect 643 13623 695 13675
rect 751 13623 803 13675
rect 859 13623 911 13675
rect 643 13515 695 13567
rect 751 13515 803 13567
rect 859 13515 911 13567
rect 643 13407 695 13459
rect 751 13407 803 13459
rect 859 13407 911 13459
rect 643 13299 695 13351
rect 751 13299 803 13351
rect 859 13299 911 13351
rect 643 13191 695 13243
rect 751 13191 803 13243
rect 859 13191 911 13243
rect 643 13083 695 13135
rect 751 13083 803 13135
rect 859 13083 911 13135
rect 643 12975 695 13027
rect 751 12975 803 13027
rect 859 12975 911 13027
rect 643 12867 695 12919
rect 751 12867 803 12919
rect 859 12867 911 12919
rect 643 12759 695 12811
rect 751 12759 803 12811
rect 859 12759 911 12811
rect 1760 18076 1812 18079
rect 1868 18076 1920 18079
rect 1976 18076 2028 18079
rect 2084 18076 2136 18079
rect 2192 18076 2244 18079
rect 2300 18076 2352 18079
rect 2408 18076 2460 18079
rect 2516 18076 2568 18079
rect 2624 18076 2676 18079
rect 2732 18076 2784 18079
rect 2840 18076 2892 18079
rect 2948 18076 3000 18079
rect 3056 18076 3108 18079
rect 3164 18076 3216 18079
rect 3272 18076 3324 18079
rect 3380 18076 3432 18079
rect 3488 18076 3540 18079
rect 3596 18076 3648 18079
rect 3704 18076 3756 18079
rect 4130 18076 4182 18079
rect 4238 18076 4290 18079
rect 4346 18076 4398 18079
rect 4454 18076 4506 18079
rect 4562 18076 4614 18079
rect 4670 18076 4722 18079
rect 4778 18076 4830 18079
rect 4886 18076 4938 18079
rect 4994 18076 5046 18079
rect 5102 18076 5154 18079
rect 5210 18076 5262 18079
rect 5318 18076 5370 18079
rect 5426 18076 5478 18079
rect 5534 18076 5586 18079
rect 5642 18076 5694 18079
rect 5750 18076 5802 18079
rect 5858 18076 5910 18079
rect 5966 18076 6018 18079
rect 6074 18076 6126 18079
rect 6836 18076 6888 18079
rect 6944 18076 6996 18079
rect 7052 18076 7104 18079
rect 7160 18076 7212 18079
rect 7268 18076 7320 18079
rect 7376 18076 7428 18079
rect 7484 18076 7536 18079
rect 7592 18076 7644 18079
rect 7700 18076 7752 18079
rect 7808 18076 7860 18079
rect 7916 18076 7968 18079
rect 8024 18076 8076 18079
rect 8132 18076 8184 18079
rect 8240 18076 8292 18079
rect 8348 18076 8400 18079
rect 8456 18076 8508 18079
rect 8564 18076 8616 18079
rect 8672 18076 8724 18079
rect 8780 18076 8832 18079
rect 9206 18076 9258 18079
rect 9314 18076 9366 18079
rect 9422 18076 9474 18079
rect 9530 18076 9582 18079
rect 9638 18076 9690 18079
rect 9746 18076 9798 18079
rect 9854 18076 9906 18079
rect 9962 18076 10014 18079
rect 10070 18076 10122 18079
rect 10178 18076 10230 18079
rect 10286 18076 10338 18079
rect 10394 18076 10446 18079
rect 10502 18076 10554 18079
rect 10610 18076 10662 18079
rect 10718 18076 10770 18079
rect 10826 18076 10878 18079
rect 10934 18076 10986 18079
rect 11042 18076 11094 18079
rect 11150 18076 11202 18079
rect 1760 18030 1812 18076
rect 1868 18030 1920 18076
rect 1976 18030 2028 18076
rect 2084 18030 2136 18076
rect 2192 18030 2244 18076
rect 2300 18030 2352 18076
rect 2408 18030 2460 18076
rect 2516 18030 2568 18076
rect 2624 18030 2676 18076
rect 2732 18030 2784 18076
rect 2840 18030 2892 18076
rect 2948 18030 3000 18076
rect 3056 18030 3108 18076
rect 3164 18030 3216 18076
rect 3272 18030 3324 18076
rect 3380 18030 3432 18076
rect 3488 18030 3540 18076
rect 3596 18030 3648 18076
rect 3704 18030 3756 18076
rect 4130 18030 4182 18076
rect 4238 18030 4290 18076
rect 4346 18030 4398 18076
rect 4454 18030 4506 18076
rect 4562 18030 4614 18076
rect 4670 18030 4722 18076
rect 4778 18030 4830 18076
rect 4886 18030 4938 18076
rect 4994 18030 5046 18076
rect 5102 18030 5154 18076
rect 5210 18030 5262 18076
rect 5318 18030 5370 18076
rect 5426 18030 5478 18076
rect 5534 18030 5586 18076
rect 5642 18030 5694 18076
rect 5750 18030 5802 18076
rect 5858 18030 5910 18076
rect 5966 18030 6018 18076
rect 6074 18030 6126 18076
rect 6836 18030 6888 18076
rect 6944 18030 6996 18076
rect 7052 18030 7104 18076
rect 7160 18030 7212 18076
rect 7268 18030 7320 18076
rect 7376 18030 7428 18076
rect 7484 18030 7536 18076
rect 7592 18030 7644 18076
rect 7700 18030 7752 18076
rect 7808 18030 7860 18076
rect 7916 18030 7968 18076
rect 8024 18030 8076 18076
rect 8132 18030 8184 18076
rect 8240 18030 8292 18076
rect 8348 18030 8400 18076
rect 8456 18030 8508 18076
rect 8564 18030 8616 18076
rect 8672 18030 8724 18076
rect 8780 18030 8832 18076
rect 9206 18030 9258 18076
rect 9314 18030 9366 18076
rect 9422 18030 9474 18076
rect 9530 18030 9582 18076
rect 9638 18030 9690 18076
rect 9746 18030 9798 18076
rect 9854 18030 9906 18076
rect 9962 18030 10014 18076
rect 10070 18030 10122 18076
rect 10178 18030 10230 18076
rect 10286 18030 10338 18076
rect 10394 18030 10446 18076
rect 10502 18030 10554 18076
rect 10610 18030 10662 18076
rect 10718 18030 10770 18076
rect 10826 18030 10878 18076
rect 10934 18030 10986 18076
rect 11042 18030 11094 18076
rect 11150 18030 11202 18076
rect 1760 18027 1812 18030
rect 1868 18027 1920 18030
rect 1976 18027 2028 18030
rect 2084 18027 2136 18030
rect 2192 18027 2244 18030
rect 2300 18027 2352 18030
rect 2408 18027 2460 18030
rect 2516 18027 2568 18030
rect 2624 18027 2676 18030
rect 2732 18027 2784 18030
rect 2840 18027 2892 18030
rect 2948 18027 3000 18030
rect 3056 18027 3108 18030
rect 3164 18027 3216 18030
rect 3272 18027 3324 18030
rect 3380 18027 3432 18030
rect 3488 18027 3540 18030
rect 3596 18027 3648 18030
rect 3704 18027 3756 18030
rect 4130 18027 4182 18030
rect 4238 18027 4290 18030
rect 4346 18027 4398 18030
rect 4454 18027 4506 18030
rect 4562 18027 4614 18030
rect 4670 18027 4722 18030
rect 4778 18027 4830 18030
rect 4886 18027 4938 18030
rect 4994 18027 5046 18030
rect 5102 18027 5154 18030
rect 5210 18027 5262 18030
rect 5318 18027 5370 18030
rect 5426 18027 5478 18030
rect 5534 18027 5586 18030
rect 5642 18027 5694 18030
rect 5750 18027 5802 18030
rect 5858 18027 5910 18030
rect 5966 18027 6018 18030
rect 6074 18027 6126 18030
rect 6836 18027 6888 18030
rect 6944 18027 6996 18030
rect 7052 18027 7104 18030
rect 7160 18027 7212 18030
rect 7268 18027 7320 18030
rect 7376 18027 7428 18030
rect 7484 18027 7536 18030
rect 7592 18027 7644 18030
rect 7700 18027 7752 18030
rect 7808 18027 7860 18030
rect 7916 18027 7968 18030
rect 8024 18027 8076 18030
rect 8132 18027 8184 18030
rect 8240 18027 8292 18030
rect 8348 18027 8400 18030
rect 8456 18027 8508 18030
rect 8564 18027 8616 18030
rect 8672 18027 8724 18030
rect 8780 18027 8832 18030
rect 9206 18027 9258 18030
rect 9314 18027 9366 18030
rect 9422 18027 9474 18030
rect 9530 18027 9582 18030
rect 9638 18027 9690 18030
rect 9746 18027 9798 18030
rect 9854 18027 9906 18030
rect 9962 18027 10014 18030
rect 10070 18027 10122 18030
rect 10178 18027 10230 18030
rect 10286 18027 10338 18030
rect 10394 18027 10446 18030
rect 10502 18027 10554 18030
rect 10610 18027 10662 18030
rect 10718 18027 10770 18030
rect 10826 18027 10878 18030
rect 10934 18027 10986 18030
rect 11042 18027 11094 18030
rect 11150 18027 11202 18030
rect 1233 17963 1285 18015
rect 1341 17963 1393 18015
rect 1233 17855 1256 17907
rect 1256 17855 1285 17907
rect 1341 17855 1393 17907
rect 1233 17747 1256 17799
rect 1256 17747 1285 17799
rect 1341 17747 1393 17799
rect 1233 17639 1256 17691
rect 1256 17639 1285 17691
rect 1341 17639 1393 17691
rect 1233 17531 1256 17583
rect 1256 17531 1285 17583
rect 1341 17531 1393 17583
rect 1233 17423 1256 17475
rect 1256 17423 1285 17475
rect 1341 17423 1393 17475
rect 1233 17315 1256 17367
rect 1256 17315 1285 17367
rect 1341 17315 1393 17367
rect 1233 17207 1256 17259
rect 1256 17207 1285 17259
rect 1341 17207 1393 17259
rect 1233 17099 1256 17151
rect 1256 17099 1285 17151
rect 1341 17099 1393 17151
rect 1233 16991 1256 17043
rect 1256 16991 1285 17043
rect 1341 16991 1393 17043
rect 1233 16883 1256 16935
rect 1256 16883 1285 16935
rect 1341 16883 1393 16935
rect 1233 16775 1256 16827
rect 1256 16775 1285 16827
rect 1341 16775 1393 16827
rect 1233 16667 1256 16719
rect 1256 16667 1285 16719
rect 1341 16667 1393 16719
rect 1233 16559 1256 16611
rect 1256 16559 1285 16611
rect 1341 16559 1393 16611
rect 1233 16451 1256 16503
rect 1256 16451 1285 16503
rect 1341 16451 1393 16503
rect 1233 16343 1256 16395
rect 1256 16343 1285 16395
rect 1341 16343 1393 16395
rect 1233 16235 1256 16287
rect 1256 16235 1285 16287
rect 1341 16235 1393 16287
rect 1233 16127 1256 16179
rect 1256 16127 1285 16179
rect 1341 16127 1393 16179
rect 1233 16019 1256 16071
rect 1256 16019 1285 16071
rect 1341 16019 1393 16071
rect 1233 15911 1256 15963
rect 1256 15911 1285 15963
rect 1341 15911 1393 15963
rect 1233 15803 1256 15855
rect 1256 15803 1285 15855
rect 1341 15803 1393 15855
rect 1233 15695 1256 15747
rect 1256 15695 1285 15747
rect 1341 15695 1393 15747
rect 1233 15587 1256 15639
rect 1256 15587 1285 15639
rect 1341 15587 1393 15639
rect 1233 15479 1256 15531
rect 1256 15479 1285 15531
rect 1341 15479 1393 15531
rect 1233 15371 1256 15423
rect 1256 15371 1285 15423
rect 1341 15371 1393 15423
rect 1233 15263 1256 15315
rect 1256 15263 1285 15315
rect 1341 15263 1393 15315
rect 1233 15155 1256 15207
rect 1256 15155 1285 15207
rect 1341 15155 1393 15207
rect 1233 15047 1256 15099
rect 1256 15047 1285 15099
rect 1341 15047 1393 15099
rect 1233 14939 1256 14991
rect 1256 14939 1285 14991
rect 1341 14939 1393 14991
rect 1233 14831 1256 14883
rect 1256 14831 1285 14883
rect 1341 14831 1393 14883
rect 1233 14723 1256 14775
rect 1256 14723 1285 14775
rect 1341 14723 1393 14775
rect 1233 14615 1256 14667
rect 1256 14615 1285 14667
rect 1341 14615 1393 14667
rect 1233 14507 1256 14559
rect 1256 14507 1285 14559
rect 1341 14507 1393 14559
rect 1233 14399 1256 14451
rect 1256 14399 1285 14451
rect 1341 14399 1393 14451
rect 1233 14291 1256 14343
rect 1256 14291 1285 14343
rect 1341 14291 1393 14343
rect 1233 14183 1256 14235
rect 1256 14183 1285 14235
rect 1341 14183 1393 14235
rect 1233 14075 1256 14127
rect 1256 14075 1285 14127
rect 1341 14075 1393 14127
rect 1233 13967 1256 14019
rect 1256 13967 1285 14019
rect 1341 13967 1393 14019
rect 1233 13859 1256 13911
rect 1256 13859 1285 13911
rect 1341 13859 1393 13911
rect 1233 13751 1256 13803
rect 1256 13751 1285 13803
rect 1341 13751 1393 13803
rect 1233 13643 1256 13695
rect 1256 13643 1285 13695
rect 1341 13643 1393 13695
rect 1233 13535 1256 13587
rect 1256 13535 1285 13587
rect 1341 13535 1393 13587
rect 1233 13427 1256 13479
rect 1256 13427 1285 13479
rect 1341 13427 1393 13479
rect 1233 13319 1256 13371
rect 1256 13319 1285 13371
rect 1341 13319 1393 13371
rect 11569 17963 11621 18015
rect 11677 17963 11729 18015
rect 1493 17832 1545 17835
rect 1601 17832 1653 17835
rect 3863 17832 3915 17835
rect 3971 17832 4023 17835
rect 6239 17832 6291 17835
rect 6347 17832 6399 17835
rect 6455 17832 6507 17835
rect 6563 17832 6615 17835
rect 6671 17832 6723 17835
rect 8939 17832 8991 17835
rect 9047 17832 9099 17835
rect 11309 17832 11361 17835
rect 11417 17832 11469 17835
rect 1493 17786 1494 17832
rect 1494 17786 1545 17832
rect 1601 17786 1653 17832
rect 3863 17786 3915 17832
rect 3971 17786 4023 17832
rect 6239 17786 6291 17832
rect 6347 17786 6399 17832
rect 6455 17786 6507 17832
rect 6563 17786 6615 17832
rect 6671 17786 6723 17832
rect 8939 17786 8991 17832
rect 9047 17786 9099 17832
rect 11309 17786 11361 17832
rect 11417 17786 11468 17832
rect 11468 17786 11469 17832
rect 1493 17783 1545 17786
rect 1601 17783 1653 17786
rect 3863 17783 3915 17786
rect 3971 17783 4023 17786
rect 6239 17783 6291 17786
rect 6347 17783 6399 17786
rect 6455 17783 6507 17786
rect 6563 17783 6615 17786
rect 6671 17783 6723 17786
rect 8939 17783 8991 17786
rect 9047 17783 9099 17786
rect 11309 17783 11361 17786
rect 11417 17783 11469 17786
rect 1760 17588 1812 17591
rect 1868 17588 1920 17591
rect 1976 17588 2028 17591
rect 2084 17588 2136 17591
rect 2192 17588 2244 17591
rect 2300 17588 2352 17591
rect 2408 17588 2460 17591
rect 2516 17588 2568 17591
rect 2624 17588 2676 17591
rect 2732 17588 2784 17591
rect 2840 17588 2892 17591
rect 2948 17588 3000 17591
rect 3056 17588 3108 17591
rect 3164 17588 3216 17591
rect 3272 17588 3324 17591
rect 3380 17588 3432 17591
rect 3488 17588 3540 17591
rect 3596 17588 3648 17591
rect 3704 17588 3756 17591
rect 4130 17588 4182 17591
rect 4238 17588 4290 17591
rect 4346 17588 4398 17591
rect 4454 17588 4506 17591
rect 4562 17588 4614 17591
rect 4670 17588 4722 17591
rect 4778 17588 4830 17591
rect 4886 17588 4938 17591
rect 4994 17588 5046 17591
rect 5102 17588 5154 17591
rect 5210 17588 5262 17591
rect 5318 17588 5370 17591
rect 5426 17588 5478 17591
rect 5534 17588 5586 17591
rect 5642 17588 5694 17591
rect 5750 17588 5802 17591
rect 5858 17588 5910 17591
rect 5966 17588 6018 17591
rect 6074 17588 6126 17591
rect 6836 17588 6888 17591
rect 6944 17588 6996 17591
rect 7052 17588 7104 17591
rect 7160 17588 7212 17591
rect 7268 17588 7320 17591
rect 7376 17588 7428 17591
rect 7484 17588 7536 17591
rect 7592 17588 7644 17591
rect 7700 17588 7752 17591
rect 7808 17588 7860 17591
rect 7916 17588 7968 17591
rect 8024 17588 8076 17591
rect 8132 17588 8184 17591
rect 8240 17588 8292 17591
rect 8348 17588 8400 17591
rect 8456 17588 8508 17591
rect 8564 17588 8616 17591
rect 8672 17588 8724 17591
rect 8780 17588 8832 17591
rect 9206 17588 9258 17591
rect 9314 17588 9366 17591
rect 9422 17588 9474 17591
rect 9530 17588 9582 17591
rect 9638 17588 9690 17591
rect 9746 17588 9798 17591
rect 9854 17588 9906 17591
rect 9962 17588 10014 17591
rect 10070 17588 10122 17591
rect 10178 17588 10230 17591
rect 10286 17588 10338 17591
rect 10394 17588 10446 17591
rect 10502 17588 10554 17591
rect 10610 17588 10662 17591
rect 10718 17588 10770 17591
rect 10826 17588 10878 17591
rect 10934 17588 10986 17591
rect 11042 17588 11094 17591
rect 11150 17588 11202 17591
rect 1760 17542 1812 17588
rect 1868 17542 1920 17588
rect 1976 17542 2028 17588
rect 2084 17542 2136 17588
rect 2192 17542 2244 17588
rect 2300 17542 2352 17588
rect 2408 17542 2460 17588
rect 2516 17542 2568 17588
rect 2624 17542 2676 17588
rect 2732 17542 2784 17588
rect 2840 17542 2892 17588
rect 2948 17542 3000 17588
rect 3056 17542 3108 17588
rect 3164 17542 3216 17588
rect 3272 17542 3324 17588
rect 3380 17542 3432 17588
rect 3488 17542 3540 17588
rect 3596 17542 3648 17588
rect 3704 17542 3756 17588
rect 4130 17542 4182 17588
rect 4238 17542 4290 17588
rect 4346 17542 4398 17588
rect 4454 17542 4506 17588
rect 4562 17542 4614 17588
rect 4670 17542 4722 17588
rect 4778 17542 4830 17588
rect 4886 17542 4938 17588
rect 4994 17542 5046 17588
rect 5102 17542 5154 17588
rect 5210 17542 5262 17588
rect 5318 17542 5370 17588
rect 5426 17542 5478 17588
rect 5534 17542 5586 17588
rect 5642 17542 5694 17588
rect 5750 17542 5802 17588
rect 5858 17542 5910 17588
rect 5966 17542 6018 17588
rect 6074 17542 6126 17588
rect 6836 17542 6888 17588
rect 6944 17542 6996 17588
rect 7052 17542 7104 17588
rect 7160 17542 7212 17588
rect 7268 17542 7320 17588
rect 7376 17542 7428 17588
rect 7484 17542 7536 17588
rect 7592 17542 7644 17588
rect 7700 17542 7752 17588
rect 7808 17542 7860 17588
rect 7916 17542 7968 17588
rect 8024 17542 8076 17588
rect 8132 17542 8184 17588
rect 8240 17542 8292 17588
rect 8348 17542 8400 17588
rect 8456 17542 8508 17588
rect 8564 17542 8616 17588
rect 8672 17542 8724 17588
rect 8780 17542 8832 17588
rect 9206 17542 9258 17588
rect 9314 17542 9366 17588
rect 9422 17542 9474 17588
rect 9530 17542 9582 17588
rect 9638 17542 9690 17588
rect 9746 17542 9798 17588
rect 9854 17542 9906 17588
rect 9962 17542 10014 17588
rect 10070 17542 10122 17588
rect 10178 17542 10230 17588
rect 10286 17542 10338 17588
rect 10394 17542 10446 17588
rect 10502 17542 10554 17588
rect 10610 17542 10662 17588
rect 10718 17542 10770 17588
rect 10826 17542 10878 17588
rect 10934 17542 10986 17588
rect 11042 17542 11094 17588
rect 11150 17542 11202 17588
rect 1760 17539 1812 17542
rect 1868 17539 1920 17542
rect 1976 17539 2028 17542
rect 2084 17539 2136 17542
rect 2192 17539 2244 17542
rect 2300 17539 2352 17542
rect 2408 17539 2460 17542
rect 2516 17539 2568 17542
rect 2624 17539 2676 17542
rect 2732 17539 2784 17542
rect 2840 17539 2892 17542
rect 2948 17539 3000 17542
rect 3056 17539 3108 17542
rect 3164 17539 3216 17542
rect 3272 17539 3324 17542
rect 3380 17539 3432 17542
rect 3488 17539 3540 17542
rect 3596 17539 3648 17542
rect 3704 17539 3756 17542
rect 4130 17539 4182 17542
rect 4238 17539 4290 17542
rect 4346 17539 4398 17542
rect 4454 17539 4506 17542
rect 4562 17539 4614 17542
rect 4670 17539 4722 17542
rect 4778 17539 4830 17542
rect 4886 17539 4938 17542
rect 4994 17539 5046 17542
rect 5102 17539 5154 17542
rect 5210 17539 5262 17542
rect 5318 17539 5370 17542
rect 5426 17539 5478 17542
rect 5534 17539 5586 17542
rect 5642 17539 5694 17542
rect 5750 17539 5802 17542
rect 5858 17539 5910 17542
rect 5966 17539 6018 17542
rect 6074 17539 6126 17542
rect 6836 17539 6888 17542
rect 6944 17539 6996 17542
rect 7052 17539 7104 17542
rect 7160 17539 7212 17542
rect 7268 17539 7320 17542
rect 7376 17539 7428 17542
rect 7484 17539 7536 17542
rect 7592 17539 7644 17542
rect 7700 17539 7752 17542
rect 7808 17539 7860 17542
rect 7916 17539 7968 17542
rect 8024 17539 8076 17542
rect 8132 17539 8184 17542
rect 8240 17539 8292 17542
rect 8348 17539 8400 17542
rect 8456 17539 8508 17542
rect 8564 17539 8616 17542
rect 8672 17539 8724 17542
rect 8780 17539 8832 17542
rect 9206 17539 9258 17542
rect 9314 17539 9366 17542
rect 9422 17539 9474 17542
rect 9530 17539 9582 17542
rect 9638 17539 9690 17542
rect 9746 17539 9798 17542
rect 9854 17539 9906 17542
rect 9962 17539 10014 17542
rect 10070 17539 10122 17542
rect 10178 17539 10230 17542
rect 10286 17539 10338 17542
rect 10394 17539 10446 17542
rect 10502 17539 10554 17542
rect 10610 17539 10662 17542
rect 10718 17539 10770 17542
rect 10826 17539 10878 17542
rect 10934 17539 10986 17542
rect 11042 17539 11094 17542
rect 11150 17539 11202 17542
rect 1493 17344 1545 17347
rect 1601 17344 1653 17347
rect 3863 17344 3915 17347
rect 3971 17344 4023 17347
rect 6239 17344 6291 17347
rect 6347 17344 6399 17347
rect 6455 17344 6507 17347
rect 6563 17344 6615 17347
rect 6671 17344 6723 17347
rect 8939 17344 8991 17347
rect 9047 17344 9099 17347
rect 11309 17344 11361 17347
rect 11417 17344 11469 17347
rect 1493 17298 1494 17344
rect 1494 17298 1545 17344
rect 1601 17298 1653 17344
rect 3863 17298 3915 17344
rect 3971 17298 4023 17344
rect 6239 17298 6291 17344
rect 6347 17298 6399 17344
rect 6455 17298 6507 17344
rect 6563 17298 6615 17344
rect 6671 17298 6723 17344
rect 8939 17298 8991 17344
rect 9047 17298 9099 17344
rect 11309 17298 11361 17344
rect 11417 17298 11468 17344
rect 11468 17298 11469 17344
rect 1493 17295 1545 17298
rect 1601 17295 1653 17298
rect 3863 17295 3915 17298
rect 3971 17295 4023 17298
rect 6239 17295 6291 17298
rect 6347 17295 6399 17298
rect 6455 17295 6507 17298
rect 6563 17295 6615 17298
rect 6671 17295 6723 17298
rect 8939 17295 8991 17298
rect 9047 17295 9099 17298
rect 11309 17295 11361 17298
rect 11417 17295 11469 17298
rect 1760 17100 1812 17103
rect 1868 17100 1920 17103
rect 1976 17100 2028 17103
rect 2084 17100 2136 17103
rect 2192 17100 2244 17103
rect 2300 17100 2352 17103
rect 2408 17100 2460 17103
rect 2516 17100 2568 17103
rect 2624 17100 2676 17103
rect 2732 17100 2784 17103
rect 2840 17100 2892 17103
rect 2948 17100 3000 17103
rect 3056 17100 3108 17103
rect 3164 17100 3216 17103
rect 3272 17100 3324 17103
rect 3380 17100 3432 17103
rect 3488 17100 3540 17103
rect 3596 17100 3648 17103
rect 3704 17100 3756 17103
rect 4130 17100 4182 17103
rect 4238 17100 4290 17103
rect 4346 17100 4398 17103
rect 4454 17100 4506 17103
rect 4562 17100 4614 17103
rect 4670 17100 4722 17103
rect 4778 17100 4830 17103
rect 4886 17100 4938 17103
rect 4994 17100 5046 17103
rect 5102 17100 5154 17103
rect 5210 17100 5262 17103
rect 5318 17100 5370 17103
rect 5426 17100 5478 17103
rect 5534 17100 5586 17103
rect 5642 17100 5694 17103
rect 5750 17100 5802 17103
rect 5858 17100 5910 17103
rect 5966 17100 6018 17103
rect 6074 17100 6126 17103
rect 6836 17100 6888 17103
rect 6944 17100 6996 17103
rect 7052 17100 7104 17103
rect 7160 17100 7212 17103
rect 7268 17100 7320 17103
rect 7376 17100 7428 17103
rect 7484 17100 7536 17103
rect 7592 17100 7644 17103
rect 7700 17100 7752 17103
rect 7808 17100 7860 17103
rect 7916 17100 7968 17103
rect 8024 17100 8076 17103
rect 8132 17100 8184 17103
rect 8240 17100 8292 17103
rect 8348 17100 8400 17103
rect 8456 17100 8508 17103
rect 8564 17100 8616 17103
rect 8672 17100 8724 17103
rect 8780 17100 8832 17103
rect 9206 17100 9258 17103
rect 9314 17100 9366 17103
rect 9422 17100 9474 17103
rect 9530 17100 9582 17103
rect 9638 17100 9690 17103
rect 9746 17100 9798 17103
rect 9854 17100 9906 17103
rect 9962 17100 10014 17103
rect 10070 17100 10122 17103
rect 10178 17100 10230 17103
rect 10286 17100 10338 17103
rect 10394 17100 10446 17103
rect 10502 17100 10554 17103
rect 10610 17100 10662 17103
rect 10718 17100 10770 17103
rect 10826 17100 10878 17103
rect 10934 17100 10986 17103
rect 11042 17100 11094 17103
rect 11150 17100 11202 17103
rect 1760 17054 1812 17100
rect 1868 17054 1920 17100
rect 1976 17054 2028 17100
rect 2084 17054 2136 17100
rect 2192 17054 2244 17100
rect 2300 17054 2352 17100
rect 2408 17054 2460 17100
rect 2516 17054 2568 17100
rect 2624 17054 2676 17100
rect 2732 17054 2784 17100
rect 2840 17054 2892 17100
rect 2948 17054 3000 17100
rect 3056 17054 3108 17100
rect 3164 17054 3216 17100
rect 3272 17054 3324 17100
rect 3380 17054 3432 17100
rect 3488 17054 3540 17100
rect 3596 17054 3648 17100
rect 3704 17054 3756 17100
rect 4130 17054 4182 17100
rect 4238 17054 4290 17100
rect 4346 17054 4398 17100
rect 4454 17054 4506 17100
rect 4562 17054 4614 17100
rect 4670 17054 4722 17100
rect 4778 17054 4830 17100
rect 4886 17054 4938 17100
rect 4994 17054 5046 17100
rect 5102 17054 5154 17100
rect 5210 17054 5262 17100
rect 5318 17054 5370 17100
rect 5426 17054 5478 17100
rect 5534 17054 5586 17100
rect 5642 17054 5694 17100
rect 5750 17054 5802 17100
rect 5858 17054 5910 17100
rect 5966 17054 6018 17100
rect 6074 17054 6126 17100
rect 6836 17054 6888 17100
rect 6944 17054 6996 17100
rect 7052 17054 7104 17100
rect 7160 17054 7212 17100
rect 7268 17054 7320 17100
rect 7376 17054 7428 17100
rect 7484 17054 7536 17100
rect 7592 17054 7644 17100
rect 7700 17054 7752 17100
rect 7808 17054 7860 17100
rect 7916 17054 7968 17100
rect 8024 17054 8076 17100
rect 8132 17054 8184 17100
rect 8240 17054 8292 17100
rect 8348 17054 8400 17100
rect 8456 17054 8508 17100
rect 8564 17054 8616 17100
rect 8672 17054 8724 17100
rect 8780 17054 8832 17100
rect 9206 17054 9258 17100
rect 9314 17054 9366 17100
rect 9422 17054 9474 17100
rect 9530 17054 9582 17100
rect 9638 17054 9690 17100
rect 9746 17054 9798 17100
rect 9854 17054 9906 17100
rect 9962 17054 10014 17100
rect 10070 17054 10122 17100
rect 10178 17054 10230 17100
rect 10286 17054 10338 17100
rect 10394 17054 10446 17100
rect 10502 17054 10554 17100
rect 10610 17054 10662 17100
rect 10718 17054 10770 17100
rect 10826 17054 10878 17100
rect 10934 17054 10986 17100
rect 11042 17054 11094 17100
rect 11150 17054 11202 17100
rect 1760 17051 1812 17054
rect 1868 17051 1920 17054
rect 1976 17051 2028 17054
rect 2084 17051 2136 17054
rect 2192 17051 2244 17054
rect 2300 17051 2352 17054
rect 2408 17051 2460 17054
rect 2516 17051 2568 17054
rect 2624 17051 2676 17054
rect 2732 17051 2784 17054
rect 2840 17051 2892 17054
rect 2948 17051 3000 17054
rect 3056 17051 3108 17054
rect 3164 17051 3216 17054
rect 3272 17051 3324 17054
rect 3380 17051 3432 17054
rect 3488 17051 3540 17054
rect 3596 17051 3648 17054
rect 3704 17051 3756 17054
rect 4130 17051 4182 17054
rect 4238 17051 4290 17054
rect 4346 17051 4398 17054
rect 4454 17051 4506 17054
rect 4562 17051 4614 17054
rect 4670 17051 4722 17054
rect 4778 17051 4830 17054
rect 4886 17051 4938 17054
rect 4994 17051 5046 17054
rect 5102 17051 5154 17054
rect 5210 17051 5262 17054
rect 5318 17051 5370 17054
rect 5426 17051 5478 17054
rect 5534 17051 5586 17054
rect 5642 17051 5694 17054
rect 5750 17051 5802 17054
rect 5858 17051 5910 17054
rect 5966 17051 6018 17054
rect 6074 17051 6126 17054
rect 6836 17051 6888 17054
rect 6944 17051 6996 17054
rect 7052 17051 7104 17054
rect 7160 17051 7212 17054
rect 7268 17051 7320 17054
rect 7376 17051 7428 17054
rect 7484 17051 7536 17054
rect 7592 17051 7644 17054
rect 7700 17051 7752 17054
rect 7808 17051 7860 17054
rect 7916 17051 7968 17054
rect 8024 17051 8076 17054
rect 8132 17051 8184 17054
rect 8240 17051 8292 17054
rect 8348 17051 8400 17054
rect 8456 17051 8508 17054
rect 8564 17051 8616 17054
rect 8672 17051 8724 17054
rect 8780 17051 8832 17054
rect 9206 17051 9258 17054
rect 9314 17051 9366 17054
rect 9422 17051 9474 17054
rect 9530 17051 9582 17054
rect 9638 17051 9690 17054
rect 9746 17051 9798 17054
rect 9854 17051 9906 17054
rect 9962 17051 10014 17054
rect 10070 17051 10122 17054
rect 10178 17051 10230 17054
rect 10286 17051 10338 17054
rect 10394 17051 10446 17054
rect 10502 17051 10554 17054
rect 10610 17051 10662 17054
rect 10718 17051 10770 17054
rect 10826 17051 10878 17054
rect 10934 17051 10986 17054
rect 11042 17051 11094 17054
rect 11150 17051 11202 17054
rect 1493 16856 1545 16859
rect 1601 16856 1653 16859
rect 3863 16856 3915 16859
rect 3971 16856 4023 16859
rect 6239 16856 6291 16859
rect 6347 16856 6399 16859
rect 6455 16856 6507 16859
rect 6563 16856 6615 16859
rect 6671 16856 6723 16859
rect 8939 16856 8991 16859
rect 9047 16856 9099 16859
rect 11309 16856 11361 16859
rect 11417 16856 11469 16859
rect 1493 16810 1494 16856
rect 1494 16810 1545 16856
rect 1601 16810 1653 16856
rect 3863 16810 3915 16856
rect 3971 16810 4023 16856
rect 6239 16810 6291 16856
rect 6347 16810 6399 16856
rect 6455 16810 6507 16856
rect 6563 16810 6615 16856
rect 6671 16810 6723 16856
rect 8939 16810 8991 16856
rect 9047 16810 9099 16856
rect 11309 16810 11361 16856
rect 11417 16810 11468 16856
rect 11468 16810 11469 16856
rect 1493 16807 1545 16810
rect 1601 16807 1653 16810
rect 3863 16807 3915 16810
rect 3971 16807 4023 16810
rect 6239 16807 6291 16810
rect 6347 16807 6399 16810
rect 6455 16807 6507 16810
rect 6563 16807 6615 16810
rect 6671 16807 6723 16810
rect 8939 16807 8991 16810
rect 9047 16807 9099 16810
rect 11309 16807 11361 16810
rect 11417 16807 11469 16810
rect 1760 16612 1812 16615
rect 1868 16612 1920 16615
rect 1976 16612 2028 16615
rect 2084 16612 2136 16615
rect 2192 16612 2244 16615
rect 2300 16612 2352 16615
rect 2408 16612 2460 16615
rect 2516 16612 2568 16615
rect 2624 16612 2676 16615
rect 2732 16612 2784 16615
rect 2840 16612 2892 16615
rect 2948 16612 3000 16615
rect 3056 16612 3108 16615
rect 3164 16612 3216 16615
rect 3272 16612 3324 16615
rect 3380 16612 3432 16615
rect 3488 16612 3540 16615
rect 3596 16612 3648 16615
rect 3704 16612 3756 16615
rect 4130 16612 4182 16615
rect 4238 16612 4290 16615
rect 4346 16612 4398 16615
rect 4454 16612 4506 16615
rect 4562 16612 4614 16615
rect 4670 16612 4722 16615
rect 4778 16612 4830 16615
rect 4886 16612 4938 16615
rect 4994 16612 5046 16615
rect 5102 16612 5154 16615
rect 5210 16612 5262 16615
rect 5318 16612 5370 16615
rect 5426 16612 5478 16615
rect 5534 16612 5586 16615
rect 5642 16612 5694 16615
rect 5750 16612 5802 16615
rect 5858 16612 5910 16615
rect 5966 16612 6018 16615
rect 6074 16612 6126 16615
rect 6836 16612 6888 16615
rect 6944 16612 6996 16615
rect 7052 16612 7104 16615
rect 7160 16612 7212 16615
rect 7268 16612 7320 16615
rect 7376 16612 7428 16615
rect 7484 16612 7536 16615
rect 7592 16612 7644 16615
rect 7700 16612 7752 16615
rect 7808 16612 7860 16615
rect 7916 16612 7968 16615
rect 8024 16612 8076 16615
rect 8132 16612 8184 16615
rect 8240 16612 8292 16615
rect 8348 16612 8400 16615
rect 8456 16612 8508 16615
rect 8564 16612 8616 16615
rect 8672 16612 8724 16615
rect 8780 16612 8832 16615
rect 9206 16612 9258 16615
rect 9314 16612 9366 16615
rect 9422 16612 9474 16615
rect 9530 16612 9582 16615
rect 9638 16612 9690 16615
rect 9746 16612 9798 16615
rect 9854 16612 9906 16615
rect 9962 16612 10014 16615
rect 10070 16612 10122 16615
rect 10178 16612 10230 16615
rect 10286 16612 10338 16615
rect 10394 16612 10446 16615
rect 10502 16612 10554 16615
rect 10610 16612 10662 16615
rect 10718 16612 10770 16615
rect 10826 16612 10878 16615
rect 10934 16612 10986 16615
rect 11042 16612 11094 16615
rect 11150 16612 11202 16615
rect 1760 16566 1812 16612
rect 1868 16566 1920 16612
rect 1976 16566 2028 16612
rect 2084 16566 2136 16612
rect 2192 16566 2244 16612
rect 2300 16566 2352 16612
rect 2408 16566 2460 16612
rect 2516 16566 2568 16612
rect 2624 16566 2676 16612
rect 2732 16566 2784 16612
rect 2840 16566 2892 16612
rect 2948 16566 3000 16612
rect 3056 16566 3108 16612
rect 3164 16566 3216 16612
rect 3272 16566 3324 16612
rect 3380 16566 3432 16612
rect 3488 16566 3540 16612
rect 3596 16566 3648 16612
rect 3704 16566 3756 16612
rect 4130 16566 4182 16612
rect 4238 16566 4290 16612
rect 4346 16566 4398 16612
rect 4454 16566 4506 16612
rect 4562 16566 4614 16612
rect 4670 16566 4722 16612
rect 4778 16566 4830 16612
rect 4886 16566 4938 16612
rect 4994 16566 5046 16612
rect 5102 16566 5154 16612
rect 5210 16566 5262 16612
rect 5318 16566 5370 16612
rect 5426 16566 5478 16612
rect 5534 16566 5586 16612
rect 5642 16566 5694 16612
rect 5750 16566 5802 16612
rect 5858 16566 5910 16612
rect 5966 16566 6018 16612
rect 6074 16566 6126 16612
rect 6836 16566 6888 16612
rect 6944 16566 6996 16612
rect 7052 16566 7104 16612
rect 7160 16566 7212 16612
rect 7268 16566 7320 16612
rect 7376 16566 7428 16612
rect 7484 16566 7536 16612
rect 7592 16566 7644 16612
rect 7700 16566 7752 16612
rect 7808 16566 7860 16612
rect 7916 16566 7968 16612
rect 8024 16566 8076 16612
rect 8132 16566 8184 16612
rect 8240 16566 8292 16612
rect 8348 16566 8400 16612
rect 8456 16566 8508 16612
rect 8564 16566 8616 16612
rect 8672 16566 8724 16612
rect 8780 16566 8832 16612
rect 9206 16566 9258 16612
rect 9314 16566 9366 16612
rect 9422 16566 9474 16612
rect 9530 16566 9582 16612
rect 9638 16566 9690 16612
rect 9746 16566 9798 16612
rect 9854 16566 9906 16612
rect 9962 16566 10014 16612
rect 10070 16566 10122 16612
rect 10178 16566 10230 16612
rect 10286 16566 10338 16612
rect 10394 16566 10446 16612
rect 10502 16566 10554 16612
rect 10610 16566 10662 16612
rect 10718 16566 10770 16612
rect 10826 16566 10878 16612
rect 10934 16566 10986 16612
rect 11042 16566 11094 16612
rect 11150 16566 11202 16612
rect 1760 16563 1812 16566
rect 1868 16563 1920 16566
rect 1976 16563 2028 16566
rect 2084 16563 2136 16566
rect 2192 16563 2244 16566
rect 2300 16563 2352 16566
rect 2408 16563 2460 16566
rect 2516 16563 2568 16566
rect 2624 16563 2676 16566
rect 2732 16563 2784 16566
rect 2840 16563 2892 16566
rect 2948 16563 3000 16566
rect 3056 16563 3108 16566
rect 3164 16563 3216 16566
rect 3272 16563 3324 16566
rect 3380 16563 3432 16566
rect 3488 16563 3540 16566
rect 3596 16563 3648 16566
rect 3704 16563 3756 16566
rect 4130 16563 4182 16566
rect 4238 16563 4290 16566
rect 4346 16563 4398 16566
rect 4454 16563 4506 16566
rect 4562 16563 4614 16566
rect 4670 16563 4722 16566
rect 4778 16563 4830 16566
rect 4886 16563 4938 16566
rect 4994 16563 5046 16566
rect 5102 16563 5154 16566
rect 5210 16563 5262 16566
rect 5318 16563 5370 16566
rect 5426 16563 5478 16566
rect 5534 16563 5586 16566
rect 5642 16563 5694 16566
rect 5750 16563 5802 16566
rect 5858 16563 5910 16566
rect 5966 16563 6018 16566
rect 6074 16563 6126 16566
rect 6836 16563 6888 16566
rect 6944 16563 6996 16566
rect 7052 16563 7104 16566
rect 7160 16563 7212 16566
rect 7268 16563 7320 16566
rect 7376 16563 7428 16566
rect 7484 16563 7536 16566
rect 7592 16563 7644 16566
rect 7700 16563 7752 16566
rect 7808 16563 7860 16566
rect 7916 16563 7968 16566
rect 8024 16563 8076 16566
rect 8132 16563 8184 16566
rect 8240 16563 8292 16566
rect 8348 16563 8400 16566
rect 8456 16563 8508 16566
rect 8564 16563 8616 16566
rect 8672 16563 8724 16566
rect 8780 16563 8832 16566
rect 9206 16563 9258 16566
rect 9314 16563 9366 16566
rect 9422 16563 9474 16566
rect 9530 16563 9582 16566
rect 9638 16563 9690 16566
rect 9746 16563 9798 16566
rect 9854 16563 9906 16566
rect 9962 16563 10014 16566
rect 10070 16563 10122 16566
rect 10178 16563 10230 16566
rect 10286 16563 10338 16566
rect 10394 16563 10446 16566
rect 10502 16563 10554 16566
rect 10610 16563 10662 16566
rect 10718 16563 10770 16566
rect 10826 16563 10878 16566
rect 10934 16563 10986 16566
rect 11042 16563 11094 16566
rect 11150 16563 11202 16566
rect 1493 16368 1545 16371
rect 1601 16368 1653 16371
rect 3863 16368 3915 16371
rect 3971 16368 4023 16371
rect 6239 16368 6291 16371
rect 6347 16368 6399 16371
rect 6455 16368 6507 16371
rect 6563 16368 6615 16371
rect 6671 16368 6723 16371
rect 8939 16368 8991 16371
rect 9047 16368 9099 16371
rect 11309 16368 11361 16371
rect 11417 16368 11469 16371
rect 1493 16322 1494 16368
rect 1494 16322 1545 16368
rect 1601 16322 1653 16368
rect 3863 16322 3915 16368
rect 3971 16322 4023 16368
rect 6239 16322 6291 16368
rect 6347 16322 6399 16368
rect 6455 16322 6507 16368
rect 6563 16322 6615 16368
rect 6671 16322 6723 16368
rect 8939 16322 8991 16368
rect 9047 16322 9099 16368
rect 11309 16322 11361 16368
rect 11417 16322 11468 16368
rect 11468 16322 11469 16368
rect 1493 16319 1545 16322
rect 1601 16319 1653 16322
rect 3863 16319 3915 16322
rect 3971 16319 4023 16322
rect 6239 16319 6291 16322
rect 6347 16319 6399 16322
rect 6455 16319 6507 16322
rect 6563 16319 6615 16322
rect 6671 16319 6723 16322
rect 8939 16319 8991 16322
rect 9047 16319 9099 16322
rect 11309 16319 11361 16322
rect 11417 16319 11469 16322
rect 1760 16124 1812 16127
rect 1868 16124 1920 16127
rect 1976 16124 2028 16127
rect 2084 16124 2136 16127
rect 2192 16124 2244 16127
rect 2300 16124 2352 16127
rect 2408 16124 2460 16127
rect 2516 16124 2568 16127
rect 2624 16124 2676 16127
rect 2732 16124 2784 16127
rect 2840 16124 2892 16127
rect 2948 16124 3000 16127
rect 3056 16124 3108 16127
rect 3164 16124 3216 16127
rect 3272 16124 3324 16127
rect 3380 16124 3432 16127
rect 3488 16124 3540 16127
rect 3596 16124 3648 16127
rect 3704 16124 3756 16127
rect 4130 16124 4182 16127
rect 4238 16124 4290 16127
rect 4346 16124 4398 16127
rect 4454 16124 4506 16127
rect 4562 16124 4614 16127
rect 4670 16124 4722 16127
rect 4778 16124 4830 16127
rect 4886 16124 4938 16127
rect 4994 16124 5046 16127
rect 5102 16124 5154 16127
rect 5210 16124 5262 16127
rect 5318 16124 5370 16127
rect 5426 16124 5478 16127
rect 5534 16124 5586 16127
rect 5642 16124 5694 16127
rect 5750 16124 5802 16127
rect 5858 16124 5910 16127
rect 5966 16124 6018 16127
rect 6074 16124 6126 16127
rect 6836 16124 6888 16127
rect 6944 16124 6996 16127
rect 7052 16124 7104 16127
rect 7160 16124 7212 16127
rect 7268 16124 7320 16127
rect 7376 16124 7428 16127
rect 7484 16124 7536 16127
rect 7592 16124 7644 16127
rect 7700 16124 7752 16127
rect 7808 16124 7860 16127
rect 7916 16124 7968 16127
rect 8024 16124 8076 16127
rect 8132 16124 8184 16127
rect 8240 16124 8292 16127
rect 8348 16124 8400 16127
rect 8456 16124 8508 16127
rect 8564 16124 8616 16127
rect 8672 16124 8724 16127
rect 8780 16124 8832 16127
rect 9206 16124 9258 16127
rect 9314 16124 9366 16127
rect 9422 16124 9474 16127
rect 9530 16124 9582 16127
rect 9638 16124 9690 16127
rect 9746 16124 9798 16127
rect 9854 16124 9906 16127
rect 9962 16124 10014 16127
rect 10070 16124 10122 16127
rect 10178 16124 10230 16127
rect 10286 16124 10338 16127
rect 10394 16124 10446 16127
rect 10502 16124 10554 16127
rect 10610 16124 10662 16127
rect 10718 16124 10770 16127
rect 10826 16124 10878 16127
rect 10934 16124 10986 16127
rect 11042 16124 11094 16127
rect 11150 16124 11202 16127
rect 1760 16078 1812 16124
rect 1868 16078 1920 16124
rect 1976 16078 2028 16124
rect 2084 16078 2136 16124
rect 2192 16078 2244 16124
rect 2300 16078 2352 16124
rect 2408 16078 2460 16124
rect 2516 16078 2568 16124
rect 2624 16078 2676 16124
rect 2732 16078 2784 16124
rect 2840 16078 2892 16124
rect 2948 16078 3000 16124
rect 3056 16078 3108 16124
rect 3164 16078 3216 16124
rect 3272 16078 3324 16124
rect 3380 16078 3432 16124
rect 3488 16078 3540 16124
rect 3596 16078 3648 16124
rect 3704 16078 3756 16124
rect 4130 16078 4182 16124
rect 4238 16078 4290 16124
rect 4346 16078 4398 16124
rect 4454 16078 4506 16124
rect 4562 16078 4614 16124
rect 4670 16078 4722 16124
rect 4778 16078 4830 16124
rect 4886 16078 4938 16124
rect 4994 16078 5046 16124
rect 5102 16078 5154 16124
rect 5210 16078 5262 16124
rect 5318 16078 5370 16124
rect 5426 16078 5478 16124
rect 5534 16078 5586 16124
rect 5642 16078 5694 16124
rect 5750 16078 5802 16124
rect 5858 16078 5910 16124
rect 5966 16078 6018 16124
rect 6074 16078 6126 16124
rect 6836 16078 6888 16124
rect 6944 16078 6996 16124
rect 7052 16078 7104 16124
rect 7160 16078 7212 16124
rect 7268 16078 7320 16124
rect 7376 16078 7428 16124
rect 7484 16078 7536 16124
rect 7592 16078 7644 16124
rect 7700 16078 7752 16124
rect 7808 16078 7860 16124
rect 7916 16078 7968 16124
rect 8024 16078 8076 16124
rect 8132 16078 8184 16124
rect 8240 16078 8292 16124
rect 8348 16078 8400 16124
rect 8456 16078 8508 16124
rect 8564 16078 8616 16124
rect 8672 16078 8724 16124
rect 8780 16078 8832 16124
rect 9206 16078 9258 16124
rect 9314 16078 9366 16124
rect 9422 16078 9474 16124
rect 9530 16078 9582 16124
rect 9638 16078 9690 16124
rect 9746 16078 9798 16124
rect 9854 16078 9906 16124
rect 9962 16078 10014 16124
rect 10070 16078 10122 16124
rect 10178 16078 10230 16124
rect 10286 16078 10338 16124
rect 10394 16078 10446 16124
rect 10502 16078 10554 16124
rect 10610 16078 10662 16124
rect 10718 16078 10770 16124
rect 10826 16078 10878 16124
rect 10934 16078 10986 16124
rect 11042 16078 11094 16124
rect 11150 16078 11202 16124
rect 1760 16075 1812 16078
rect 1868 16075 1920 16078
rect 1976 16075 2028 16078
rect 2084 16075 2136 16078
rect 2192 16075 2244 16078
rect 2300 16075 2352 16078
rect 2408 16075 2460 16078
rect 2516 16075 2568 16078
rect 2624 16075 2676 16078
rect 2732 16075 2784 16078
rect 2840 16075 2892 16078
rect 2948 16075 3000 16078
rect 3056 16075 3108 16078
rect 3164 16075 3216 16078
rect 3272 16075 3324 16078
rect 3380 16075 3432 16078
rect 3488 16075 3540 16078
rect 3596 16075 3648 16078
rect 3704 16075 3756 16078
rect 4130 16075 4182 16078
rect 4238 16075 4290 16078
rect 4346 16075 4398 16078
rect 4454 16075 4506 16078
rect 4562 16075 4614 16078
rect 4670 16075 4722 16078
rect 4778 16075 4830 16078
rect 4886 16075 4938 16078
rect 4994 16075 5046 16078
rect 5102 16075 5154 16078
rect 5210 16075 5262 16078
rect 5318 16075 5370 16078
rect 5426 16075 5478 16078
rect 5534 16075 5586 16078
rect 5642 16075 5694 16078
rect 5750 16075 5802 16078
rect 5858 16075 5910 16078
rect 5966 16075 6018 16078
rect 6074 16075 6126 16078
rect 6836 16075 6888 16078
rect 6944 16075 6996 16078
rect 7052 16075 7104 16078
rect 7160 16075 7212 16078
rect 7268 16075 7320 16078
rect 7376 16075 7428 16078
rect 7484 16075 7536 16078
rect 7592 16075 7644 16078
rect 7700 16075 7752 16078
rect 7808 16075 7860 16078
rect 7916 16075 7968 16078
rect 8024 16075 8076 16078
rect 8132 16075 8184 16078
rect 8240 16075 8292 16078
rect 8348 16075 8400 16078
rect 8456 16075 8508 16078
rect 8564 16075 8616 16078
rect 8672 16075 8724 16078
rect 8780 16075 8832 16078
rect 9206 16075 9258 16078
rect 9314 16075 9366 16078
rect 9422 16075 9474 16078
rect 9530 16075 9582 16078
rect 9638 16075 9690 16078
rect 9746 16075 9798 16078
rect 9854 16075 9906 16078
rect 9962 16075 10014 16078
rect 10070 16075 10122 16078
rect 10178 16075 10230 16078
rect 10286 16075 10338 16078
rect 10394 16075 10446 16078
rect 10502 16075 10554 16078
rect 10610 16075 10662 16078
rect 10718 16075 10770 16078
rect 10826 16075 10878 16078
rect 10934 16075 10986 16078
rect 11042 16075 11094 16078
rect 11150 16075 11202 16078
rect 1493 15880 1545 15883
rect 1601 15880 1653 15883
rect 3863 15880 3915 15883
rect 3971 15880 4023 15883
rect 6239 15880 6291 15883
rect 6347 15880 6399 15883
rect 6455 15880 6507 15883
rect 6563 15880 6615 15883
rect 6671 15880 6723 15883
rect 8939 15880 8991 15883
rect 9047 15880 9099 15883
rect 11309 15880 11361 15883
rect 11417 15880 11469 15883
rect 1493 15834 1494 15880
rect 1494 15834 1545 15880
rect 1601 15834 1653 15880
rect 3863 15834 3915 15880
rect 3971 15834 4023 15880
rect 6239 15834 6291 15880
rect 6347 15834 6399 15880
rect 6455 15834 6507 15880
rect 6563 15834 6615 15880
rect 6671 15834 6723 15880
rect 8939 15834 8991 15880
rect 9047 15834 9099 15880
rect 11309 15834 11361 15880
rect 11417 15834 11468 15880
rect 11468 15834 11469 15880
rect 1493 15831 1545 15834
rect 1601 15831 1653 15834
rect 3863 15831 3915 15834
rect 3971 15831 4023 15834
rect 6239 15831 6291 15834
rect 6347 15831 6399 15834
rect 6455 15831 6507 15834
rect 6563 15831 6615 15834
rect 6671 15831 6723 15834
rect 8939 15831 8991 15834
rect 9047 15831 9099 15834
rect 11309 15831 11361 15834
rect 11417 15831 11469 15834
rect 1760 15636 1812 15639
rect 1868 15636 1920 15639
rect 1976 15636 2028 15639
rect 2084 15636 2136 15639
rect 2192 15636 2244 15639
rect 2300 15636 2352 15639
rect 2408 15636 2460 15639
rect 2516 15636 2568 15639
rect 2624 15636 2676 15639
rect 2732 15636 2784 15639
rect 2840 15636 2892 15639
rect 2948 15636 3000 15639
rect 3056 15636 3108 15639
rect 3164 15636 3216 15639
rect 3272 15636 3324 15639
rect 3380 15636 3432 15639
rect 3488 15636 3540 15639
rect 3596 15636 3648 15639
rect 3704 15636 3756 15639
rect 4130 15636 4182 15639
rect 4238 15636 4290 15639
rect 4346 15636 4398 15639
rect 4454 15636 4506 15639
rect 4562 15636 4614 15639
rect 4670 15636 4722 15639
rect 4778 15636 4830 15639
rect 4886 15636 4938 15639
rect 4994 15636 5046 15639
rect 5102 15636 5154 15639
rect 5210 15636 5262 15639
rect 5318 15636 5370 15639
rect 5426 15636 5478 15639
rect 5534 15636 5586 15639
rect 5642 15636 5694 15639
rect 5750 15636 5802 15639
rect 5858 15636 5910 15639
rect 5966 15636 6018 15639
rect 6074 15636 6126 15639
rect 6836 15636 6888 15639
rect 6944 15636 6996 15639
rect 7052 15636 7104 15639
rect 7160 15636 7212 15639
rect 7268 15636 7320 15639
rect 7376 15636 7428 15639
rect 7484 15636 7536 15639
rect 7592 15636 7644 15639
rect 7700 15636 7752 15639
rect 7808 15636 7860 15639
rect 7916 15636 7968 15639
rect 8024 15636 8076 15639
rect 8132 15636 8184 15639
rect 8240 15636 8292 15639
rect 8348 15636 8400 15639
rect 8456 15636 8508 15639
rect 8564 15636 8616 15639
rect 8672 15636 8724 15639
rect 8780 15636 8832 15639
rect 9206 15636 9258 15639
rect 9314 15636 9366 15639
rect 9422 15636 9474 15639
rect 9530 15636 9582 15639
rect 9638 15636 9690 15639
rect 9746 15636 9798 15639
rect 9854 15636 9906 15639
rect 9962 15636 10014 15639
rect 10070 15636 10122 15639
rect 10178 15636 10230 15639
rect 10286 15636 10338 15639
rect 10394 15636 10446 15639
rect 10502 15636 10554 15639
rect 10610 15636 10662 15639
rect 10718 15636 10770 15639
rect 10826 15636 10878 15639
rect 10934 15636 10986 15639
rect 11042 15636 11094 15639
rect 11150 15636 11202 15639
rect 1760 15590 1812 15636
rect 1868 15590 1920 15636
rect 1976 15590 2028 15636
rect 2084 15590 2136 15636
rect 2192 15590 2244 15636
rect 2300 15590 2352 15636
rect 2408 15590 2460 15636
rect 2516 15590 2568 15636
rect 2624 15590 2676 15636
rect 2732 15590 2784 15636
rect 2840 15590 2892 15636
rect 2948 15590 3000 15636
rect 3056 15590 3108 15636
rect 3164 15590 3216 15636
rect 3272 15590 3324 15636
rect 3380 15590 3432 15636
rect 3488 15590 3540 15636
rect 3596 15590 3648 15636
rect 3704 15590 3756 15636
rect 4130 15590 4182 15636
rect 4238 15590 4290 15636
rect 4346 15590 4398 15636
rect 4454 15590 4506 15636
rect 4562 15590 4614 15636
rect 4670 15590 4722 15636
rect 4778 15590 4830 15636
rect 4886 15590 4938 15636
rect 4994 15590 5046 15636
rect 5102 15590 5154 15636
rect 5210 15590 5262 15636
rect 5318 15590 5370 15636
rect 5426 15590 5478 15636
rect 5534 15590 5586 15636
rect 5642 15590 5694 15636
rect 5750 15590 5802 15636
rect 5858 15590 5910 15636
rect 5966 15590 6018 15636
rect 6074 15590 6126 15636
rect 6836 15590 6888 15636
rect 6944 15590 6996 15636
rect 7052 15590 7104 15636
rect 7160 15590 7212 15636
rect 7268 15590 7320 15636
rect 7376 15590 7428 15636
rect 7484 15590 7536 15636
rect 7592 15590 7644 15636
rect 7700 15590 7752 15636
rect 7808 15590 7860 15636
rect 7916 15590 7968 15636
rect 8024 15590 8076 15636
rect 8132 15590 8184 15636
rect 8240 15590 8292 15636
rect 8348 15590 8400 15636
rect 8456 15590 8508 15636
rect 8564 15590 8616 15636
rect 8672 15590 8724 15636
rect 8780 15590 8832 15636
rect 9206 15590 9258 15636
rect 9314 15590 9366 15636
rect 9422 15590 9474 15636
rect 9530 15590 9582 15636
rect 9638 15590 9690 15636
rect 9746 15590 9798 15636
rect 9854 15590 9906 15636
rect 9962 15590 10014 15636
rect 10070 15590 10122 15636
rect 10178 15590 10230 15636
rect 10286 15590 10338 15636
rect 10394 15590 10446 15636
rect 10502 15590 10554 15636
rect 10610 15590 10662 15636
rect 10718 15590 10770 15636
rect 10826 15590 10878 15636
rect 10934 15590 10986 15636
rect 11042 15590 11094 15636
rect 11150 15590 11202 15636
rect 1760 15587 1812 15590
rect 1868 15587 1920 15590
rect 1976 15587 2028 15590
rect 2084 15587 2136 15590
rect 2192 15587 2244 15590
rect 2300 15587 2352 15590
rect 2408 15587 2460 15590
rect 2516 15587 2568 15590
rect 2624 15587 2676 15590
rect 2732 15587 2784 15590
rect 2840 15587 2892 15590
rect 2948 15587 3000 15590
rect 3056 15587 3108 15590
rect 3164 15587 3216 15590
rect 3272 15587 3324 15590
rect 3380 15587 3432 15590
rect 3488 15587 3540 15590
rect 3596 15587 3648 15590
rect 3704 15587 3756 15590
rect 4130 15587 4182 15590
rect 4238 15587 4290 15590
rect 4346 15587 4398 15590
rect 4454 15587 4506 15590
rect 4562 15587 4614 15590
rect 4670 15587 4722 15590
rect 4778 15587 4830 15590
rect 4886 15587 4938 15590
rect 4994 15587 5046 15590
rect 5102 15587 5154 15590
rect 5210 15587 5262 15590
rect 5318 15587 5370 15590
rect 5426 15587 5478 15590
rect 5534 15587 5586 15590
rect 5642 15587 5694 15590
rect 5750 15587 5802 15590
rect 5858 15587 5910 15590
rect 5966 15587 6018 15590
rect 6074 15587 6126 15590
rect 6836 15587 6888 15590
rect 6944 15587 6996 15590
rect 7052 15587 7104 15590
rect 7160 15587 7212 15590
rect 7268 15587 7320 15590
rect 7376 15587 7428 15590
rect 7484 15587 7536 15590
rect 7592 15587 7644 15590
rect 7700 15587 7752 15590
rect 7808 15587 7860 15590
rect 7916 15587 7968 15590
rect 8024 15587 8076 15590
rect 8132 15587 8184 15590
rect 8240 15587 8292 15590
rect 8348 15587 8400 15590
rect 8456 15587 8508 15590
rect 8564 15587 8616 15590
rect 8672 15587 8724 15590
rect 8780 15587 8832 15590
rect 9206 15587 9258 15590
rect 9314 15587 9366 15590
rect 9422 15587 9474 15590
rect 9530 15587 9582 15590
rect 9638 15587 9690 15590
rect 9746 15587 9798 15590
rect 9854 15587 9906 15590
rect 9962 15587 10014 15590
rect 10070 15587 10122 15590
rect 10178 15587 10230 15590
rect 10286 15587 10338 15590
rect 10394 15587 10446 15590
rect 10502 15587 10554 15590
rect 10610 15587 10662 15590
rect 10718 15587 10770 15590
rect 10826 15587 10878 15590
rect 10934 15587 10986 15590
rect 11042 15587 11094 15590
rect 11150 15587 11202 15590
rect 1493 15392 1545 15395
rect 1601 15392 1653 15395
rect 3863 15392 3915 15395
rect 3971 15392 4023 15395
rect 6239 15392 6291 15395
rect 6347 15392 6399 15395
rect 6455 15392 6507 15395
rect 6563 15392 6615 15395
rect 6671 15392 6723 15395
rect 8939 15392 8991 15395
rect 9047 15392 9099 15395
rect 11309 15392 11361 15395
rect 11417 15392 11469 15395
rect 1493 15346 1494 15392
rect 1494 15346 1545 15392
rect 1601 15346 1653 15392
rect 3863 15346 3915 15392
rect 3971 15346 4023 15392
rect 6239 15346 6291 15392
rect 6347 15346 6399 15392
rect 6455 15346 6507 15392
rect 6563 15346 6615 15392
rect 6671 15346 6723 15392
rect 8939 15346 8991 15392
rect 9047 15346 9099 15392
rect 11309 15346 11361 15392
rect 11417 15346 11468 15392
rect 11468 15346 11469 15392
rect 1493 15343 1545 15346
rect 1601 15343 1653 15346
rect 3863 15343 3915 15346
rect 3971 15343 4023 15346
rect 6239 15343 6291 15346
rect 6347 15343 6399 15346
rect 6455 15343 6507 15346
rect 6563 15343 6615 15346
rect 6671 15343 6723 15346
rect 8939 15343 8991 15346
rect 9047 15343 9099 15346
rect 11309 15343 11361 15346
rect 11417 15343 11469 15346
rect 1760 15148 1812 15151
rect 1868 15148 1920 15151
rect 1976 15148 2028 15151
rect 2084 15148 2136 15151
rect 2192 15148 2244 15151
rect 2300 15148 2352 15151
rect 2408 15148 2460 15151
rect 2516 15148 2568 15151
rect 2624 15148 2676 15151
rect 2732 15148 2784 15151
rect 2840 15148 2892 15151
rect 2948 15148 3000 15151
rect 3056 15148 3108 15151
rect 3164 15148 3216 15151
rect 3272 15148 3324 15151
rect 3380 15148 3432 15151
rect 3488 15148 3540 15151
rect 3596 15148 3648 15151
rect 3704 15148 3756 15151
rect 4130 15148 4182 15151
rect 4238 15148 4290 15151
rect 4346 15148 4398 15151
rect 4454 15148 4506 15151
rect 4562 15148 4614 15151
rect 4670 15148 4722 15151
rect 4778 15148 4830 15151
rect 4886 15148 4938 15151
rect 4994 15148 5046 15151
rect 5102 15148 5154 15151
rect 5210 15148 5262 15151
rect 5318 15148 5370 15151
rect 5426 15148 5478 15151
rect 5534 15148 5586 15151
rect 5642 15148 5694 15151
rect 5750 15148 5802 15151
rect 5858 15148 5910 15151
rect 5966 15148 6018 15151
rect 6074 15148 6126 15151
rect 6836 15148 6888 15151
rect 6944 15148 6996 15151
rect 7052 15148 7104 15151
rect 7160 15148 7212 15151
rect 7268 15148 7320 15151
rect 7376 15148 7428 15151
rect 7484 15148 7536 15151
rect 7592 15148 7644 15151
rect 7700 15148 7752 15151
rect 7808 15148 7860 15151
rect 7916 15148 7968 15151
rect 8024 15148 8076 15151
rect 8132 15148 8184 15151
rect 8240 15148 8292 15151
rect 8348 15148 8400 15151
rect 8456 15148 8508 15151
rect 8564 15148 8616 15151
rect 8672 15148 8724 15151
rect 8780 15148 8832 15151
rect 9206 15148 9258 15151
rect 9314 15148 9366 15151
rect 9422 15148 9474 15151
rect 9530 15148 9582 15151
rect 9638 15148 9690 15151
rect 9746 15148 9798 15151
rect 9854 15148 9906 15151
rect 9962 15148 10014 15151
rect 10070 15148 10122 15151
rect 10178 15148 10230 15151
rect 10286 15148 10338 15151
rect 10394 15148 10446 15151
rect 10502 15148 10554 15151
rect 10610 15148 10662 15151
rect 10718 15148 10770 15151
rect 10826 15148 10878 15151
rect 10934 15148 10986 15151
rect 11042 15148 11094 15151
rect 11150 15148 11202 15151
rect 1760 15102 1812 15148
rect 1868 15102 1920 15148
rect 1976 15102 2028 15148
rect 2084 15102 2136 15148
rect 2192 15102 2244 15148
rect 2300 15102 2352 15148
rect 2408 15102 2460 15148
rect 2516 15102 2568 15148
rect 2624 15102 2676 15148
rect 2732 15102 2784 15148
rect 2840 15102 2892 15148
rect 2948 15102 3000 15148
rect 3056 15102 3108 15148
rect 3164 15102 3216 15148
rect 3272 15102 3324 15148
rect 3380 15102 3432 15148
rect 3488 15102 3540 15148
rect 3596 15102 3648 15148
rect 3704 15102 3756 15148
rect 4130 15102 4182 15148
rect 4238 15102 4290 15148
rect 4346 15102 4398 15148
rect 4454 15102 4506 15148
rect 4562 15102 4614 15148
rect 4670 15102 4722 15148
rect 4778 15102 4830 15148
rect 4886 15102 4938 15148
rect 4994 15102 5046 15148
rect 5102 15102 5154 15148
rect 5210 15102 5262 15148
rect 5318 15102 5370 15148
rect 5426 15102 5478 15148
rect 5534 15102 5586 15148
rect 5642 15102 5694 15148
rect 5750 15102 5802 15148
rect 5858 15102 5910 15148
rect 5966 15102 6018 15148
rect 6074 15102 6126 15148
rect 6836 15102 6888 15148
rect 6944 15102 6996 15148
rect 7052 15102 7104 15148
rect 7160 15102 7212 15148
rect 7268 15102 7320 15148
rect 7376 15102 7428 15148
rect 7484 15102 7536 15148
rect 7592 15102 7644 15148
rect 7700 15102 7752 15148
rect 7808 15102 7860 15148
rect 7916 15102 7968 15148
rect 8024 15102 8076 15148
rect 8132 15102 8184 15148
rect 8240 15102 8292 15148
rect 8348 15102 8400 15148
rect 8456 15102 8508 15148
rect 8564 15102 8616 15148
rect 8672 15102 8724 15148
rect 8780 15102 8832 15148
rect 9206 15102 9258 15148
rect 9314 15102 9366 15148
rect 9422 15102 9474 15148
rect 9530 15102 9582 15148
rect 9638 15102 9690 15148
rect 9746 15102 9798 15148
rect 9854 15102 9906 15148
rect 9962 15102 10014 15148
rect 10070 15102 10122 15148
rect 10178 15102 10230 15148
rect 10286 15102 10338 15148
rect 10394 15102 10446 15148
rect 10502 15102 10554 15148
rect 10610 15102 10662 15148
rect 10718 15102 10770 15148
rect 10826 15102 10878 15148
rect 10934 15102 10986 15148
rect 11042 15102 11094 15148
rect 11150 15102 11202 15148
rect 1760 15099 1812 15102
rect 1868 15099 1920 15102
rect 1976 15099 2028 15102
rect 2084 15099 2136 15102
rect 2192 15099 2244 15102
rect 2300 15099 2352 15102
rect 2408 15099 2460 15102
rect 2516 15099 2568 15102
rect 2624 15099 2676 15102
rect 2732 15099 2784 15102
rect 2840 15099 2892 15102
rect 2948 15099 3000 15102
rect 3056 15099 3108 15102
rect 3164 15099 3216 15102
rect 3272 15099 3324 15102
rect 3380 15099 3432 15102
rect 3488 15099 3540 15102
rect 3596 15099 3648 15102
rect 3704 15099 3756 15102
rect 4130 15099 4182 15102
rect 4238 15099 4290 15102
rect 4346 15099 4398 15102
rect 4454 15099 4506 15102
rect 4562 15099 4614 15102
rect 4670 15099 4722 15102
rect 4778 15099 4830 15102
rect 4886 15099 4938 15102
rect 4994 15099 5046 15102
rect 5102 15099 5154 15102
rect 5210 15099 5262 15102
rect 5318 15099 5370 15102
rect 5426 15099 5478 15102
rect 5534 15099 5586 15102
rect 5642 15099 5694 15102
rect 5750 15099 5802 15102
rect 5858 15099 5910 15102
rect 5966 15099 6018 15102
rect 6074 15099 6126 15102
rect 6836 15099 6888 15102
rect 6944 15099 6996 15102
rect 7052 15099 7104 15102
rect 7160 15099 7212 15102
rect 7268 15099 7320 15102
rect 7376 15099 7428 15102
rect 7484 15099 7536 15102
rect 7592 15099 7644 15102
rect 7700 15099 7752 15102
rect 7808 15099 7860 15102
rect 7916 15099 7968 15102
rect 8024 15099 8076 15102
rect 8132 15099 8184 15102
rect 8240 15099 8292 15102
rect 8348 15099 8400 15102
rect 8456 15099 8508 15102
rect 8564 15099 8616 15102
rect 8672 15099 8724 15102
rect 8780 15099 8832 15102
rect 9206 15099 9258 15102
rect 9314 15099 9366 15102
rect 9422 15099 9474 15102
rect 9530 15099 9582 15102
rect 9638 15099 9690 15102
rect 9746 15099 9798 15102
rect 9854 15099 9906 15102
rect 9962 15099 10014 15102
rect 10070 15099 10122 15102
rect 10178 15099 10230 15102
rect 10286 15099 10338 15102
rect 10394 15099 10446 15102
rect 10502 15099 10554 15102
rect 10610 15099 10662 15102
rect 10718 15099 10770 15102
rect 10826 15099 10878 15102
rect 10934 15099 10986 15102
rect 11042 15099 11094 15102
rect 11150 15099 11202 15102
rect 1493 14904 1545 14907
rect 1601 14904 1653 14907
rect 3863 14904 3915 14907
rect 3971 14904 4023 14907
rect 6239 14904 6291 14907
rect 6347 14904 6399 14907
rect 6455 14904 6507 14907
rect 6563 14904 6615 14907
rect 6671 14904 6723 14907
rect 8939 14904 8991 14907
rect 9047 14904 9099 14907
rect 11309 14904 11361 14907
rect 11417 14904 11469 14907
rect 1493 14858 1494 14904
rect 1494 14858 1545 14904
rect 1601 14858 1653 14904
rect 3863 14858 3915 14904
rect 3971 14858 4023 14904
rect 6239 14858 6291 14904
rect 6347 14858 6399 14904
rect 6455 14858 6507 14904
rect 6563 14858 6615 14904
rect 6671 14858 6723 14904
rect 8939 14858 8991 14904
rect 9047 14858 9099 14904
rect 11309 14858 11361 14904
rect 11417 14858 11468 14904
rect 11468 14858 11469 14904
rect 1493 14855 1545 14858
rect 1601 14855 1653 14858
rect 3863 14855 3915 14858
rect 3971 14855 4023 14858
rect 6239 14855 6291 14858
rect 6347 14855 6399 14858
rect 6455 14855 6507 14858
rect 6563 14855 6615 14858
rect 6671 14855 6723 14858
rect 8939 14855 8991 14858
rect 9047 14855 9099 14858
rect 11309 14855 11361 14858
rect 11417 14855 11469 14858
rect 1760 14660 1812 14663
rect 1868 14660 1920 14663
rect 1976 14660 2028 14663
rect 2084 14660 2136 14663
rect 2192 14660 2244 14663
rect 2300 14660 2352 14663
rect 2408 14660 2460 14663
rect 2516 14660 2568 14663
rect 2624 14660 2676 14663
rect 2732 14660 2784 14663
rect 2840 14660 2892 14663
rect 2948 14660 3000 14663
rect 3056 14660 3108 14663
rect 3164 14660 3216 14663
rect 3272 14660 3324 14663
rect 3380 14660 3432 14663
rect 3488 14660 3540 14663
rect 3596 14660 3648 14663
rect 3704 14660 3756 14663
rect 4130 14660 4182 14663
rect 4238 14660 4290 14663
rect 4346 14660 4398 14663
rect 4454 14660 4506 14663
rect 4562 14660 4614 14663
rect 4670 14660 4722 14663
rect 4778 14660 4830 14663
rect 4886 14660 4938 14663
rect 4994 14660 5046 14663
rect 5102 14660 5154 14663
rect 5210 14660 5262 14663
rect 5318 14660 5370 14663
rect 5426 14660 5478 14663
rect 5534 14660 5586 14663
rect 5642 14660 5694 14663
rect 5750 14660 5802 14663
rect 5858 14660 5910 14663
rect 5966 14660 6018 14663
rect 6074 14660 6126 14663
rect 6836 14660 6888 14663
rect 6944 14660 6996 14663
rect 7052 14660 7104 14663
rect 7160 14660 7212 14663
rect 7268 14660 7320 14663
rect 7376 14660 7428 14663
rect 7484 14660 7536 14663
rect 7592 14660 7644 14663
rect 7700 14660 7752 14663
rect 7808 14660 7860 14663
rect 7916 14660 7968 14663
rect 8024 14660 8076 14663
rect 8132 14660 8184 14663
rect 8240 14660 8292 14663
rect 8348 14660 8400 14663
rect 8456 14660 8508 14663
rect 8564 14660 8616 14663
rect 8672 14660 8724 14663
rect 8780 14660 8832 14663
rect 9206 14660 9258 14663
rect 9314 14660 9366 14663
rect 9422 14660 9474 14663
rect 9530 14660 9582 14663
rect 9638 14660 9690 14663
rect 9746 14660 9798 14663
rect 9854 14660 9906 14663
rect 9962 14660 10014 14663
rect 10070 14660 10122 14663
rect 10178 14660 10230 14663
rect 10286 14660 10338 14663
rect 10394 14660 10446 14663
rect 10502 14660 10554 14663
rect 10610 14660 10662 14663
rect 10718 14660 10770 14663
rect 10826 14660 10878 14663
rect 10934 14660 10986 14663
rect 11042 14660 11094 14663
rect 11150 14660 11202 14663
rect 1760 14614 1812 14660
rect 1868 14614 1920 14660
rect 1976 14614 2028 14660
rect 2084 14614 2136 14660
rect 2192 14614 2244 14660
rect 2300 14614 2352 14660
rect 2408 14614 2460 14660
rect 2516 14614 2568 14660
rect 2624 14614 2676 14660
rect 2732 14614 2784 14660
rect 2840 14614 2892 14660
rect 2948 14614 3000 14660
rect 3056 14614 3108 14660
rect 3164 14614 3216 14660
rect 3272 14614 3324 14660
rect 3380 14614 3432 14660
rect 3488 14614 3540 14660
rect 3596 14614 3648 14660
rect 3704 14614 3756 14660
rect 4130 14614 4182 14660
rect 4238 14614 4290 14660
rect 4346 14614 4398 14660
rect 4454 14614 4506 14660
rect 4562 14614 4614 14660
rect 4670 14614 4722 14660
rect 4778 14614 4830 14660
rect 4886 14614 4938 14660
rect 4994 14614 5046 14660
rect 5102 14614 5154 14660
rect 5210 14614 5262 14660
rect 5318 14614 5370 14660
rect 5426 14614 5478 14660
rect 5534 14614 5586 14660
rect 5642 14614 5694 14660
rect 5750 14614 5802 14660
rect 5858 14614 5910 14660
rect 5966 14614 6018 14660
rect 6074 14614 6126 14660
rect 6836 14614 6888 14660
rect 6944 14614 6996 14660
rect 7052 14614 7104 14660
rect 7160 14614 7212 14660
rect 7268 14614 7320 14660
rect 7376 14614 7428 14660
rect 7484 14614 7536 14660
rect 7592 14614 7644 14660
rect 7700 14614 7752 14660
rect 7808 14614 7860 14660
rect 7916 14614 7968 14660
rect 8024 14614 8076 14660
rect 8132 14614 8184 14660
rect 8240 14614 8292 14660
rect 8348 14614 8400 14660
rect 8456 14614 8508 14660
rect 8564 14614 8616 14660
rect 8672 14614 8724 14660
rect 8780 14614 8832 14660
rect 9206 14614 9258 14660
rect 9314 14614 9366 14660
rect 9422 14614 9474 14660
rect 9530 14614 9582 14660
rect 9638 14614 9690 14660
rect 9746 14614 9798 14660
rect 9854 14614 9906 14660
rect 9962 14614 10014 14660
rect 10070 14614 10122 14660
rect 10178 14614 10230 14660
rect 10286 14614 10338 14660
rect 10394 14614 10446 14660
rect 10502 14614 10554 14660
rect 10610 14614 10662 14660
rect 10718 14614 10770 14660
rect 10826 14614 10878 14660
rect 10934 14614 10986 14660
rect 11042 14614 11094 14660
rect 11150 14614 11202 14660
rect 1760 14611 1812 14614
rect 1868 14611 1920 14614
rect 1976 14611 2028 14614
rect 2084 14611 2136 14614
rect 2192 14611 2244 14614
rect 2300 14611 2352 14614
rect 2408 14611 2460 14614
rect 2516 14611 2568 14614
rect 2624 14611 2676 14614
rect 2732 14611 2784 14614
rect 2840 14611 2892 14614
rect 2948 14611 3000 14614
rect 3056 14611 3108 14614
rect 3164 14611 3216 14614
rect 3272 14611 3324 14614
rect 3380 14611 3432 14614
rect 3488 14611 3540 14614
rect 3596 14611 3648 14614
rect 3704 14611 3756 14614
rect 4130 14611 4182 14614
rect 4238 14611 4290 14614
rect 4346 14611 4398 14614
rect 4454 14611 4506 14614
rect 4562 14611 4614 14614
rect 4670 14611 4722 14614
rect 4778 14611 4830 14614
rect 4886 14611 4938 14614
rect 4994 14611 5046 14614
rect 5102 14611 5154 14614
rect 5210 14611 5262 14614
rect 5318 14611 5370 14614
rect 5426 14611 5478 14614
rect 5534 14611 5586 14614
rect 5642 14611 5694 14614
rect 5750 14611 5802 14614
rect 5858 14611 5910 14614
rect 5966 14611 6018 14614
rect 6074 14611 6126 14614
rect 6836 14611 6888 14614
rect 6944 14611 6996 14614
rect 7052 14611 7104 14614
rect 7160 14611 7212 14614
rect 7268 14611 7320 14614
rect 7376 14611 7428 14614
rect 7484 14611 7536 14614
rect 7592 14611 7644 14614
rect 7700 14611 7752 14614
rect 7808 14611 7860 14614
rect 7916 14611 7968 14614
rect 8024 14611 8076 14614
rect 8132 14611 8184 14614
rect 8240 14611 8292 14614
rect 8348 14611 8400 14614
rect 8456 14611 8508 14614
rect 8564 14611 8616 14614
rect 8672 14611 8724 14614
rect 8780 14611 8832 14614
rect 9206 14611 9258 14614
rect 9314 14611 9366 14614
rect 9422 14611 9474 14614
rect 9530 14611 9582 14614
rect 9638 14611 9690 14614
rect 9746 14611 9798 14614
rect 9854 14611 9906 14614
rect 9962 14611 10014 14614
rect 10070 14611 10122 14614
rect 10178 14611 10230 14614
rect 10286 14611 10338 14614
rect 10394 14611 10446 14614
rect 10502 14611 10554 14614
rect 10610 14611 10662 14614
rect 10718 14611 10770 14614
rect 10826 14611 10878 14614
rect 10934 14611 10986 14614
rect 11042 14611 11094 14614
rect 11150 14611 11202 14614
rect 1493 14416 1545 14419
rect 1601 14416 1653 14419
rect 3863 14416 3915 14419
rect 3971 14416 4023 14419
rect 6239 14416 6291 14419
rect 6347 14416 6399 14419
rect 6455 14416 6507 14419
rect 6563 14416 6615 14419
rect 6671 14416 6723 14419
rect 8939 14416 8991 14419
rect 9047 14416 9099 14419
rect 11309 14416 11361 14419
rect 11417 14416 11469 14419
rect 1493 14370 1494 14416
rect 1494 14370 1545 14416
rect 1601 14370 1653 14416
rect 3863 14370 3915 14416
rect 3971 14370 4023 14416
rect 6239 14370 6291 14416
rect 6347 14370 6399 14416
rect 6455 14370 6507 14416
rect 6563 14370 6615 14416
rect 6671 14370 6723 14416
rect 8939 14370 8991 14416
rect 9047 14370 9099 14416
rect 11309 14370 11361 14416
rect 11417 14370 11468 14416
rect 11468 14370 11469 14416
rect 1493 14367 1545 14370
rect 1601 14367 1653 14370
rect 3863 14367 3915 14370
rect 3971 14367 4023 14370
rect 6239 14367 6291 14370
rect 6347 14367 6399 14370
rect 6455 14367 6507 14370
rect 6563 14367 6615 14370
rect 6671 14367 6723 14370
rect 8939 14367 8991 14370
rect 9047 14367 9099 14370
rect 11309 14367 11361 14370
rect 11417 14367 11469 14370
rect 1760 14172 1812 14175
rect 1868 14172 1920 14175
rect 1976 14172 2028 14175
rect 2084 14172 2136 14175
rect 2192 14172 2244 14175
rect 2300 14172 2352 14175
rect 2408 14172 2460 14175
rect 2516 14172 2568 14175
rect 2624 14172 2676 14175
rect 2732 14172 2784 14175
rect 2840 14172 2892 14175
rect 2948 14172 3000 14175
rect 3056 14172 3108 14175
rect 3164 14172 3216 14175
rect 3272 14172 3324 14175
rect 3380 14172 3432 14175
rect 3488 14172 3540 14175
rect 3596 14172 3648 14175
rect 3704 14172 3756 14175
rect 4130 14172 4182 14175
rect 4238 14172 4290 14175
rect 4346 14172 4398 14175
rect 4454 14172 4506 14175
rect 4562 14172 4614 14175
rect 4670 14172 4722 14175
rect 4778 14172 4830 14175
rect 4886 14172 4938 14175
rect 4994 14172 5046 14175
rect 5102 14172 5154 14175
rect 5210 14172 5262 14175
rect 5318 14172 5370 14175
rect 5426 14172 5478 14175
rect 5534 14172 5586 14175
rect 5642 14172 5694 14175
rect 5750 14172 5802 14175
rect 5858 14172 5910 14175
rect 5966 14172 6018 14175
rect 6074 14172 6126 14175
rect 6836 14172 6888 14175
rect 6944 14172 6996 14175
rect 7052 14172 7104 14175
rect 7160 14172 7212 14175
rect 7268 14172 7320 14175
rect 7376 14172 7428 14175
rect 7484 14172 7536 14175
rect 7592 14172 7644 14175
rect 7700 14172 7752 14175
rect 7808 14172 7860 14175
rect 7916 14172 7968 14175
rect 8024 14172 8076 14175
rect 8132 14172 8184 14175
rect 8240 14172 8292 14175
rect 8348 14172 8400 14175
rect 8456 14172 8508 14175
rect 8564 14172 8616 14175
rect 8672 14172 8724 14175
rect 8780 14172 8832 14175
rect 9206 14172 9258 14175
rect 9314 14172 9366 14175
rect 9422 14172 9474 14175
rect 9530 14172 9582 14175
rect 9638 14172 9690 14175
rect 9746 14172 9798 14175
rect 9854 14172 9906 14175
rect 9962 14172 10014 14175
rect 10070 14172 10122 14175
rect 10178 14172 10230 14175
rect 10286 14172 10338 14175
rect 10394 14172 10446 14175
rect 10502 14172 10554 14175
rect 10610 14172 10662 14175
rect 10718 14172 10770 14175
rect 10826 14172 10878 14175
rect 10934 14172 10986 14175
rect 11042 14172 11094 14175
rect 11150 14172 11202 14175
rect 1760 14126 1812 14172
rect 1868 14126 1920 14172
rect 1976 14126 2028 14172
rect 2084 14126 2136 14172
rect 2192 14126 2244 14172
rect 2300 14126 2352 14172
rect 2408 14126 2460 14172
rect 2516 14126 2568 14172
rect 2624 14126 2676 14172
rect 2732 14126 2784 14172
rect 2840 14126 2892 14172
rect 2948 14126 3000 14172
rect 3056 14126 3108 14172
rect 3164 14126 3216 14172
rect 3272 14126 3324 14172
rect 3380 14126 3432 14172
rect 3488 14126 3540 14172
rect 3596 14126 3648 14172
rect 3704 14126 3756 14172
rect 4130 14126 4182 14172
rect 4238 14126 4290 14172
rect 4346 14126 4398 14172
rect 4454 14126 4506 14172
rect 4562 14126 4614 14172
rect 4670 14126 4722 14172
rect 4778 14126 4830 14172
rect 4886 14126 4938 14172
rect 4994 14126 5046 14172
rect 5102 14126 5154 14172
rect 5210 14126 5262 14172
rect 5318 14126 5370 14172
rect 5426 14126 5478 14172
rect 5534 14126 5586 14172
rect 5642 14126 5694 14172
rect 5750 14126 5802 14172
rect 5858 14126 5910 14172
rect 5966 14126 6018 14172
rect 6074 14126 6126 14172
rect 6836 14126 6888 14172
rect 6944 14126 6996 14172
rect 7052 14126 7104 14172
rect 7160 14126 7212 14172
rect 7268 14126 7320 14172
rect 7376 14126 7428 14172
rect 7484 14126 7536 14172
rect 7592 14126 7644 14172
rect 7700 14126 7752 14172
rect 7808 14126 7860 14172
rect 7916 14126 7968 14172
rect 8024 14126 8076 14172
rect 8132 14126 8184 14172
rect 8240 14126 8292 14172
rect 8348 14126 8400 14172
rect 8456 14126 8508 14172
rect 8564 14126 8616 14172
rect 8672 14126 8724 14172
rect 8780 14126 8832 14172
rect 9206 14126 9258 14172
rect 9314 14126 9366 14172
rect 9422 14126 9474 14172
rect 9530 14126 9582 14172
rect 9638 14126 9690 14172
rect 9746 14126 9798 14172
rect 9854 14126 9906 14172
rect 9962 14126 10014 14172
rect 10070 14126 10122 14172
rect 10178 14126 10230 14172
rect 10286 14126 10338 14172
rect 10394 14126 10446 14172
rect 10502 14126 10554 14172
rect 10610 14126 10662 14172
rect 10718 14126 10770 14172
rect 10826 14126 10878 14172
rect 10934 14126 10986 14172
rect 11042 14126 11094 14172
rect 11150 14126 11202 14172
rect 1760 14123 1812 14126
rect 1868 14123 1920 14126
rect 1976 14123 2028 14126
rect 2084 14123 2136 14126
rect 2192 14123 2244 14126
rect 2300 14123 2352 14126
rect 2408 14123 2460 14126
rect 2516 14123 2568 14126
rect 2624 14123 2676 14126
rect 2732 14123 2784 14126
rect 2840 14123 2892 14126
rect 2948 14123 3000 14126
rect 3056 14123 3108 14126
rect 3164 14123 3216 14126
rect 3272 14123 3324 14126
rect 3380 14123 3432 14126
rect 3488 14123 3540 14126
rect 3596 14123 3648 14126
rect 3704 14123 3756 14126
rect 4130 14123 4182 14126
rect 4238 14123 4290 14126
rect 4346 14123 4398 14126
rect 4454 14123 4506 14126
rect 4562 14123 4614 14126
rect 4670 14123 4722 14126
rect 4778 14123 4830 14126
rect 4886 14123 4938 14126
rect 4994 14123 5046 14126
rect 5102 14123 5154 14126
rect 5210 14123 5262 14126
rect 5318 14123 5370 14126
rect 5426 14123 5478 14126
rect 5534 14123 5586 14126
rect 5642 14123 5694 14126
rect 5750 14123 5802 14126
rect 5858 14123 5910 14126
rect 5966 14123 6018 14126
rect 6074 14123 6126 14126
rect 6836 14123 6888 14126
rect 6944 14123 6996 14126
rect 7052 14123 7104 14126
rect 7160 14123 7212 14126
rect 7268 14123 7320 14126
rect 7376 14123 7428 14126
rect 7484 14123 7536 14126
rect 7592 14123 7644 14126
rect 7700 14123 7752 14126
rect 7808 14123 7860 14126
rect 7916 14123 7968 14126
rect 8024 14123 8076 14126
rect 8132 14123 8184 14126
rect 8240 14123 8292 14126
rect 8348 14123 8400 14126
rect 8456 14123 8508 14126
rect 8564 14123 8616 14126
rect 8672 14123 8724 14126
rect 8780 14123 8832 14126
rect 9206 14123 9258 14126
rect 9314 14123 9366 14126
rect 9422 14123 9474 14126
rect 9530 14123 9582 14126
rect 9638 14123 9690 14126
rect 9746 14123 9798 14126
rect 9854 14123 9906 14126
rect 9962 14123 10014 14126
rect 10070 14123 10122 14126
rect 10178 14123 10230 14126
rect 10286 14123 10338 14126
rect 10394 14123 10446 14126
rect 10502 14123 10554 14126
rect 10610 14123 10662 14126
rect 10718 14123 10770 14126
rect 10826 14123 10878 14126
rect 10934 14123 10986 14126
rect 11042 14123 11094 14126
rect 11150 14123 11202 14126
rect 1493 13928 1545 13931
rect 1601 13928 1653 13931
rect 3863 13928 3915 13931
rect 3971 13928 4023 13931
rect 6239 13928 6291 13931
rect 6347 13928 6399 13931
rect 6455 13928 6507 13931
rect 6563 13928 6615 13931
rect 6671 13928 6723 13931
rect 8939 13928 8991 13931
rect 9047 13928 9099 13931
rect 11309 13928 11361 13931
rect 11417 13928 11469 13931
rect 1493 13882 1494 13928
rect 1494 13882 1545 13928
rect 1601 13882 1653 13928
rect 3863 13882 3915 13928
rect 3971 13882 4023 13928
rect 6239 13882 6291 13928
rect 6347 13882 6399 13928
rect 6455 13882 6507 13928
rect 6563 13882 6615 13928
rect 6671 13882 6723 13928
rect 8939 13882 8991 13928
rect 9047 13882 9099 13928
rect 11309 13882 11361 13928
rect 11417 13882 11468 13928
rect 11468 13882 11469 13928
rect 1493 13879 1545 13882
rect 1601 13879 1653 13882
rect 3863 13879 3915 13882
rect 3971 13879 4023 13882
rect 6239 13879 6291 13882
rect 6347 13879 6399 13882
rect 6455 13879 6507 13882
rect 6563 13879 6615 13882
rect 6671 13879 6723 13882
rect 8939 13879 8991 13882
rect 9047 13879 9099 13882
rect 11309 13879 11361 13882
rect 11417 13879 11469 13882
rect 1760 13684 1812 13687
rect 1868 13684 1920 13687
rect 1976 13684 2028 13687
rect 2084 13684 2136 13687
rect 2192 13684 2244 13687
rect 2300 13684 2352 13687
rect 2408 13684 2460 13687
rect 2516 13684 2568 13687
rect 2624 13684 2676 13687
rect 2732 13684 2784 13687
rect 2840 13684 2892 13687
rect 2948 13684 3000 13687
rect 3056 13684 3108 13687
rect 3164 13684 3216 13687
rect 3272 13684 3324 13687
rect 3380 13684 3432 13687
rect 3488 13684 3540 13687
rect 3596 13684 3648 13687
rect 3704 13684 3756 13687
rect 4130 13684 4182 13687
rect 4238 13684 4290 13687
rect 4346 13684 4398 13687
rect 4454 13684 4506 13687
rect 4562 13684 4614 13687
rect 4670 13684 4722 13687
rect 4778 13684 4830 13687
rect 4886 13684 4938 13687
rect 4994 13684 5046 13687
rect 5102 13684 5154 13687
rect 5210 13684 5262 13687
rect 5318 13684 5370 13687
rect 5426 13684 5478 13687
rect 5534 13684 5586 13687
rect 5642 13684 5694 13687
rect 5750 13684 5802 13687
rect 5858 13684 5910 13687
rect 5966 13684 6018 13687
rect 6074 13684 6126 13687
rect 6836 13684 6888 13687
rect 6944 13684 6996 13687
rect 7052 13684 7104 13687
rect 7160 13684 7212 13687
rect 7268 13684 7320 13687
rect 7376 13684 7428 13687
rect 7484 13684 7536 13687
rect 7592 13684 7644 13687
rect 7700 13684 7752 13687
rect 7808 13684 7860 13687
rect 7916 13684 7968 13687
rect 8024 13684 8076 13687
rect 8132 13684 8184 13687
rect 8240 13684 8292 13687
rect 8348 13684 8400 13687
rect 8456 13684 8508 13687
rect 8564 13684 8616 13687
rect 8672 13684 8724 13687
rect 8780 13684 8832 13687
rect 9206 13684 9258 13687
rect 9314 13684 9366 13687
rect 9422 13684 9474 13687
rect 9530 13684 9582 13687
rect 9638 13684 9690 13687
rect 9746 13684 9798 13687
rect 9854 13684 9906 13687
rect 9962 13684 10014 13687
rect 10070 13684 10122 13687
rect 10178 13684 10230 13687
rect 10286 13684 10338 13687
rect 10394 13684 10446 13687
rect 10502 13684 10554 13687
rect 10610 13684 10662 13687
rect 10718 13684 10770 13687
rect 10826 13684 10878 13687
rect 10934 13684 10986 13687
rect 11042 13684 11094 13687
rect 11150 13684 11202 13687
rect 1760 13638 1812 13684
rect 1868 13638 1920 13684
rect 1976 13638 2028 13684
rect 2084 13638 2136 13684
rect 2192 13638 2244 13684
rect 2300 13638 2352 13684
rect 2408 13638 2460 13684
rect 2516 13638 2568 13684
rect 2624 13638 2676 13684
rect 2732 13638 2784 13684
rect 2840 13638 2892 13684
rect 2948 13638 3000 13684
rect 3056 13638 3108 13684
rect 3164 13638 3216 13684
rect 3272 13638 3324 13684
rect 3380 13638 3432 13684
rect 3488 13638 3540 13684
rect 3596 13638 3648 13684
rect 3704 13638 3756 13684
rect 4130 13638 4182 13684
rect 4238 13638 4290 13684
rect 4346 13638 4398 13684
rect 4454 13638 4506 13684
rect 4562 13638 4614 13684
rect 4670 13638 4722 13684
rect 4778 13638 4830 13684
rect 4886 13638 4938 13684
rect 4994 13638 5046 13684
rect 5102 13638 5154 13684
rect 5210 13638 5262 13684
rect 5318 13638 5370 13684
rect 5426 13638 5478 13684
rect 5534 13638 5586 13684
rect 5642 13638 5694 13684
rect 5750 13638 5802 13684
rect 5858 13638 5910 13684
rect 5966 13638 6018 13684
rect 6074 13638 6126 13684
rect 6836 13638 6888 13684
rect 6944 13638 6996 13684
rect 7052 13638 7104 13684
rect 7160 13638 7212 13684
rect 7268 13638 7320 13684
rect 7376 13638 7428 13684
rect 7484 13638 7536 13684
rect 7592 13638 7644 13684
rect 7700 13638 7752 13684
rect 7808 13638 7860 13684
rect 7916 13638 7968 13684
rect 8024 13638 8076 13684
rect 8132 13638 8184 13684
rect 8240 13638 8292 13684
rect 8348 13638 8400 13684
rect 8456 13638 8508 13684
rect 8564 13638 8616 13684
rect 8672 13638 8724 13684
rect 8780 13638 8832 13684
rect 9206 13638 9258 13684
rect 9314 13638 9366 13684
rect 9422 13638 9474 13684
rect 9530 13638 9582 13684
rect 9638 13638 9690 13684
rect 9746 13638 9798 13684
rect 9854 13638 9906 13684
rect 9962 13638 10014 13684
rect 10070 13638 10122 13684
rect 10178 13638 10230 13684
rect 10286 13638 10338 13684
rect 10394 13638 10446 13684
rect 10502 13638 10554 13684
rect 10610 13638 10662 13684
rect 10718 13638 10770 13684
rect 10826 13638 10878 13684
rect 10934 13638 10986 13684
rect 11042 13638 11094 13684
rect 11150 13638 11202 13684
rect 1760 13635 1812 13638
rect 1868 13635 1920 13638
rect 1976 13635 2028 13638
rect 2084 13635 2136 13638
rect 2192 13635 2244 13638
rect 2300 13635 2352 13638
rect 2408 13635 2460 13638
rect 2516 13635 2568 13638
rect 2624 13635 2676 13638
rect 2732 13635 2784 13638
rect 2840 13635 2892 13638
rect 2948 13635 3000 13638
rect 3056 13635 3108 13638
rect 3164 13635 3216 13638
rect 3272 13635 3324 13638
rect 3380 13635 3432 13638
rect 3488 13635 3540 13638
rect 3596 13635 3648 13638
rect 3704 13635 3756 13638
rect 4130 13635 4182 13638
rect 4238 13635 4290 13638
rect 4346 13635 4398 13638
rect 4454 13635 4506 13638
rect 4562 13635 4614 13638
rect 4670 13635 4722 13638
rect 4778 13635 4830 13638
rect 4886 13635 4938 13638
rect 4994 13635 5046 13638
rect 5102 13635 5154 13638
rect 5210 13635 5262 13638
rect 5318 13635 5370 13638
rect 5426 13635 5478 13638
rect 5534 13635 5586 13638
rect 5642 13635 5694 13638
rect 5750 13635 5802 13638
rect 5858 13635 5910 13638
rect 5966 13635 6018 13638
rect 6074 13635 6126 13638
rect 6836 13635 6888 13638
rect 6944 13635 6996 13638
rect 7052 13635 7104 13638
rect 7160 13635 7212 13638
rect 7268 13635 7320 13638
rect 7376 13635 7428 13638
rect 7484 13635 7536 13638
rect 7592 13635 7644 13638
rect 7700 13635 7752 13638
rect 7808 13635 7860 13638
rect 7916 13635 7968 13638
rect 8024 13635 8076 13638
rect 8132 13635 8184 13638
rect 8240 13635 8292 13638
rect 8348 13635 8400 13638
rect 8456 13635 8508 13638
rect 8564 13635 8616 13638
rect 8672 13635 8724 13638
rect 8780 13635 8832 13638
rect 9206 13635 9258 13638
rect 9314 13635 9366 13638
rect 9422 13635 9474 13638
rect 9530 13635 9582 13638
rect 9638 13635 9690 13638
rect 9746 13635 9798 13638
rect 9854 13635 9906 13638
rect 9962 13635 10014 13638
rect 10070 13635 10122 13638
rect 10178 13635 10230 13638
rect 10286 13635 10338 13638
rect 10394 13635 10446 13638
rect 10502 13635 10554 13638
rect 10610 13635 10662 13638
rect 10718 13635 10770 13638
rect 10826 13635 10878 13638
rect 10934 13635 10986 13638
rect 11042 13635 11094 13638
rect 11150 13635 11202 13638
rect 1493 13440 1545 13443
rect 1601 13440 1653 13443
rect 3863 13440 3915 13443
rect 3971 13440 4023 13443
rect 6239 13440 6291 13443
rect 6347 13440 6399 13443
rect 6455 13440 6507 13443
rect 6563 13440 6615 13443
rect 6671 13440 6723 13443
rect 8939 13440 8991 13443
rect 9047 13440 9099 13443
rect 11309 13440 11361 13443
rect 11417 13440 11469 13443
rect 1493 13394 1494 13440
rect 1494 13394 1545 13440
rect 1601 13394 1653 13440
rect 3863 13394 3915 13440
rect 3971 13394 4023 13440
rect 6239 13394 6291 13440
rect 6347 13394 6399 13440
rect 6455 13394 6507 13440
rect 6563 13394 6615 13440
rect 6671 13394 6723 13440
rect 8939 13394 8991 13440
rect 9047 13394 9099 13440
rect 11309 13394 11361 13440
rect 11417 13394 11468 13440
rect 11468 13394 11469 13440
rect 1493 13391 1545 13394
rect 1601 13391 1653 13394
rect 3863 13391 3915 13394
rect 3971 13391 4023 13394
rect 6239 13391 6291 13394
rect 6347 13391 6399 13394
rect 6455 13391 6507 13394
rect 6563 13391 6615 13394
rect 6671 13391 6723 13394
rect 8939 13391 8991 13394
rect 9047 13391 9099 13394
rect 11309 13391 11361 13394
rect 11417 13391 11469 13394
rect 1233 13211 1285 13263
rect 1341 13211 1393 13263
rect 11569 17855 11621 17907
rect 11677 17855 11706 17907
rect 11706 17855 11729 17907
rect 11569 17747 11621 17799
rect 11677 17747 11706 17799
rect 11706 17747 11729 17799
rect 11569 17639 11621 17691
rect 11677 17639 11706 17691
rect 11706 17639 11729 17691
rect 11569 17531 11621 17583
rect 11677 17531 11706 17583
rect 11706 17531 11729 17583
rect 11569 17423 11621 17475
rect 11677 17423 11706 17475
rect 11706 17423 11729 17475
rect 11569 17315 11621 17367
rect 11677 17315 11706 17367
rect 11706 17315 11729 17367
rect 11569 17207 11621 17259
rect 11677 17207 11706 17259
rect 11706 17207 11729 17259
rect 11569 17099 11621 17151
rect 11677 17099 11706 17151
rect 11706 17099 11729 17151
rect 11569 16991 11621 17043
rect 11677 16991 11706 17043
rect 11706 16991 11729 17043
rect 11569 16883 11621 16935
rect 11677 16883 11706 16935
rect 11706 16883 11729 16935
rect 11569 16775 11621 16827
rect 11677 16775 11706 16827
rect 11706 16775 11729 16827
rect 11569 16667 11621 16719
rect 11677 16667 11706 16719
rect 11706 16667 11729 16719
rect 11569 16559 11621 16611
rect 11677 16559 11706 16611
rect 11706 16559 11729 16611
rect 11569 16451 11621 16503
rect 11677 16451 11706 16503
rect 11706 16451 11729 16503
rect 11569 16343 11621 16395
rect 11677 16343 11706 16395
rect 11706 16343 11729 16395
rect 11569 16235 11621 16287
rect 11677 16235 11706 16287
rect 11706 16235 11729 16287
rect 11569 16127 11621 16179
rect 11677 16127 11706 16179
rect 11706 16127 11729 16179
rect 11569 16019 11621 16071
rect 11677 16019 11706 16071
rect 11706 16019 11729 16071
rect 11569 15911 11621 15963
rect 11677 15911 11706 15963
rect 11706 15911 11729 15963
rect 11569 15803 11621 15855
rect 11677 15803 11706 15855
rect 11706 15803 11729 15855
rect 11569 15695 11621 15747
rect 11677 15695 11706 15747
rect 11706 15695 11729 15747
rect 11569 15587 11621 15639
rect 11677 15587 11706 15639
rect 11706 15587 11729 15639
rect 11569 15479 11621 15531
rect 11677 15479 11706 15531
rect 11706 15479 11729 15531
rect 11569 15371 11621 15423
rect 11677 15371 11706 15423
rect 11706 15371 11729 15423
rect 11569 15263 11621 15315
rect 11677 15263 11706 15315
rect 11706 15263 11729 15315
rect 11569 15155 11621 15207
rect 11677 15155 11706 15207
rect 11706 15155 11729 15207
rect 11569 15047 11621 15099
rect 11677 15047 11706 15099
rect 11706 15047 11729 15099
rect 11569 14939 11621 14991
rect 11677 14939 11706 14991
rect 11706 14939 11729 14991
rect 11569 14831 11621 14883
rect 11677 14831 11706 14883
rect 11706 14831 11729 14883
rect 11569 14723 11621 14775
rect 11677 14723 11706 14775
rect 11706 14723 11729 14775
rect 11569 14615 11621 14667
rect 11677 14615 11706 14667
rect 11706 14615 11729 14667
rect 11569 14507 11621 14559
rect 11677 14507 11706 14559
rect 11706 14507 11729 14559
rect 11569 14399 11621 14451
rect 11677 14399 11706 14451
rect 11706 14399 11729 14451
rect 11569 14291 11621 14343
rect 11677 14291 11706 14343
rect 11706 14291 11729 14343
rect 11569 14183 11621 14235
rect 11677 14183 11706 14235
rect 11706 14183 11729 14235
rect 11569 14075 11621 14127
rect 11677 14075 11706 14127
rect 11706 14075 11729 14127
rect 11569 13967 11621 14019
rect 11677 13967 11706 14019
rect 11706 13967 11729 14019
rect 11569 13859 11621 13911
rect 11677 13859 11706 13911
rect 11706 13859 11729 13911
rect 11569 13751 11621 13803
rect 11677 13751 11706 13803
rect 11706 13751 11729 13803
rect 11569 13643 11621 13695
rect 11677 13643 11706 13695
rect 11706 13643 11729 13695
rect 11569 13535 11621 13587
rect 11677 13535 11706 13587
rect 11706 13535 11729 13587
rect 11569 13427 11621 13479
rect 11677 13427 11706 13479
rect 11706 13427 11729 13479
rect 11569 13319 11621 13371
rect 11677 13319 11706 13371
rect 11706 13319 11729 13371
rect 11569 13211 11621 13263
rect 11677 13211 11729 13263
rect 1760 13196 1812 13199
rect 1868 13196 1920 13199
rect 1976 13196 2028 13199
rect 2084 13196 2136 13199
rect 2192 13196 2244 13199
rect 2300 13196 2352 13199
rect 2408 13196 2460 13199
rect 2516 13196 2568 13199
rect 2624 13196 2676 13199
rect 2732 13196 2784 13199
rect 2840 13196 2892 13199
rect 2948 13196 3000 13199
rect 3056 13196 3108 13199
rect 3164 13196 3216 13199
rect 3272 13196 3324 13199
rect 3380 13196 3432 13199
rect 3488 13196 3540 13199
rect 3596 13196 3648 13199
rect 3704 13196 3756 13199
rect 4130 13196 4182 13199
rect 4238 13196 4290 13199
rect 4346 13196 4398 13199
rect 4454 13196 4506 13199
rect 4562 13196 4614 13199
rect 4670 13196 4722 13199
rect 4778 13196 4830 13199
rect 4886 13196 4938 13199
rect 4994 13196 5046 13199
rect 5102 13196 5154 13199
rect 5210 13196 5262 13199
rect 5318 13196 5370 13199
rect 5426 13196 5478 13199
rect 5534 13196 5586 13199
rect 5642 13196 5694 13199
rect 5750 13196 5802 13199
rect 5858 13196 5910 13199
rect 5966 13196 6018 13199
rect 6074 13196 6126 13199
rect 6836 13196 6888 13199
rect 6944 13196 6996 13199
rect 7052 13196 7104 13199
rect 7160 13196 7212 13199
rect 7268 13196 7320 13199
rect 7376 13196 7428 13199
rect 7484 13196 7536 13199
rect 7592 13196 7644 13199
rect 7700 13196 7752 13199
rect 7808 13196 7860 13199
rect 7916 13196 7968 13199
rect 8024 13196 8076 13199
rect 8132 13196 8184 13199
rect 8240 13196 8292 13199
rect 8348 13196 8400 13199
rect 8456 13196 8508 13199
rect 8564 13196 8616 13199
rect 8672 13196 8724 13199
rect 8780 13196 8832 13199
rect 9206 13196 9258 13199
rect 9314 13196 9366 13199
rect 9422 13196 9474 13199
rect 9530 13196 9582 13199
rect 9638 13196 9690 13199
rect 9746 13196 9798 13199
rect 9854 13196 9906 13199
rect 9962 13196 10014 13199
rect 10070 13196 10122 13199
rect 10178 13196 10230 13199
rect 10286 13196 10338 13199
rect 10394 13196 10446 13199
rect 10502 13196 10554 13199
rect 10610 13196 10662 13199
rect 10718 13196 10770 13199
rect 10826 13196 10878 13199
rect 10934 13196 10986 13199
rect 11042 13196 11094 13199
rect 11150 13196 11202 13199
rect 1760 13150 1812 13196
rect 1868 13150 1920 13196
rect 1976 13150 2028 13196
rect 2084 13150 2136 13196
rect 2192 13150 2244 13196
rect 2300 13150 2352 13196
rect 2408 13150 2460 13196
rect 2516 13150 2568 13196
rect 2624 13150 2676 13196
rect 2732 13150 2784 13196
rect 2840 13150 2892 13196
rect 2948 13150 3000 13196
rect 3056 13150 3108 13196
rect 3164 13150 3216 13196
rect 3272 13150 3324 13196
rect 3380 13150 3432 13196
rect 3488 13150 3540 13196
rect 3596 13150 3648 13196
rect 3704 13150 3756 13196
rect 4130 13150 4182 13196
rect 4238 13150 4290 13196
rect 4346 13150 4398 13196
rect 4454 13150 4506 13196
rect 4562 13150 4614 13196
rect 4670 13150 4722 13196
rect 4778 13150 4830 13196
rect 4886 13150 4938 13196
rect 4994 13150 5046 13196
rect 5102 13150 5154 13196
rect 5210 13150 5262 13196
rect 5318 13150 5370 13196
rect 5426 13150 5478 13196
rect 5534 13150 5586 13196
rect 5642 13150 5694 13196
rect 5750 13150 5802 13196
rect 5858 13150 5910 13196
rect 5966 13150 6018 13196
rect 6074 13150 6126 13196
rect 6836 13150 6888 13196
rect 6944 13150 6996 13196
rect 7052 13150 7104 13196
rect 7160 13150 7212 13196
rect 7268 13150 7320 13196
rect 7376 13150 7428 13196
rect 7484 13150 7536 13196
rect 7592 13150 7644 13196
rect 7700 13150 7752 13196
rect 7808 13150 7860 13196
rect 7916 13150 7968 13196
rect 8024 13150 8076 13196
rect 8132 13150 8184 13196
rect 8240 13150 8292 13196
rect 8348 13150 8400 13196
rect 8456 13150 8508 13196
rect 8564 13150 8616 13196
rect 8672 13150 8724 13196
rect 8780 13150 8832 13196
rect 9206 13150 9258 13196
rect 9314 13150 9366 13196
rect 9422 13150 9474 13196
rect 9530 13150 9582 13196
rect 9638 13150 9690 13196
rect 9746 13150 9798 13196
rect 9854 13150 9906 13196
rect 9962 13150 10014 13196
rect 10070 13150 10122 13196
rect 10178 13150 10230 13196
rect 10286 13150 10338 13196
rect 10394 13150 10446 13196
rect 10502 13150 10554 13196
rect 10610 13150 10662 13196
rect 10718 13150 10770 13196
rect 10826 13150 10878 13196
rect 10934 13150 10986 13196
rect 11042 13150 11094 13196
rect 11150 13150 11202 13196
rect 1760 13147 1812 13150
rect 1868 13147 1920 13150
rect 1976 13147 2028 13150
rect 2084 13147 2136 13150
rect 2192 13147 2244 13150
rect 2300 13147 2352 13150
rect 2408 13147 2460 13150
rect 2516 13147 2568 13150
rect 2624 13147 2676 13150
rect 2732 13147 2784 13150
rect 2840 13147 2892 13150
rect 2948 13147 3000 13150
rect 3056 13147 3108 13150
rect 3164 13147 3216 13150
rect 3272 13147 3324 13150
rect 3380 13147 3432 13150
rect 3488 13147 3540 13150
rect 3596 13147 3648 13150
rect 3704 13147 3756 13150
rect 4130 13147 4182 13150
rect 4238 13147 4290 13150
rect 4346 13147 4398 13150
rect 4454 13147 4506 13150
rect 4562 13147 4614 13150
rect 4670 13147 4722 13150
rect 4778 13147 4830 13150
rect 4886 13147 4938 13150
rect 4994 13147 5046 13150
rect 5102 13147 5154 13150
rect 5210 13147 5262 13150
rect 5318 13147 5370 13150
rect 5426 13147 5478 13150
rect 5534 13147 5586 13150
rect 5642 13147 5694 13150
rect 5750 13147 5802 13150
rect 5858 13147 5910 13150
rect 5966 13147 6018 13150
rect 6074 13147 6126 13150
rect 6836 13147 6888 13150
rect 6944 13147 6996 13150
rect 7052 13147 7104 13150
rect 7160 13147 7212 13150
rect 7268 13147 7320 13150
rect 7376 13147 7428 13150
rect 7484 13147 7536 13150
rect 7592 13147 7644 13150
rect 7700 13147 7752 13150
rect 7808 13147 7860 13150
rect 7916 13147 7968 13150
rect 8024 13147 8076 13150
rect 8132 13147 8184 13150
rect 8240 13147 8292 13150
rect 8348 13147 8400 13150
rect 8456 13147 8508 13150
rect 8564 13147 8616 13150
rect 8672 13147 8724 13150
rect 8780 13147 8832 13150
rect 9206 13147 9258 13150
rect 9314 13147 9366 13150
rect 9422 13147 9474 13150
rect 9530 13147 9582 13150
rect 9638 13147 9690 13150
rect 9746 13147 9798 13150
rect 9854 13147 9906 13150
rect 9962 13147 10014 13150
rect 10070 13147 10122 13150
rect 10178 13147 10230 13150
rect 10286 13147 10338 13150
rect 10394 13147 10446 13150
rect 10502 13147 10554 13150
rect 10610 13147 10662 13150
rect 10718 13147 10770 13150
rect 10826 13147 10878 13150
rect 10934 13147 10986 13150
rect 11042 13147 11094 13150
rect 11150 13147 11202 13150
rect 12051 18375 12103 18427
rect 12159 18375 12211 18427
rect 12267 18375 12319 18427
rect 12051 18267 12103 18319
rect 12159 18267 12211 18319
rect 12267 18267 12319 18319
rect 12051 18159 12103 18211
rect 12159 18159 12211 18211
rect 12267 18159 12319 18211
rect 12051 18051 12103 18103
rect 12159 18051 12211 18103
rect 12267 18051 12319 18103
rect 12051 17943 12103 17995
rect 12159 17943 12211 17995
rect 12267 17943 12319 17995
rect 12051 17835 12103 17887
rect 12159 17835 12211 17887
rect 12267 17835 12319 17887
rect 12051 17727 12103 17779
rect 12159 17727 12211 17779
rect 12267 17727 12319 17779
rect 12051 17619 12103 17671
rect 12159 17619 12211 17671
rect 12267 17619 12319 17671
rect 12051 17511 12103 17563
rect 12159 17511 12211 17563
rect 12267 17511 12319 17563
rect 12051 17403 12103 17455
rect 12159 17403 12211 17455
rect 12267 17403 12319 17455
rect 12051 17295 12103 17347
rect 12159 17295 12211 17347
rect 12267 17295 12319 17347
rect 12051 17187 12103 17239
rect 12159 17187 12211 17239
rect 12267 17187 12319 17239
rect 12051 17079 12103 17131
rect 12159 17079 12211 17131
rect 12267 17079 12319 17131
rect 12051 16971 12103 17023
rect 12159 16971 12211 17023
rect 12267 16971 12319 17023
rect 12051 16863 12103 16915
rect 12159 16863 12211 16915
rect 12267 16863 12319 16915
rect 12051 16755 12103 16807
rect 12159 16755 12211 16807
rect 12267 16755 12319 16807
rect 12051 16647 12103 16699
rect 12159 16647 12211 16699
rect 12267 16647 12319 16699
rect 12051 16539 12103 16591
rect 12159 16539 12211 16591
rect 12267 16539 12319 16591
rect 12051 16431 12103 16483
rect 12159 16431 12211 16483
rect 12267 16431 12319 16483
rect 12051 16323 12103 16375
rect 12159 16323 12211 16375
rect 12267 16323 12319 16375
rect 12051 16215 12103 16267
rect 12159 16215 12211 16267
rect 12267 16215 12319 16267
rect 12051 16107 12103 16159
rect 12159 16107 12211 16159
rect 12267 16107 12319 16159
rect 12051 15999 12103 16051
rect 12159 15999 12211 16051
rect 12267 15999 12319 16051
rect 12051 15891 12103 15943
rect 12159 15891 12211 15943
rect 12267 15891 12319 15943
rect 12051 15783 12103 15835
rect 12159 15783 12211 15835
rect 12267 15783 12319 15835
rect 12051 15675 12103 15727
rect 12159 15675 12211 15727
rect 12267 15675 12319 15727
rect 12051 15567 12103 15619
rect 12159 15567 12211 15619
rect 12267 15567 12319 15619
rect 12051 15459 12103 15511
rect 12159 15459 12211 15511
rect 12267 15459 12319 15511
rect 12051 15351 12103 15403
rect 12159 15351 12211 15403
rect 12267 15351 12319 15403
rect 12051 15243 12103 15295
rect 12159 15243 12211 15295
rect 12267 15243 12319 15295
rect 12051 15135 12103 15187
rect 12159 15135 12211 15187
rect 12267 15135 12319 15187
rect 12051 15027 12103 15079
rect 12159 15027 12211 15079
rect 12267 15027 12319 15079
rect 12051 14919 12103 14971
rect 12159 14919 12211 14971
rect 12267 14919 12319 14971
rect 12051 14811 12103 14863
rect 12159 14811 12211 14863
rect 12267 14811 12319 14863
rect 12051 14703 12103 14755
rect 12159 14703 12211 14755
rect 12267 14703 12319 14755
rect 12051 14595 12103 14647
rect 12159 14595 12211 14647
rect 12267 14595 12319 14647
rect 12051 14487 12103 14539
rect 12159 14487 12211 14539
rect 12267 14487 12319 14539
rect 12051 14379 12103 14431
rect 12159 14379 12211 14431
rect 12267 14379 12319 14431
rect 12051 14271 12103 14323
rect 12159 14271 12211 14323
rect 12267 14271 12319 14323
rect 12051 14163 12103 14215
rect 12159 14163 12211 14215
rect 12267 14163 12319 14215
rect 12051 14055 12103 14107
rect 12159 14055 12211 14107
rect 12267 14055 12319 14107
rect 12051 13947 12103 13999
rect 12159 13947 12211 13999
rect 12267 13947 12319 13999
rect 12051 13839 12103 13891
rect 12159 13839 12211 13891
rect 12267 13839 12319 13891
rect 12051 13731 12103 13783
rect 12159 13731 12211 13783
rect 12267 13731 12319 13783
rect 12051 13623 12103 13675
rect 12159 13623 12211 13675
rect 12267 13623 12319 13675
rect 12051 13515 12103 13567
rect 12159 13515 12211 13567
rect 12267 13515 12319 13567
rect 12051 13407 12103 13459
rect 12159 13407 12211 13459
rect 12267 13407 12319 13459
rect 12051 13299 12103 13351
rect 12159 13299 12211 13351
rect 12267 13299 12319 13351
rect 12051 13191 12103 13243
rect 12159 13191 12211 13243
rect 12267 13191 12319 13243
rect 12051 13083 12103 13135
rect 12159 13083 12211 13135
rect 12267 13083 12319 13135
rect 12051 12975 12103 13027
rect 12159 12975 12211 13027
rect 12267 12975 12319 13027
rect 12051 12867 12103 12919
rect 12159 12867 12211 12919
rect 12267 12867 12319 12919
rect 12051 12759 12103 12811
rect 12159 12759 12211 12811
rect 12267 12759 12319 12811
rect 1760 12750 1812 12757
rect 1868 12750 1920 12757
rect 1976 12750 2028 12757
rect 2084 12750 2136 12757
rect 2192 12750 2244 12757
rect 2300 12750 2352 12757
rect 2408 12750 2460 12757
rect 2516 12750 2568 12757
rect 2624 12750 2676 12757
rect 2732 12750 2784 12757
rect 2840 12750 2892 12757
rect 2948 12750 3000 12757
rect 3056 12750 3108 12757
rect 3164 12750 3216 12757
rect 3272 12750 3324 12757
rect 3380 12750 3432 12757
rect 3488 12750 3540 12757
rect 3596 12750 3648 12757
rect 3704 12750 3756 12757
rect 4130 12750 4182 12757
rect 4238 12750 4290 12757
rect 4346 12750 4398 12757
rect 4454 12750 4506 12757
rect 4562 12750 4614 12757
rect 4670 12750 4722 12757
rect 4778 12750 4830 12757
rect 4886 12750 4938 12757
rect 4994 12750 5046 12757
rect 5102 12750 5154 12757
rect 5210 12750 5262 12757
rect 5318 12750 5370 12757
rect 5426 12750 5478 12757
rect 5534 12750 5586 12757
rect 5642 12750 5694 12757
rect 5750 12750 5802 12757
rect 5858 12750 5910 12757
rect 5966 12750 6018 12757
rect 6074 12750 6126 12757
rect 6836 12750 6888 12757
rect 6944 12750 6996 12757
rect 7052 12750 7104 12757
rect 7160 12750 7212 12757
rect 7268 12750 7320 12757
rect 7376 12750 7428 12757
rect 7484 12750 7536 12757
rect 7592 12750 7644 12757
rect 7700 12750 7752 12757
rect 7808 12750 7860 12757
rect 7916 12750 7968 12757
rect 8024 12750 8076 12757
rect 8132 12750 8184 12757
rect 8240 12750 8292 12757
rect 8348 12750 8400 12757
rect 8456 12750 8508 12757
rect 8564 12750 8616 12757
rect 8672 12750 8724 12757
rect 8780 12750 8832 12757
rect 9206 12750 9258 12757
rect 9314 12750 9366 12757
rect 9422 12750 9474 12757
rect 9530 12750 9582 12757
rect 9638 12750 9690 12757
rect 9746 12750 9798 12757
rect 9854 12750 9906 12757
rect 9962 12750 10014 12757
rect 10070 12750 10122 12757
rect 10178 12750 10230 12757
rect 10286 12750 10338 12757
rect 10394 12750 10446 12757
rect 10502 12750 10554 12757
rect 10610 12750 10662 12757
rect 10718 12750 10770 12757
rect 10826 12750 10878 12757
rect 10934 12750 10986 12757
rect 11042 12750 11094 12757
rect 11150 12750 11202 12757
rect 643 12651 695 12703
rect 751 12651 803 12703
rect 859 12651 911 12703
rect 1760 12705 1812 12750
rect 1868 12705 1920 12750
rect 1976 12705 2028 12750
rect 2084 12705 2136 12750
rect 2192 12705 2244 12750
rect 2300 12705 2352 12750
rect 2408 12705 2460 12750
rect 2516 12705 2568 12750
rect 2624 12705 2676 12750
rect 2732 12705 2784 12750
rect 2840 12705 2892 12750
rect 2948 12705 3000 12750
rect 3056 12705 3108 12750
rect 3164 12705 3216 12750
rect 3272 12705 3324 12750
rect 3380 12705 3432 12750
rect 3488 12705 3540 12750
rect 3596 12705 3648 12750
rect 3704 12705 3756 12750
rect 4130 12705 4182 12750
rect 4238 12705 4290 12750
rect 4346 12705 4398 12750
rect 4454 12705 4506 12750
rect 4562 12705 4614 12750
rect 4670 12705 4722 12750
rect 4778 12705 4830 12750
rect 4886 12705 4938 12750
rect 4994 12705 5046 12750
rect 5102 12705 5154 12750
rect 5210 12705 5262 12750
rect 5318 12705 5370 12750
rect 5426 12705 5478 12750
rect 5534 12705 5586 12750
rect 5642 12705 5694 12750
rect 5750 12705 5802 12750
rect 5858 12705 5910 12750
rect 5966 12705 6018 12750
rect 6074 12705 6126 12750
rect 6836 12705 6888 12750
rect 6944 12705 6996 12750
rect 7052 12705 7104 12750
rect 7160 12705 7212 12750
rect 7268 12705 7320 12750
rect 7376 12705 7428 12750
rect 7484 12705 7536 12750
rect 7592 12705 7644 12750
rect 7700 12705 7752 12750
rect 7808 12705 7860 12750
rect 7916 12705 7968 12750
rect 8024 12705 8076 12750
rect 8132 12705 8184 12750
rect 8240 12705 8292 12750
rect 8348 12705 8400 12750
rect 8456 12705 8508 12750
rect 8564 12705 8616 12750
rect 8672 12705 8724 12750
rect 8780 12705 8832 12750
rect 9206 12705 9258 12750
rect 9314 12705 9366 12750
rect 9422 12705 9474 12750
rect 9530 12705 9582 12750
rect 9638 12705 9690 12750
rect 9746 12705 9798 12750
rect 9854 12705 9906 12750
rect 9962 12705 10014 12750
rect 10070 12705 10122 12750
rect 10178 12705 10230 12750
rect 10286 12705 10338 12750
rect 10394 12705 10446 12750
rect 10502 12705 10554 12750
rect 10610 12705 10662 12750
rect 10718 12705 10770 12750
rect 10826 12705 10878 12750
rect 10934 12705 10986 12750
rect 11042 12705 11094 12750
rect 11150 12705 11202 12750
rect 1760 12604 1812 12649
rect 1868 12604 1920 12649
rect 1976 12604 2028 12649
rect 2084 12604 2136 12649
rect 2192 12604 2244 12649
rect 2300 12604 2352 12649
rect 2408 12604 2460 12649
rect 2516 12604 2568 12649
rect 2624 12604 2676 12649
rect 2732 12604 2784 12649
rect 2840 12604 2892 12649
rect 2948 12604 3000 12649
rect 3056 12604 3108 12649
rect 3164 12604 3216 12649
rect 3272 12604 3324 12649
rect 3380 12604 3432 12649
rect 3488 12604 3540 12649
rect 3596 12604 3648 12649
rect 3704 12604 3756 12649
rect 4130 12604 4182 12649
rect 4238 12604 4290 12649
rect 4346 12604 4398 12649
rect 4454 12604 4506 12649
rect 4562 12604 4614 12649
rect 4670 12604 4722 12649
rect 4778 12604 4830 12649
rect 4886 12604 4938 12649
rect 4994 12604 5046 12649
rect 5102 12604 5154 12649
rect 5210 12604 5262 12649
rect 5318 12604 5370 12649
rect 5426 12604 5478 12649
rect 5534 12604 5586 12649
rect 5642 12604 5694 12649
rect 5750 12604 5802 12649
rect 5858 12604 5910 12649
rect 5966 12604 6018 12649
rect 6074 12604 6126 12649
rect 6836 12604 6888 12649
rect 6944 12604 6996 12649
rect 7052 12604 7104 12649
rect 7160 12604 7212 12649
rect 7268 12604 7320 12649
rect 7376 12604 7428 12649
rect 7484 12604 7536 12649
rect 7592 12604 7644 12649
rect 7700 12604 7752 12649
rect 7808 12604 7860 12649
rect 7916 12604 7968 12649
rect 8024 12604 8076 12649
rect 8132 12604 8184 12649
rect 8240 12604 8292 12649
rect 8348 12604 8400 12649
rect 8456 12604 8508 12649
rect 8564 12604 8616 12649
rect 8672 12604 8724 12649
rect 8780 12604 8832 12649
rect 9206 12604 9258 12649
rect 9314 12604 9366 12649
rect 9422 12604 9474 12649
rect 9530 12604 9582 12649
rect 9638 12604 9690 12649
rect 9746 12604 9798 12649
rect 9854 12604 9906 12649
rect 9962 12604 10014 12649
rect 10070 12604 10122 12649
rect 10178 12604 10230 12649
rect 10286 12604 10338 12649
rect 10394 12604 10446 12649
rect 10502 12604 10554 12649
rect 10610 12604 10662 12649
rect 10718 12604 10770 12649
rect 10826 12604 10878 12649
rect 10934 12604 10986 12649
rect 11042 12604 11094 12649
rect 11150 12604 11202 12649
rect 12051 12651 12103 12703
rect 12159 12651 12211 12703
rect 12267 12651 12319 12703
rect 1760 12597 1812 12604
rect 1868 12597 1920 12604
rect 1976 12597 2028 12604
rect 2084 12597 2136 12604
rect 2192 12597 2244 12604
rect 2300 12597 2352 12604
rect 2408 12597 2460 12604
rect 2516 12597 2568 12604
rect 2624 12597 2676 12604
rect 2732 12597 2784 12604
rect 2840 12597 2892 12604
rect 2948 12597 3000 12604
rect 3056 12597 3108 12604
rect 3164 12597 3216 12604
rect 3272 12597 3324 12604
rect 3380 12597 3432 12604
rect 3488 12597 3540 12604
rect 3596 12597 3648 12604
rect 3704 12597 3756 12604
rect 4130 12597 4182 12604
rect 4238 12597 4290 12604
rect 4346 12597 4398 12604
rect 4454 12597 4506 12604
rect 4562 12597 4614 12604
rect 4670 12597 4722 12604
rect 4778 12597 4830 12604
rect 4886 12597 4938 12604
rect 4994 12597 5046 12604
rect 5102 12597 5154 12604
rect 5210 12597 5262 12604
rect 5318 12597 5370 12604
rect 5426 12597 5478 12604
rect 5534 12597 5586 12604
rect 5642 12597 5694 12604
rect 5750 12597 5802 12604
rect 5858 12597 5910 12604
rect 5966 12597 6018 12604
rect 6074 12597 6126 12604
rect 6836 12597 6888 12604
rect 6944 12597 6996 12604
rect 7052 12597 7104 12604
rect 7160 12597 7212 12604
rect 7268 12597 7320 12604
rect 7376 12597 7428 12604
rect 7484 12597 7536 12604
rect 7592 12597 7644 12604
rect 7700 12597 7752 12604
rect 7808 12597 7860 12604
rect 7916 12597 7968 12604
rect 8024 12597 8076 12604
rect 8132 12597 8184 12604
rect 8240 12597 8292 12604
rect 8348 12597 8400 12604
rect 8456 12597 8508 12604
rect 8564 12597 8616 12604
rect 8672 12597 8724 12604
rect 8780 12597 8832 12604
rect 9206 12597 9258 12604
rect 9314 12597 9366 12604
rect 9422 12597 9474 12604
rect 9530 12597 9582 12604
rect 9638 12597 9690 12604
rect 9746 12597 9798 12604
rect 9854 12597 9906 12604
rect 9962 12597 10014 12604
rect 10070 12597 10122 12604
rect 10178 12597 10230 12604
rect 10286 12597 10338 12604
rect 10394 12597 10446 12604
rect 10502 12597 10554 12604
rect 10610 12597 10662 12604
rect 10718 12597 10770 12604
rect 10826 12597 10878 12604
rect 10934 12597 10986 12604
rect 11042 12597 11094 12604
rect 11150 12597 11202 12604
rect 643 12543 695 12595
rect 751 12543 803 12595
rect 859 12543 911 12595
rect 643 12435 695 12487
rect 751 12435 803 12487
rect 859 12435 911 12487
rect 643 12327 695 12379
rect 751 12327 803 12379
rect 859 12327 911 12379
rect 643 12219 695 12271
rect 751 12219 803 12271
rect 859 12219 911 12271
rect 643 12111 695 12163
rect 751 12111 803 12163
rect 859 12111 911 12163
rect 643 12003 695 12055
rect 751 12003 803 12055
rect 859 12003 911 12055
rect 643 11895 695 11947
rect 751 11895 803 11947
rect 859 11895 911 11947
rect 643 11787 695 11839
rect 751 11787 803 11839
rect 859 11787 911 11839
rect 643 11679 695 11731
rect 751 11679 803 11731
rect 859 11679 911 11731
rect 643 11571 695 11623
rect 751 11571 803 11623
rect 859 11571 911 11623
rect 643 11463 695 11515
rect 751 11463 803 11515
rect 859 11463 911 11515
rect 643 11355 695 11407
rect 751 11355 803 11407
rect 859 11355 911 11407
rect 643 11247 695 11299
rect 751 11247 803 11299
rect 859 11247 911 11299
rect 643 11139 695 11191
rect 751 11139 803 11191
rect 859 11139 911 11191
rect 643 11031 695 11083
rect 751 11031 803 11083
rect 859 11031 911 11083
rect 643 10923 695 10975
rect 751 10923 803 10975
rect 859 10923 911 10975
rect 643 10815 695 10867
rect 751 10815 803 10867
rect 859 10815 911 10867
rect 643 10707 695 10759
rect 751 10707 803 10759
rect 859 10707 911 10759
rect 643 10599 695 10651
rect 751 10599 803 10651
rect 859 10599 911 10651
rect 643 10491 695 10543
rect 751 10491 803 10543
rect 859 10491 911 10543
rect 643 10383 695 10435
rect 751 10383 803 10435
rect 859 10383 911 10435
rect 643 10275 695 10327
rect 751 10275 803 10327
rect 859 10275 911 10327
rect 643 10167 695 10219
rect 751 10167 803 10219
rect 859 10167 911 10219
rect 643 10059 695 10111
rect 751 10059 803 10111
rect 859 10059 911 10111
rect 643 9951 695 10003
rect 751 9951 803 10003
rect 859 9951 911 10003
rect 643 9843 695 9895
rect 751 9843 803 9895
rect 859 9843 911 9895
rect 643 9735 695 9787
rect 751 9735 803 9787
rect 859 9735 911 9787
rect 643 9627 695 9679
rect 751 9627 803 9679
rect 859 9627 911 9679
rect 643 9519 695 9571
rect 751 9519 803 9571
rect 859 9519 911 9571
rect 643 9411 695 9463
rect 751 9411 803 9463
rect 859 9411 911 9463
rect 643 9303 695 9355
rect 751 9303 803 9355
rect 859 9303 911 9355
rect 643 9195 695 9247
rect 751 9195 803 9247
rect 859 9195 911 9247
rect 643 9087 695 9139
rect 751 9087 803 9139
rect 859 9087 911 9139
rect 643 8979 695 9031
rect 751 8979 803 9031
rect 859 8979 911 9031
rect 643 8871 695 8923
rect 751 8871 803 8923
rect 859 8871 911 8923
rect 643 8763 695 8815
rect 751 8763 803 8815
rect 859 8763 911 8815
rect 643 8655 695 8707
rect 751 8655 803 8707
rect 859 8655 911 8707
rect 643 8547 695 8599
rect 751 8547 803 8599
rect 859 8547 911 8599
rect 643 8439 695 8491
rect 751 8439 803 8491
rect 859 8439 911 8491
rect 643 8331 695 8383
rect 751 8331 803 8383
rect 859 8331 911 8383
rect 643 8223 695 8275
rect 751 8223 803 8275
rect 859 8223 911 8275
rect 643 8115 695 8167
rect 751 8115 803 8167
rect 859 8115 911 8167
rect 643 8007 695 8059
rect 751 8007 803 8059
rect 859 8007 911 8059
rect 643 7899 695 7951
rect 751 7899 803 7951
rect 859 7899 911 7951
rect 643 7791 695 7843
rect 751 7791 803 7843
rect 859 7791 911 7843
rect 643 7683 695 7735
rect 751 7683 803 7735
rect 859 7683 911 7735
rect 643 7575 695 7627
rect 751 7575 803 7627
rect 859 7575 911 7627
rect 643 7467 695 7519
rect 751 7467 803 7519
rect 859 7467 911 7519
rect 643 7359 695 7411
rect 751 7359 803 7411
rect 859 7359 911 7411
rect 643 7251 695 7303
rect 751 7251 803 7303
rect 859 7251 911 7303
rect 643 7143 695 7195
rect 751 7143 803 7195
rect 859 7143 911 7195
rect 643 7035 695 7087
rect 751 7035 803 7087
rect 859 7035 911 7087
rect 643 6927 695 6979
rect 751 6927 803 6979
rect 859 6927 911 6979
rect 1760 12204 1812 12207
rect 1868 12204 1920 12207
rect 1976 12204 2028 12207
rect 2084 12204 2136 12207
rect 2192 12204 2244 12207
rect 2300 12204 2352 12207
rect 2408 12204 2460 12207
rect 2516 12204 2568 12207
rect 2624 12204 2676 12207
rect 2732 12204 2784 12207
rect 2840 12204 2892 12207
rect 2948 12204 3000 12207
rect 3056 12204 3108 12207
rect 3164 12204 3216 12207
rect 3272 12204 3324 12207
rect 3380 12204 3432 12207
rect 3488 12204 3540 12207
rect 3596 12204 3648 12207
rect 3704 12204 3756 12207
rect 4130 12204 4182 12207
rect 4238 12204 4290 12207
rect 4346 12204 4398 12207
rect 4454 12204 4506 12207
rect 4562 12204 4614 12207
rect 4670 12204 4722 12207
rect 4778 12204 4830 12207
rect 4886 12204 4938 12207
rect 4994 12204 5046 12207
rect 5102 12204 5154 12207
rect 5210 12204 5262 12207
rect 5318 12204 5370 12207
rect 5426 12204 5478 12207
rect 5534 12204 5586 12207
rect 5642 12204 5694 12207
rect 5750 12204 5802 12207
rect 5858 12204 5910 12207
rect 5966 12204 6018 12207
rect 6074 12204 6126 12207
rect 6836 12204 6888 12207
rect 6944 12204 6996 12207
rect 7052 12204 7104 12207
rect 7160 12204 7212 12207
rect 7268 12204 7320 12207
rect 7376 12204 7428 12207
rect 7484 12204 7536 12207
rect 7592 12204 7644 12207
rect 7700 12204 7752 12207
rect 7808 12204 7860 12207
rect 7916 12204 7968 12207
rect 8024 12204 8076 12207
rect 8132 12204 8184 12207
rect 8240 12204 8292 12207
rect 8348 12204 8400 12207
rect 8456 12204 8508 12207
rect 8564 12204 8616 12207
rect 8672 12204 8724 12207
rect 8780 12204 8832 12207
rect 9206 12204 9258 12207
rect 9314 12204 9366 12207
rect 9422 12204 9474 12207
rect 9530 12204 9582 12207
rect 9638 12204 9690 12207
rect 9746 12204 9798 12207
rect 9854 12204 9906 12207
rect 9962 12204 10014 12207
rect 10070 12204 10122 12207
rect 10178 12204 10230 12207
rect 10286 12204 10338 12207
rect 10394 12204 10446 12207
rect 10502 12204 10554 12207
rect 10610 12204 10662 12207
rect 10718 12204 10770 12207
rect 10826 12204 10878 12207
rect 10934 12204 10986 12207
rect 11042 12204 11094 12207
rect 11150 12204 11202 12207
rect 1760 12158 1812 12204
rect 1868 12158 1920 12204
rect 1976 12158 2028 12204
rect 2084 12158 2136 12204
rect 2192 12158 2244 12204
rect 2300 12158 2352 12204
rect 2408 12158 2460 12204
rect 2516 12158 2568 12204
rect 2624 12158 2676 12204
rect 2732 12158 2784 12204
rect 2840 12158 2892 12204
rect 2948 12158 3000 12204
rect 3056 12158 3108 12204
rect 3164 12158 3216 12204
rect 3272 12158 3324 12204
rect 3380 12158 3432 12204
rect 3488 12158 3540 12204
rect 3596 12158 3648 12204
rect 3704 12158 3756 12204
rect 4130 12158 4182 12204
rect 4238 12158 4290 12204
rect 4346 12158 4398 12204
rect 4454 12158 4506 12204
rect 4562 12158 4614 12204
rect 4670 12158 4722 12204
rect 4778 12158 4830 12204
rect 4886 12158 4938 12204
rect 4994 12158 5046 12204
rect 5102 12158 5154 12204
rect 5210 12158 5262 12204
rect 5318 12158 5370 12204
rect 5426 12158 5478 12204
rect 5534 12158 5586 12204
rect 5642 12158 5694 12204
rect 5750 12158 5802 12204
rect 5858 12158 5910 12204
rect 5966 12158 6018 12204
rect 6074 12158 6126 12204
rect 6836 12158 6888 12204
rect 6944 12158 6996 12204
rect 7052 12158 7104 12204
rect 7160 12158 7212 12204
rect 7268 12158 7320 12204
rect 7376 12158 7428 12204
rect 7484 12158 7536 12204
rect 7592 12158 7644 12204
rect 7700 12158 7752 12204
rect 7808 12158 7860 12204
rect 7916 12158 7968 12204
rect 8024 12158 8076 12204
rect 8132 12158 8184 12204
rect 8240 12158 8292 12204
rect 8348 12158 8400 12204
rect 8456 12158 8508 12204
rect 8564 12158 8616 12204
rect 8672 12158 8724 12204
rect 8780 12158 8832 12204
rect 9206 12158 9258 12204
rect 9314 12158 9366 12204
rect 9422 12158 9474 12204
rect 9530 12158 9582 12204
rect 9638 12158 9690 12204
rect 9746 12158 9798 12204
rect 9854 12158 9906 12204
rect 9962 12158 10014 12204
rect 10070 12158 10122 12204
rect 10178 12158 10230 12204
rect 10286 12158 10338 12204
rect 10394 12158 10446 12204
rect 10502 12158 10554 12204
rect 10610 12158 10662 12204
rect 10718 12158 10770 12204
rect 10826 12158 10878 12204
rect 10934 12158 10986 12204
rect 11042 12158 11094 12204
rect 11150 12158 11202 12204
rect 1760 12155 1812 12158
rect 1868 12155 1920 12158
rect 1976 12155 2028 12158
rect 2084 12155 2136 12158
rect 2192 12155 2244 12158
rect 2300 12155 2352 12158
rect 2408 12155 2460 12158
rect 2516 12155 2568 12158
rect 2624 12155 2676 12158
rect 2732 12155 2784 12158
rect 2840 12155 2892 12158
rect 2948 12155 3000 12158
rect 3056 12155 3108 12158
rect 3164 12155 3216 12158
rect 3272 12155 3324 12158
rect 3380 12155 3432 12158
rect 3488 12155 3540 12158
rect 3596 12155 3648 12158
rect 3704 12155 3756 12158
rect 4130 12155 4182 12158
rect 4238 12155 4290 12158
rect 4346 12155 4398 12158
rect 4454 12155 4506 12158
rect 4562 12155 4614 12158
rect 4670 12155 4722 12158
rect 4778 12155 4830 12158
rect 4886 12155 4938 12158
rect 4994 12155 5046 12158
rect 5102 12155 5154 12158
rect 5210 12155 5262 12158
rect 5318 12155 5370 12158
rect 5426 12155 5478 12158
rect 5534 12155 5586 12158
rect 5642 12155 5694 12158
rect 5750 12155 5802 12158
rect 5858 12155 5910 12158
rect 5966 12155 6018 12158
rect 6074 12155 6126 12158
rect 6836 12155 6888 12158
rect 6944 12155 6996 12158
rect 7052 12155 7104 12158
rect 7160 12155 7212 12158
rect 7268 12155 7320 12158
rect 7376 12155 7428 12158
rect 7484 12155 7536 12158
rect 7592 12155 7644 12158
rect 7700 12155 7752 12158
rect 7808 12155 7860 12158
rect 7916 12155 7968 12158
rect 8024 12155 8076 12158
rect 8132 12155 8184 12158
rect 8240 12155 8292 12158
rect 8348 12155 8400 12158
rect 8456 12155 8508 12158
rect 8564 12155 8616 12158
rect 8672 12155 8724 12158
rect 8780 12155 8832 12158
rect 9206 12155 9258 12158
rect 9314 12155 9366 12158
rect 9422 12155 9474 12158
rect 9530 12155 9582 12158
rect 9638 12155 9690 12158
rect 9746 12155 9798 12158
rect 9854 12155 9906 12158
rect 9962 12155 10014 12158
rect 10070 12155 10122 12158
rect 10178 12155 10230 12158
rect 10286 12155 10338 12158
rect 10394 12155 10446 12158
rect 10502 12155 10554 12158
rect 10610 12155 10662 12158
rect 10718 12155 10770 12158
rect 10826 12155 10878 12158
rect 10934 12155 10986 12158
rect 11042 12155 11094 12158
rect 11150 12155 11202 12158
rect 1233 12091 1285 12143
rect 1341 12091 1393 12143
rect 1233 11983 1256 12035
rect 1256 11983 1285 12035
rect 1341 11983 1393 12035
rect 1233 11875 1256 11927
rect 1256 11875 1285 11927
rect 1341 11875 1393 11927
rect 1233 11767 1256 11819
rect 1256 11767 1285 11819
rect 1341 11767 1393 11819
rect 1233 11659 1256 11711
rect 1256 11659 1285 11711
rect 1341 11659 1393 11711
rect 1233 11551 1256 11603
rect 1256 11551 1285 11603
rect 1341 11551 1393 11603
rect 1233 11443 1256 11495
rect 1256 11443 1285 11495
rect 1341 11443 1393 11495
rect 1233 11335 1256 11387
rect 1256 11335 1285 11387
rect 1341 11335 1393 11387
rect 1233 11227 1256 11279
rect 1256 11227 1285 11279
rect 1341 11227 1393 11279
rect 1233 11119 1256 11171
rect 1256 11119 1285 11171
rect 1341 11119 1393 11171
rect 1233 11011 1256 11063
rect 1256 11011 1285 11063
rect 1341 11011 1393 11063
rect 1233 10903 1256 10955
rect 1256 10903 1285 10955
rect 1341 10903 1393 10955
rect 1233 10795 1256 10847
rect 1256 10795 1285 10847
rect 1341 10795 1393 10847
rect 1233 10687 1256 10739
rect 1256 10687 1285 10739
rect 1341 10687 1393 10739
rect 1233 10579 1256 10631
rect 1256 10579 1285 10631
rect 1341 10579 1393 10631
rect 1233 10471 1256 10523
rect 1256 10471 1285 10523
rect 1341 10471 1393 10523
rect 1233 10363 1256 10415
rect 1256 10363 1285 10415
rect 1341 10363 1393 10415
rect 1233 10255 1256 10307
rect 1256 10255 1285 10307
rect 1341 10255 1393 10307
rect 1233 10147 1256 10199
rect 1256 10147 1285 10199
rect 1341 10147 1393 10199
rect 1233 10039 1256 10091
rect 1256 10039 1285 10091
rect 1341 10039 1393 10091
rect 1233 9931 1256 9983
rect 1256 9931 1285 9983
rect 1341 9931 1393 9983
rect 1233 9823 1256 9875
rect 1256 9823 1285 9875
rect 1341 9823 1393 9875
rect 1233 9715 1256 9767
rect 1256 9715 1285 9767
rect 1341 9715 1393 9767
rect 1233 9607 1256 9659
rect 1256 9607 1285 9659
rect 1341 9607 1393 9659
rect 1233 9499 1256 9551
rect 1256 9499 1285 9551
rect 1341 9499 1393 9551
rect 1233 9391 1256 9443
rect 1256 9391 1285 9443
rect 1341 9391 1393 9443
rect 1233 9283 1256 9335
rect 1256 9283 1285 9335
rect 1341 9283 1393 9335
rect 1233 9175 1256 9227
rect 1256 9175 1285 9227
rect 1341 9175 1393 9227
rect 1233 9067 1256 9119
rect 1256 9067 1285 9119
rect 1341 9067 1393 9119
rect 1233 8959 1256 9011
rect 1256 8959 1285 9011
rect 1341 8959 1393 9011
rect 1233 8851 1256 8903
rect 1256 8851 1285 8903
rect 1341 8851 1393 8903
rect 1233 8743 1256 8795
rect 1256 8743 1285 8795
rect 1341 8743 1393 8795
rect 1233 8635 1256 8687
rect 1256 8635 1285 8687
rect 1341 8635 1393 8687
rect 1233 8527 1256 8579
rect 1256 8527 1285 8579
rect 1341 8527 1393 8579
rect 1233 8419 1256 8471
rect 1256 8419 1285 8471
rect 1341 8419 1393 8471
rect 1233 8311 1256 8363
rect 1256 8311 1285 8363
rect 1341 8311 1393 8363
rect 1233 8203 1256 8255
rect 1256 8203 1285 8255
rect 1341 8203 1393 8255
rect 1233 8095 1256 8147
rect 1256 8095 1285 8147
rect 1341 8095 1393 8147
rect 1233 7987 1256 8039
rect 1256 7987 1285 8039
rect 1341 7987 1393 8039
rect 1233 7879 1256 7931
rect 1256 7879 1285 7931
rect 1341 7879 1393 7931
rect 1233 7771 1256 7823
rect 1256 7771 1285 7823
rect 1341 7771 1393 7823
rect 1233 7663 1256 7715
rect 1256 7663 1285 7715
rect 1341 7663 1393 7715
rect 1233 7555 1256 7607
rect 1256 7555 1285 7607
rect 1341 7555 1393 7607
rect 1233 7447 1256 7499
rect 1256 7447 1285 7499
rect 1341 7447 1393 7499
rect 11569 12091 11621 12143
rect 11677 12091 11729 12143
rect 1493 11960 1545 11963
rect 1601 11960 1653 11963
rect 3863 11960 3915 11963
rect 3971 11960 4023 11963
rect 6239 11960 6291 11963
rect 6347 11960 6399 11963
rect 6455 11960 6507 11963
rect 6563 11960 6615 11963
rect 6671 11960 6723 11963
rect 8939 11960 8991 11963
rect 9047 11960 9099 11963
rect 11309 11960 11361 11963
rect 11417 11960 11469 11963
rect 1493 11914 1494 11960
rect 1494 11914 1545 11960
rect 1601 11914 1653 11960
rect 3863 11914 3915 11960
rect 3971 11914 4023 11960
rect 6239 11914 6291 11960
rect 6347 11914 6399 11960
rect 6455 11914 6507 11960
rect 6563 11914 6615 11960
rect 6671 11914 6723 11960
rect 8939 11914 8991 11960
rect 9047 11914 9099 11960
rect 11309 11914 11361 11960
rect 11417 11914 11468 11960
rect 11468 11914 11469 11960
rect 1493 11911 1545 11914
rect 1601 11911 1653 11914
rect 3863 11911 3915 11914
rect 3971 11911 4023 11914
rect 6239 11911 6291 11914
rect 6347 11911 6399 11914
rect 6455 11911 6507 11914
rect 6563 11911 6615 11914
rect 6671 11911 6723 11914
rect 8939 11911 8991 11914
rect 9047 11911 9099 11914
rect 11309 11911 11361 11914
rect 11417 11911 11469 11914
rect 1760 11716 1812 11719
rect 1868 11716 1920 11719
rect 1976 11716 2028 11719
rect 2084 11716 2136 11719
rect 2192 11716 2244 11719
rect 2300 11716 2352 11719
rect 2408 11716 2460 11719
rect 2516 11716 2568 11719
rect 2624 11716 2676 11719
rect 2732 11716 2784 11719
rect 2840 11716 2892 11719
rect 2948 11716 3000 11719
rect 3056 11716 3108 11719
rect 3164 11716 3216 11719
rect 3272 11716 3324 11719
rect 3380 11716 3432 11719
rect 3488 11716 3540 11719
rect 3596 11716 3648 11719
rect 3704 11716 3756 11719
rect 4130 11716 4182 11719
rect 4238 11716 4290 11719
rect 4346 11716 4398 11719
rect 4454 11716 4506 11719
rect 4562 11716 4614 11719
rect 4670 11716 4722 11719
rect 4778 11716 4830 11719
rect 4886 11716 4938 11719
rect 4994 11716 5046 11719
rect 5102 11716 5154 11719
rect 5210 11716 5262 11719
rect 5318 11716 5370 11719
rect 5426 11716 5478 11719
rect 5534 11716 5586 11719
rect 5642 11716 5694 11719
rect 5750 11716 5802 11719
rect 5858 11716 5910 11719
rect 5966 11716 6018 11719
rect 6074 11716 6126 11719
rect 6836 11716 6888 11719
rect 6944 11716 6996 11719
rect 7052 11716 7104 11719
rect 7160 11716 7212 11719
rect 7268 11716 7320 11719
rect 7376 11716 7428 11719
rect 7484 11716 7536 11719
rect 7592 11716 7644 11719
rect 7700 11716 7752 11719
rect 7808 11716 7860 11719
rect 7916 11716 7968 11719
rect 8024 11716 8076 11719
rect 8132 11716 8184 11719
rect 8240 11716 8292 11719
rect 8348 11716 8400 11719
rect 8456 11716 8508 11719
rect 8564 11716 8616 11719
rect 8672 11716 8724 11719
rect 8780 11716 8832 11719
rect 9206 11716 9258 11719
rect 9314 11716 9366 11719
rect 9422 11716 9474 11719
rect 9530 11716 9582 11719
rect 9638 11716 9690 11719
rect 9746 11716 9798 11719
rect 9854 11716 9906 11719
rect 9962 11716 10014 11719
rect 10070 11716 10122 11719
rect 10178 11716 10230 11719
rect 10286 11716 10338 11719
rect 10394 11716 10446 11719
rect 10502 11716 10554 11719
rect 10610 11716 10662 11719
rect 10718 11716 10770 11719
rect 10826 11716 10878 11719
rect 10934 11716 10986 11719
rect 11042 11716 11094 11719
rect 11150 11716 11202 11719
rect 1760 11670 1812 11716
rect 1868 11670 1920 11716
rect 1976 11670 2028 11716
rect 2084 11670 2136 11716
rect 2192 11670 2244 11716
rect 2300 11670 2352 11716
rect 2408 11670 2460 11716
rect 2516 11670 2568 11716
rect 2624 11670 2676 11716
rect 2732 11670 2784 11716
rect 2840 11670 2892 11716
rect 2948 11670 3000 11716
rect 3056 11670 3108 11716
rect 3164 11670 3216 11716
rect 3272 11670 3324 11716
rect 3380 11670 3432 11716
rect 3488 11670 3540 11716
rect 3596 11670 3648 11716
rect 3704 11670 3756 11716
rect 4130 11670 4182 11716
rect 4238 11670 4290 11716
rect 4346 11670 4398 11716
rect 4454 11670 4506 11716
rect 4562 11670 4614 11716
rect 4670 11670 4722 11716
rect 4778 11670 4830 11716
rect 4886 11670 4938 11716
rect 4994 11670 5046 11716
rect 5102 11670 5154 11716
rect 5210 11670 5262 11716
rect 5318 11670 5370 11716
rect 5426 11670 5478 11716
rect 5534 11670 5586 11716
rect 5642 11670 5694 11716
rect 5750 11670 5802 11716
rect 5858 11670 5910 11716
rect 5966 11670 6018 11716
rect 6074 11670 6126 11716
rect 6836 11670 6888 11716
rect 6944 11670 6996 11716
rect 7052 11670 7104 11716
rect 7160 11670 7212 11716
rect 7268 11670 7320 11716
rect 7376 11670 7428 11716
rect 7484 11670 7536 11716
rect 7592 11670 7644 11716
rect 7700 11670 7752 11716
rect 7808 11670 7860 11716
rect 7916 11670 7968 11716
rect 8024 11670 8076 11716
rect 8132 11670 8184 11716
rect 8240 11670 8292 11716
rect 8348 11670 8400 11716
rect 8456 11670 8508 11716
rect 8564 11670 8616 11716
rect 8672 11670 8724 11716
rect 8780 11670 8832 11716
rect 9206 11670 9258 11716
rect 9314 11670 9366 11716
rect 9422 11670 9474 11716
rect 9530 11670 9582 11716
rect 9638 11670 9690 11716
rect 9746 11670 9798 11716
rect 9854 11670 9906 11716
rect 9962 11670 10014 11716
rect 10070 11670 10122 11716
rect 10178 11670 10230 11716
rect 10286 11670 10338 11716
rect 10394 11670 10446 11716
rect 10502 11670 10554 11716
rect 10610 11670 10662 11716
rect 10718 11670 10770 11716
rect 10826 11670 10878 11716
rect 10934 11670 10986 11716
rect 11042 11670 11094 11716
rect 11150 11670 11202 11716
rect 1760 11667 1812 11670
rect 1868 11667 1920 11670
rect 1976 11667 2028 11670
rect 2084 11667 2136 11670
rect 2192 11667 2244 11670
rect 2300 11667 2352 11670
rect 2408 11667 2460 11670
rect 2516 11667 2568 11670
rect 2624 11667 2676 11670
rect 2732 11667 2784 11670
rect 2840 11667 2892 11670
rect 2948 11667 3000 11670
rect 3056 11667 3108 11670
rect 3164 11667 3216 11670
rect 3272 11667 3324 11670
rect 3380 11667 3432 11670
rect 3488 11667 3540 11670
rect 3596 11667 3648 11670
rect 3704 11667 3756 11670
rect 4130 11667 4182 11670
rect 4238 11667 4290 11670
rect 4346 11667 4398 11670
rect 4454 11667 4506 11670
rect 4562 11667 4614 11670
rect 4670 11667 4722 11670
rect 4778 11667 4830 11670
rect 4886 11667 4938 11670
rect 4994 11667 5046 11670
rect 5102 11667 5154 11670
rect 5210 11667 5262 11670
rect 5318 11667 5370 11670
rect 5426 11667 5478 11670
rect 5534 11667 5586 11670
rect 5642 11667 5694 11670
rect 5750 11667 5802 11670
rect 5858 11667 5910 11670
rect 5966 11667 6018 11670
rect 6074 11667 6126 11670
rect 6836 11667 6888 11670
rect 6944 11667 6996 11670
rect 7052 11667 7104 11670
rect 7160 11667 7212 11670
rect 7268 11667 7320 11670
rect 7376 11667 7428 11670
rect 7484 11667 7536 11670
rect 7592 11667 7644 11670
rect 7700 11667 7752 11670
rect 7808 11667 7860 11670
rect 7916 11667 7968 11670
rect 8024 11667 8076 11670
rect 8132 11667 8184 11670
rect 8240 11667 8292 11670
rect 8348 11667 8400 11670
rect 8456 11667 8508 11670
rect 8564 11667 8616 11670
rect 8672 11667 8724 11670
rect 8780 11667 8832 11670
rect 9206 11667 9258 11670
rect 9314 11667 9366 11670
rect 9422 11667 9474 11670
rect 9530 11667 9582 11670
rect 9638 11667 9690 11670
rect 9746 11667 9798 11670
rect 9854 11667 9906 11670
rect 9962 11667 10014 11670
rect 10070 11667 10122 11670
rect 10178 11667 10230 11670
rect 10286 11667 10338 11670
rect 10394 11667 10446 11670
rect 10502 11667 10554 11670
rect 10610 11667 10662 11670
rect 10718 11667 10770 11670
rect 10826 11667 10878 11670
rect 10934 11667 10986 11670
rect 11042 11667 11094 11670
rect 11150 11667 11202 11670
rect 1493 11472 1545 11475
rect 1601 11472 1653 11475
rect 3863 11472 3915 11475
rect 3971 11472 4023 11475
rect 6239 11472 6291 11475
rect 6347 11472 6399 11475
rect 6455 11472 6507 11475
rect 6563 11472 6615 11475
rect 6671 11472 6723 11475
rect 8939 11472 8991 11475
rect 9047 11472 9099 11475
rect 11309 11472 11361 11475
rect 11417 11472 11469 11475
rect 1493 11426 1494 11472
rect 1494 11426 1545 11472
rect 1601 11426 1653 11472
rect 3863 11426 3915 11472
rect 3971 11426 4023 11472
rect 6239 11426 6291 11472
rect 6347 11426 6399 11472
rect 6455 11426 6507 11472
rect 6563 11426 6615 11472
rect 6671 11426 6723 11472
rect 8939 11426 8991 11472
rect 9047 11426 9099 11472
rect 11309 11426 11361 11472
rect 11417 11426 11468 11472
rect 11468 11426 11469 11472
rect 1493 11423 1545 11426
rect 1601 11423 1653 11426
rect 3863 11423 3915 11426
rect 3971 11423 4023 11426
rect 6239 11423 6291 11426
rect 6347 11423 6399 11426
rect 6455 11423 6507 11426
rect 6563 11423 6615 11426
rect 6671 11423 6723 11426
rect 8939 11423 8991 11426
rect 9047 11423 9099 11426
rect 11309 11423 11361 11426
rect 11417 11423 11469 11426
rect 1760 11228 1812 11231
rect 1868 11228 1920 11231
rect 1976 11228 2028 11231
rect 2084 11228 2136 11231
rect 2192 11228 2244 11231
rect 2300 11228 2352 11231
rect 2408 11228 2460 11231
rect 2516 11228 2568 11231
rect 2624 11228 2676 11231
rect 2732 11228 2784 11231
rect 2840 11228 2892 11231
rect 2948 11228 3000 11231
rect 3056 11228 3108 11231
rect 3164 11228 3216 11231
rect 3272 11228 3324 11231
rect 3380 11228 3432 11231
rect 3488 11228 3540 11231
rect 3596 11228 3648 11231
rect 3704 11228 3756 11231
rect 4130 11228 4182 11231
rect 4238 11228 4290 11231
rect 4346 11228 4398 11231
rect 4454 11228 4506 11231
rect 4562 11228 4614 11231
rect 4670 11228 4722 11231
rect 4778 11228 4830 11231
rect 4886 11228 4938 11231
rect 4994 11228 5046 11231
rect 5102 11228 5154 11231
rect 5210 11228 5262 11231
rect 5318 11228 5370 11231
rect 5426 11228 5478 11231
rect 5534 11228 5586 11231
rect 5642 11228 5694 11231
rect 5750 11228 5802 11231
rect 5858 11228 5910 11231
rect 5966 11228 6018 11231
rect 6074 11228 6126 11231
rect 6836 11228 6888 11231
rect 6944 11228 6996 11231
rect 7052 11228 7104 11231
rect 7160 11228 7212 11231
rect 7268 11228 7320 11231
rect 7376 11228 7428 11231
rect 7484 11228 7536 11231
rect 7592 11228 7644 11231
rect 7700 11228 7752 11231
rect 7808 11228 7860 11231
rect 7916 11228 7968 11231
rect 8024 11228 8076 11231
rect 8132 11228 8184 11231
rect 8240 11228 8292 11231
rect 8348 11228 8400 11231
rect 8456 11228 8508 11231
rect 8564 11228 8616 11231
rect 8672 11228 8724 11231
rect 8780 11228 8832 11231
rect 9206 11228 9258 11231
rect 9314 11228 9366 11231
rect 9422 11228 9474 11231
rect 9530 11228 9582 11231
rect 9638 11228 9690 11231
rect 9746 11228 9798 11231
rect 9854 11228 9906 11231
rect 9962 11228 10014 11231
rect 10070 11228 10122 11231
rect 10178 11228 10230 11231
rect 10286 11228 10338 11231
rect 10394 11228 10446 11231
rect 10502 11228 10554 11231
rect 10610 11228 10662 11231
rect 10718 11228 10770 11231
rect 10826 11228 10878 11231
rect 10934 11228 10986 11231
rect 11042 11228 11094 11231
rect 11150 11228 11202 11231
rect 1760 11182 1812 11228
rect 1868 11182 1920 11228
rect 1976 11182 2028 11228
rect 2084 11182 2136 11228
rect 2192 11182 2244 11228
rect 2300 11182 2352 11228
rect 2408 11182 2460 11228
rect 2516 11182 2568 11228
rect 2624 11182 2676 11228
rect 2732 11182 2784 11228
rect 2840 11182 2892 11228
rect 2948 11182 3000 11228
rect 3056 11182 3108 11228
rect 3164 11182 3216 11228
rect 3272 11182 3324 11228
rect 3380 11182 3432 11228
rect 3488 11182 3540 11228
rect 3596 11182 3648 11228
rect 3704 11182 3756 11228
rect 4130 11182 4182 11228
rect 4238 11182 4290 11228
rect 4346 11182 4398 11228
rect 4454 11182 4506 11228
rect 4562 11182 4614 11228
rect 4670 11182 4722 11228
rect 4778 11182 4830 11228
rect 4886 11182 4938 11228
rect 4994 11182 5046 11228
rect 5102 11182 5154 11228
rect 5210 11182 5262 11228
rect 5318 11182 5370 11228
rect 5426 11182 5478 11228
rect 5534 11182 5586 11228
rect 5642 11182 5694 11228
rect 5750 11182 5802 11228
rect 5858 11182 5910 11228
rect 5966 11182 6018 11228
rect 6074 11182 6126 11228
rect 6836 11182 6888 11228
rect 6944 11182 6996 11228
rect 7052 11182 7104 11228
rect 7160 11182 7212 11228
rect 7268 11182 7320 11228
rect 7376 11182 7428 11228
rect 7484 11182 7536 11228
rect 7592 11182 7644 11228
rect 7700 11182 7752 11228
rect 7808 11182 7860 11228
rect 7916 11182 7968 11228
rect 8024 11182 8076 11228
rect 8132 11182 8184 11228
rect 8240 11182 8292 11228
rect 8348 11182 8400 11228
rect 8456 11182 8508 11228
rect 8564 11182 8616 11228
rect 8672 11182 8724 11228
rect 8780 11182 8832 11228
rect 9206 11182 9258 11228
rect 9314 11182 9366 11228
rect 9422 11182 9474 11228
rect 9530 11182 9582 11228
rect 9638 11182 9690 11228
rect 9746 11182 9798 11228
rect 9854 11182 9906 11228
rect 9962 11182 10014 11228
rect 10070 11182 10122 11228
rect 10178 11182 10230 11228
rect 10286 11182 10338 11228
rect 10394 11182 10446 11228
rect 10502 11182 10554 11228
rect 10610 11182 10662 11228
rect 10718 11182 10770 11228
rect 10826 11182 10878 11228
rect 10934 11182 10986 11228
rect 11042 11182 11094 11228
rect 11150 11182 11202 11228
rect 1760 11179 1812 11182
rect 1868 11179 1920 11182
rect 1976 11179 2028 11182
rect 2084 11179 2136 11182
rect 2192 11179 2244 11182
rect 2300 11179 2352 11182
rect 2408 11179 2460 11182
rect 2516 11179 2568 11182
rect 2624 11179 2676 11182
rect 2732 11179 2784 11182
rect 2840 11179 2892 11182
rect 2948 11179 3000 11182
rect 3056 11179 3108 11182
rect 3164 11179 3216 11182
rect 3272 11179 3324 11182
rect 3380 11179 3432 11182
rect 3488 11179 3540 11182
rect 3596 11179 3648 11182
rect 3704 11179 3756 11182
rect 4130 11179 4182 11182
rect 4238 11179 4290 11182
rect 4346 11179 4398 11182
rect 4454 11179 4506 11182
rect 4562 11179 4614 11182
rect 4670 11179 4722 11182
rect 4778 11179 4830 11182
rect 4886 11179 4938 11182
rect 4994 11179 5046 11182
rect 5102 11179 5154 11182
rect 5210 11179 5262 11182
rect 5318 11179 5370 11182
rect 5426 11179 5478 11182
rect 5534 11179 5586 11182
rect 5642 11179 5694 11182
rect 5750 11179 5802 11182
rect 5858 11179 5910 11182
rect 5966 11179 6018 11182
rect 6074 11179 6126 11182
rect 6836 11179 6888 11182
rect 6944 11179 6996 11182
rect 7052 11179 7104 11182
rect 7160 11179 7212 11182
rect 7268 11179 7320 11182
rect 7376 11179 7428 11182
rect 7484 11179 7536 11182
rect 7592 11179 7644 11182
rect 7700 11179 7752 11182
rect 7808 11179 7860 11182
rect 7916 11179 7968 11182
rect 8024 11179 8076 11182
rect 8132 11179 8184 11182
rect 8240 11179 8292 11182
rect 8348 11179 8400 11182
rect 8456 11179 8508 11182
rect 8564 11179 8616 11182
rect 8672 11179 8724 11182
rect 8780 11179 8832 11182
rect 9206 11179 9258 11182
rect 9314 11179 9366 11182
rect 9422 11179 9474 11182
rect 9530 11179 9582 11182
rect 9638 11179 9690 11182
rect 9746 11179 9798 11182
rect 9854 11179 9906 11182
rect 9962 11179 10014 11182
rect 10070 11179 10122 11182
rect 10178 11179 10230 11182
rect 10286 11179 10338 11182
rect 10394 11179 10446 11182
rect 10502 11179 10554 11182
rect 10610 11179 10662 11182
rect 10718 11179 10770 11182
rect 10826 11179 10878 11182
rect 10934 11179 10986 11182
rect 11042 11179 11094 11182
rect 11150 11179 11202 11182
rect 1493 10984 1545 10987
rect 1601 10984 1653 10987
rect 3863 10984 3915 10987
rect 3971 10984 4023 10987
rect 6239 10984 6291 10987
rect 6347 10984 6399 10987
rect 6455 10984 6507 10987
rect 6563 10984 6615 10987
rect 6671 10984 6723 10987
rect 8939 10984 8991 10987
rect 9047 10984 9099 10987
rect 11309 10984 11361 10987
rect 11417 10984 11469 10987
rect 1493 10938 1494 10984
rect 1494 10938 1545 10984
rect 1601 10938 1653 10984
rect 3863 10938 3915 10984
rect 3971 10938 4023 10984
rect 6239 10938 6291 10984
rect 6347 10938 6399 10984
rect 6455 10938 6507 10984
rect 6563 10938 6615 10984
rect 6671 10938 6723 10984
rect 8939 10938 8991 10984
rect 9047 10938 9099 10984
rect 11309 10938 11361 10984
rect 11417 10938 11468 10984
rect 11468 10938 11469 10984
rect 1493 10935 1545 10938
rect 1601 10935 1653 10938
rect 3863 10935 3915 10938
rect 3971 10935 4023 10938
rect 6239 10935 6291 10938
rect 6347 10935 6399 10938
rect 6455 10935 6507 10938
rect 6563 10935 6615 10938
rect 6671 10935 6723 10938
rect 8939 10935 8991 10938
rect 9047 10935 9099 10938
rect 11309 10935 11361 10938
rect 11417 10935 11469 10938
rect 1760 10740 1812 10743
rect 1868 10740 1920 10743
rect 1976 10740 2028 10743
rect 2084 10740 2136 10743
rect 2192 10740 2244 10743
rect 2300 10740 2352 10743
rect 2408 10740 2460 10743
rect 2516 10740 2568 10743
rect 2624 10740 2676 10743
rect 2732 10740 2784 10743
rect 2840 10740 2892 10743
rect 2948 10740 3000 10743
rect 3056 10740 3108 10743
rect 3164 10740 3216 10743
rect 3272 10740 3324 10743
rect 3380 10740 3432 10743
rect 3488 10740 3540 10743
rect 3596 10740 3648 10743
rect 3704 10740 3756 10743
rect 4130 10740 4182 10743
rect 4238 10740 4290 10743
rect 4346 10740 4398 10743
rect 4454 10740 4506 10743
rect 4562 10740 4614 10743
rect 4670 10740 4722 10743
rect 4778 10740 4830 10743
rect 4886 10740 4938 10743
rect 4994 10740 5046 10743
rect 5102 10740 5154 10743
rect 5210 10740 5262 10743
rect 5318 10740 5370 10743
rect 5426 10740 5478 10743
rect 5534 10740 5586 10743
rect 5642 10740 5694 10743
rect 5750 10740 5802 10743
rect 5858 10740 5910 10743
rect 5966 10740 6018 10743
rect 6074 10740 6126 10743
rect 6836 10740 6888 10743
rect 6944 10740 6996 10743
rect 7052 10740 7104 10743
rect 7160 10740 7212 10743
rect 7268 10740 7320 10743
rect 7376 10740 7428 10743
rect 7484 10740 7536 10743
rect 7592 10740 7644 10743
rect 7700 10740 7752 10743
rect 7808 10740 7860 10743
rect 7916 10740 7968 10743
rect 8024 10740 8076 10743
rect 8132 10740 8184 10743
rect 8240 10740 8292 10743
rect 8348 10740 8400 10743
rect 8456 10740 8508 10743
rect 8564 10740 8616 10743
rect 8672 10740 8724 10743
rect 8780 10740 8832 10743
rect 9206 10740 9258 10743
rect 9314 10740 9366 10743
rect 9422 10740 9474 10743
rect 9530 10740 9582 10743
rect 9638 10740 9690 10743
rect 9746 10740 9798 10743
rect 9854 10740 9906 10743
rect 9962 10740 10014 10743
rect 10070 10740 10122 10743
rect 10178 10740 10230 10743
rect 10286 10740 10338 10743
rect 10394 10740 10446 10743
rect 10502 10740 10554 10743
rect 10610 10740 10662 10743
rect 10718 10740 10770 10743
rect 10826 10740 10878 10743
rect 10934 10740 10986 10743
rect 11042 10740 11094 10743
rect 11150 10740 11202 10743
rect 1760 10694 1812 10740
rect 1868 10694 1920 10740
rect 1976 10694 2028 10740
rect 2084 10694 2136 10740
rect 2192 10694 2244 10740
rect 2300 10694 2352 10740
rect 2408 10694 2460 10740
rect 2516 10694 2568 10740
rect 2624 10694 2676 10740
rect 2732 10694 2784 10740
rect 2840 10694 2892 10740
rect 2948 10694 3000 10740
rect 3056 10694 3108 10740
rect 3164 10694 3216 10740
rect 3272 10694 3324 10740
rect 3380 10694 3432 10740
rect 3488 10694 3540 10740
rect 3596 10694 3648 10740
rect 3704 10694 3756 10740
rect 4130 10694 4182 10740
rect 4238 10694 4290 10740
rect 4346 10694 4398 10740
rect 4454 10694 4506 10740
rect 4562 10694 4614 10740
rect 4670 10694 4722 10740
rect 4778 10694 4830 10740
rect 4886 10694 4938 10740
rect 4994 10694 5046 10740
rect 5102 10694 5154 10740
rect 5210 10694 5262 10740
rect 5318 10694 5370 10740
rect 5426 10694 5478 10740
rect 5534 10694 5586 10740
rect 5642 10694 5694 10740
rect 5750 10694 5802 10740
rect 5858 10694 5910 10740
rect 5966 10694 6018 10740
rect 6074 10694 6126 10740
rect 6836 10694 6888 10740
rect 6944 10694 6996 10740
rect 7052 10694 7104 10740
rect 7160 10694 7212 10740
rect 7268 10694 7320 10740
rect 7376 10694 7428 10740
rect 7484 10694 7536 10740
rect 7592 10694 7644 10740
rect 7700 10694 7752 10740
rect 7808 10694 7860 10740
rect 7916 10694 7968 10740
rect 8024 10694 8076 10740
rect 8132 10694 8184 10740
rect 8240 10694 8292 10740
rect 8348 10694 8400 10740
rect 8456 10694 8508 10740
rect 8564 10694 8616 10740
rect 8672 10694 8724 10740
rect 8780 10694 8832 10740
rect 9206 10694 9258 10740
rect 9314 10694 9366 10740
rect 9422 10694 9474 10740
rect 9530 10694 9582 10740
rect 9638 10694 9690 10740
rect 9746 10694 9798 10740
rect 9854 10694 9906 10740
rect 9962 10694 10014 10740
rect 10070 10694 10122 10740
rect 10178 10694 10230 10740
rect 10286 10694 10338 10740
rect 10394 10694 10446 10740
rect 10502 10694 10554 10740
rect 10610 10694 10662 10740
rect 10718 10694 10770 10740
rect 10826 10694 10878 10740
rect 10934 10694 10986 10740
rect 11042 10694 11094 10740
rect 11150 10694 11202 10740
rect 1760 10691 1812 10694
rect 1868 10691 1920 10694
rect 1976 10691 2028 10694
rect 2084 10691 2136 10694
rect 2192 10691 2244 10694
rect 2300 10691 2352 10694
rect 2408 10691 2460 10694
rect 2516 10691 2568 10694
rect 2624 10691 2676 10694
rect 2732 10691 2784 10694
rect 2840 10691 2892 10694
rect 2948 10691 3000 10694
rect 3056 10691 3108 10694
rect 3164 10691 3216 10694
rect 3272 10691 3324 10694
rect 3380 10691 3432 10694
rect 3488 10691 3540 10694
rect 3596 10691 3648 10694
rect 3704 10691 3756 10694
rect 4130 10691 4182 10694
rect 4238 10691 4290 10694
rect 4346 10691 4398 10694
rect 4454 10691 4506 10694
rect 4562 10691 4614 10694
rect 4670 10691 4722 10694
rect 4778 10691 4830 10694
rect 4886 10691 4938 10694
rect 4994 10691 5046 10694
rect 5102 10691 5154 10694
rect 5210 10691 5262 10694
rect 5318 10691 5370 10694
rect 5426 10691 5478 10694
rect 5534 10691 5586 10694
rect 5642 10691 5694 10694
rect 5750 10691 5802 10694
rect 5858 10691 5910 10694
rect 5966 10691 6018 10694
rect 6074 10691 6126 10694
rect 6836 10691 6888 10694
rect 6944 10691 6996 10694
rect 7052 10691 7104 10694
rect 7160 10691 7212 10694
rect 7268 10691 7320 10694
rect 7376 10691 7428 10694
rect 7484 10691 7536 10694
rect 7592 10691 7644 10694
rect 7700 10691 7752 10694
rect 7808 10691 7860 10694
rect 7916 10691 7968 10694
rect 8024 10691 8076 10694
rect 8132 10691 8184 10694
rect 8240 10691 8292 10694
rect 8348 10691 8400 10694
rect 8456 10691 8508 10694
rect 8564 10691 8616 10694
rect 8672 10691 8724 10694
rect 8780 10691 8832 10694
rect 9206 10691 9258 10694
rect 9314 10691 9366 10694
rect 9422 10691 9474 10694
rect 9530 10691 9582 10694
rect 9638 10691 9690 10694
rect 9746 10691 9798 10694
rect 9854 10691 9906 10694
rect 9962 10691 10014 10694
rect 10070 10691 10122 10694
rect 10178 10691 10230 10694
rect 10286 10691 10338 10694
rect 10394 10691 10446 10694
rect 10502 10691 10554 10694
rect 10610 10691 10662 10694
rect 10718 10691 10770 10694
rect 10826 10691 10878 10694
rect 10934 10691 10986 10694
rect 11042 10691 11094 10694
rect 11150 10691 11202 10694
rect 1493 10496 1545 10499
rect 1601 10496 1653 10499
rect 3863 10496 3915 10499
rect 3971 10496 4023 10499
rect 6239 10496 6291 10499
rect 6347 10496 6399 10499
rect 6455 10496 6507 10499
rect 6563 10496 6615 10499
rect 6671 10496 6723 10499
rect 8939 10496 8991 10499
rect 9047 10496 9099 10499
rect 11309 10496 11361 10499
rect 11417 10496 11469 10499
rect 1493 10450 1494 10496
rect 1494 10450 1545 10496
rect 1601 10450 1653 10496
rect 3863 10450 3915 10496
rect 3971 10450 4023 10496
rect 6239 10450 6291 10496
rect 6347 10450 6399 10496
rect 6455 10450 6507 10496
rect 6563 10450 6615 10496
rect 6671 10450 6723 10496
rect 8939 10450 8991 10496
rect 9047 10450 9099 10496
rect 11309 10450 11361 10496
rect 11417 10450 11468 10496
rect 11468 10450 11469 10496
rect 1493 10447 1545 10450
rect 1601 10447 1653 10450
rect 3863 10447 3915 10450
rect 3971 10447 4023 10450
rect 6239 10447 6291 10450
rect 6347 10447 6399 10450
rect 6455 10447 6507 10450
rect 6563 10447 6615 10450
rect 6671 10447 6723 10450
rect 8939 10447 8991 10450
rect 9047 10447 9099 10450
rect 11309 10447 11361 10450
rect 11417 10447 11469 10450
rect 1760 10252 1812 10255
rect 1868 10252 1920 10255
rect 1976 10252 2028 10255
rect 2084 10252 2136 10255
rect 2192 10252 2244 10255
rect 2300 10252 2352 10255
rect 2408 10252 2460 10255
rect 2516 10252 2568 10255
rect 2624 10252 2676 10255
rect 2732 10252 2784 10255
rect 2840 10252 2892 10255
rect 2948 10252 3000 10255
rect 3056 10252 3108 10255
rect 3164 10252 3216 10255
rect 3272 10252 3324 10255
rect 3380 10252 3432 10255
rect 3488 10252 3540 10255
rect 3596 10252 3648 10255
rect 3704 10252 3756 10255
rect 4130 10252 4182 10255
rect 4238 10252 4290 10255
rect 4346 10252 4398 10255
rect 4454 10252 4506 10255
rect 4562 10252 4614 10255
rect 4670 10252 4722 10255
rect 4778 10252 4830 10255
rect 4886 10252 4938 10255
rect 4994 10252 5046 10255
rect 5102 10252 5154 10255
rect 5210 10252 5262 10255
rect 5318 10252 5370 10255
rect 5426 10252 5478 10255
rect 5534 10252 5586 10255
rect 5642 10252 5694 10255
rect 5750 10252 5802 10255
rect 5858 10252 5910 10255
rect 5966 10252 6018 10255
rect 6074 10252 6126 10255
rect 6836 10252 6888 10255
rect 6944 10252 6996 10255
rect 7052 10252 7104 10255
rect 7160 10252 7212 10255
rect 7268 10252 7320 10255
rect 7376 10252 7428 10255
rect 7484 10252 7536 10255
rect 7592 10252 7644 10255
rect 7700 10252 7752 10255
rect 7808 10252 7860 10255
rect 7916 10252 7968 10255
rect 8024 10252 8076 10255
rect 8132 10252 8184 10255
rect 8240 10252 8292 10255
rect 8348 10252 8400 10255
rect 8456 10252 8508 10255
rect 8564 10252 8616 10255
rect 8672 10252 8724 10255
rect 8780 10252 8832 10255
rect 9206 10252 9258 10255
rect 9314 10252 9366 10255
rect 9422 10252 9474 10255
rect 9530 10252 9582 10255
rect 9638 10252 9690 10255
rect 9746 10252 9798 10255
rect 9854 10252 9906 10255
rect 9962 10252 10014 10255
rect 10070 10252 10122 10255
rect 10178 10252 10230 10255
rect 10286 10252 10338 10255
rect 10394 10252 10446 10255
rect 10502 10252 10554 10255
rect 10610 10252 10662 10255
rect 10718 10252 10770 10255
rect 10826 10252 10878 10255
rect 10934 10252 10986 10255
rect 11042 10252 11094 10255
rect 11150 10252 11202 10255
rect 1760 10206 1812 10252
rect 1868 10206 1920 10252
rect 1976 10206 2028 10252
rect 2084 10206 2136 10252
rect 2192 10206 2244 10252
rect 2300 10206 2352 10252
rect 2408 10206 2460 10252
rect 2516 10206 2568 10252
rect 2624 10206 2676 10252
rect 2732 10206 2784 10252
rect 2840 10206 2892 10252
rect 2948 10206 3000 10252
rect 3056 10206 3108 10252
rect 3164 10206 3216 10252
rect 3272 10206 3324 10252
rect 3380 10206 3432 10252
rect 3488 10206 3540 10252
rect 3596 10206 3648 10252
rect 3704 10206 3756 10252
rect 4130 10206 4182 10252
rect 4238 10206 4290 10252
rect 4346 10206 4398 10252
rect 4454 10206 4506 10252
rect 4562 10206 4614 10252
rect 4670 10206 4722 10252
rect 4778 10206 4830 10252
rect 4886 10206 4938 10252
rect 4994 10206 5046 10252
rect 5102 10206 5154 10252
rect 5210 10206 5262 10252
rect 5318 10206 5370 10252
rect 5426 10206 5478 10252
rect 5534 10206 5586 10252
rect 5642 10206 5694 10252
rect 5750 10206 5802 10252
rect 5858 10206 5910 10252
rect 5966 10206 6018 10252
rect 6074 10206 6126 10252
rect 6836 10206 6888 10252
rect 6944 10206 6996 10252
rect 7052 10206 7104 10252
rect 7160 10206 7212 10252
rect 7268 10206 7320 10252
rect 7376 10206 7428 10252
rect 7484 10206 7536 10252
rect 7592 10206 7644 10252
rect 7700 10206 7752 10252
rect 7808 10206 7860 10252
rect 7916 10206 7968 10252
rect 8024 10206 8076 10252
rect 8132 10206 8184 10252
rect 8240 10206 8292 10252
rect 8348 10206 8400 10252
rect 8456 10206 8508 10252
rect 8564 10206 8616 10252
rect 8672 10206 8724 10252
rect 8780 10206 8832 10252
rect 9206 10206 9258 10252
rect 9314 10206 9366 10252
rect 9422 10206 9474 10252
rect 9530 10206 9582 10252
rect 9638 10206 9690 10252
rect 9746 10206 9798 10252
rect 9854 10206 9906 10252
rect 9962 10206 10014 10252
rect 10070 10206 10122 10252
rect 10178 10206 10230 10252
rect 10286 10206 10338 10252
rect 10394 10206 10446 10252
rect 10502 10206 10554 10252
rect 10610 10206 10662 10252
rect 10718 10206 10770 10252
rect 10826 10206 10878 10252
rect 10934 10206 10986 10252
rect 11042 10206 11094 10252
rect 11150 10206 11202 10252
rect 1760 10203 1812 10206
rect 1868 10203 1920 10206
rect 1976 10203 2028 10206
rect 2084 10203 2136 10206
rect 2192 10203 2244 10206
rect 2300 10203 2352 10206
rect 2408 10203 2460 10206
rect 2516 10203 2568 10206
rect 2624 10203 2676 10206
rect 2732 10203 2784 10206
rect 2840 10203 2892 10206
rect 2948 10203 3000 10206
rect 3056 10203 3108 10206
rect 3164 10203 3216 10206
rect 3272 10203 3324 10206
rect 3380 10203 3432 10206
rect 3488 10203 3540 10206
rect 3596 10203 3648 10206
rect 3704 10203 3756 10206
rect 4130 10203 4182 10206
rect 4238 10203 4290 10206
rect 4346 10203 4398 10206
rect 4454 10203 4506 10206
rect 4562 10203 4614 10206
rect 4670 10203 4722 10206
rect 4778 10203 4830 10206
rect 4886 10203 4938 10206
rect 4994 10203 5046 10206
rect 5102 10203 5154 10206
rect 5210 10203 5262 10206
rect 5318 10203 5370 10206
rect 5426 10203 5478 10206
rect 5534 10203 5586 10206
rect 5642 10203 5694 10206
rect 5750 10203 5802 10206
rect 5858 10203 5910 10206
rect 5966 10203 6018 10206
rect 6074 10203 6126 10206
rect 6836 10203 6888 10206
rect 6944 10203 6996 10206
rect 7052 10203 7104 10206
rect 7160 10203 7212 10206
rect 7268 10203 7320 10206
rect 7376 10203 7428 10206
rect 7484 10203 7536 10206
rect 7592 10203 7644 10206
rect 7700 10203 7752 10206
rect 7808 10203 7860 10206
rect 7916 10203 7968 10206
rect 8024 10203 8076 10206
rect 8132 10203 8184 10206
rect 8240 10203 8292 10206
rect 8348 10203 8400 10206
rect 8456 10203 8508 10206
rect 8564 10203 8616 10206
rect 8672 10203 8724 10206
rect 8780 10203 8832 10206
rect 9206 10203 9258 10206
rect 9314 10203 9366 10206
rect 9422 10203 9474 10206
rect 9530 10203 9582 10206
rect 9638 10203 9690 10206
rect 9746 10203 9798 10206
rect 9854 10203 9906 10206
rect 9962 10203 10014 10206
rect 10070 10203 10122 10206
rect 10178 10203 10230 10206
rect 10286 10203 10338 10206
rect 10394 10203 10446 10206
rect 10502 10203 10554 10206
rect 10610 10203 10662 10206
rect 10718 10203 10770 10206
rect 10826 10203 10878 10206
rect 10934 10203 10986 10206
rect 11042 10203 11094 10206
rect 11150 10203 11202 10206
rect 1493 10008 1545 10011
rect 1601 10008 1653 10011
rect 3863 10008 3915 10011
rect 3971 10008 4023 10011
rect 6239 10008 6291 10011
rect 6347 10008 6399 10011
rect 6455 10008 6507 10011
rect 6563 10008 6615 10011
rect 6671 10008 6723 10011
rect 8939 10008 8991 10011
rect 9047 10008 9099 10011
rect 11309 10008 11361 10011
rect 11417 10008 11469 10011
rect 1493 9962 1494 10008
rect 1494 9962 1545 10008
rect 1601 9962 1653 10008
rect 3863 9962 3915 10008
rect 3971 9962 4023 10008
rect 6239 9962 6291 10008
rect 6347 9962 6399 10008
rect 6455 9962 6507 10008
rect 6563 9962 6615 10008
rect 6671 9962 6723 10008
rect 8939 9962 8991 10008
rect 9047 9962 9099 10008
rect 11309 9962 11361 10008
rect 11417 9962 11468 10008
rect 11468 9962 11469 10008
rect 1493 9959 1545 9962
rect 1601 9959 1653 9962
rect 3863 9959 3915 9962
rect 3971 9959 4023 9962
rect 6239 9959 6291 9962
rect 6347 9959 6399 9962
rect 6455 9959 6507 9962
rect 6563 9959 6615 9962
rect 6671 9959 6723 9962
rect 8939 9959 8991 9962
rect 9047 9959 9099 9962
rect 11309 9959 11361 9962
rect 11417 9959 11469 9962
rect 1760 9764 1812 9767
rect 1868 9764 1920 9767
rect 1976 9764 2028 9767
rect 2084 9764 2136 9767
rect 2192 9764 2244 9767
rect 2300 9764 2352 9767
rect 2408 9764 2460 9767
rect 2516 9764 2568 9767
rect 2624 9764 2676 9767
rect 2732 9764 2784 9767
rect 2840 9764 2892 9767
rect 2948 9764 3000 9767
rect 3056 9764 3108 9767
rect 3164 9764 3216 9767
rect 3272 9764 3324 9767
rect 3380 9764 3432 9767
rect 3488 9764 3540 9767
rect 3596 9764 3648 9767
rect 3704 9764 3756 9767
rect 4130 9764 4182 9767
rect 4238 9764 4290 9767
rect 4346 9764 4398 9767
rect 4454 9764 4506 9767
rect 4562 9764 4614 9767
rect 4670 9764 4722 9767
rect 4778 9764 4830 9767
rect 4886 9764 4938 9767
rect 4994 9764 5046 9767
rect 5102 9764 5154 9767
rect 5210 9764 5262 9767
rect 5318 9764 5370 9767
rect 5426 9764 5478 9767
rect 5534 9764 5586 9767
rect 5642 9764 5694 9767
rect 5750 9764 5802 9767
rect 5858 9764 5910 9767
rect 5966 9764 6018 9767
rect 6074 9764 6126 9767
rect 6836 9764 6888 9767
rect 6944 9764 6996 9767
rect 7052 9764 7104 9767
rect 7160 9764 7212 9767
rect 7268 9764 7320 9767
rect 7376 9764 7428 9767
rect 7484 9764 7536 9767
rect 7592 9764 7644 9767
rect 7700 9764 7752 9767
rect 7808 9764 7860 9767
rect 7916 9764 7968 9767
rect 8024 9764 8076 9767
rect 8132 9764 8184 9767
rect 8240 9764 8292 9767
rect 8348 9764 8400 9767
rect 8456 9764 8508 9767
rect 8564 9764 8616 9767
rect 8672 9764 8724 9767
rect 8780 9764 8832 9767
rect 9206 9764 9258 9767
rect 9314 9764 9366 9767
rect 9422 9764 9474 9767
rect 9530 9764 9582 9767
rect 9638 9764 9690 9767
rect 9746 9764 9798 9767
rect 9854 9764 9906 9767
rect 9962 9764 10014 9767
rect 10070 9764 10122 9767
rect 10178 9764 10230 9767
rect 10286 9764 10338 9767
rect 10394 9764 10446 9767
rect 10502 9764 10554 9767
rect 10610 9764 10662 9767
rect 10718 9764 10770 9767
rect 10826 9764 10878 9767
rect 10934 9764 10986 9767
rect 11042 9764 11094 9767
rect 11150 9764 11202 9767
rect 1760 9718 1812 9764
rect 1868 9718 1920 9764
rect 1976 9718 2028 9764
rect 2084 9718 2136 9764
rect 2192 9718 2244 9764
rect 2300 9718 2352 9764
rect 2408 9718 2460 9764
rect 2516 9718 2568 9764
rect 2624 9718 2676 9764
rect 2732 9718 2784 9764
rect 2840 9718 2892 9764
rect 2948 9718 3000 9764
rect 3056 9718 3108 9764
rect 3164 9718 3216 9764
rect 3272 9718 3324 9764
rect 3380 9718 3432 9764
rect 3488 9718 3540 9764
rect 3596 9718 3648 9764
rect 3704 9718 3756 9764
rect 4130 9718 4182 9764
rect 4238 9718 4290 9764
rect 4346 9718 4398 9764
rect 4454 9718 4506 9764
rect 4562 9718 4614 9764
rect 4670 9718 4722 9764
rect 4778 9718 4830 9764
rect 4886 9718 4938 9764
rect 4994 9718 5046 9764
rect 5102 9718 5154 9764
rect 5210 9718 5262 9764
rect 5318 9718 5370 9764
rect 5426 9718 5478 9764
rect 5534 9718 5586 9764
rect 5642 9718 5694 9764
rect 5750 9718 5802 9764
rect 5858 9718 5910 9764
rect 5966 9718 6018 9764
rect 6074 9718 6126 9764
rect 6836 9718 6888 9764
rect 6944 9718 6996 9764
rect 7052 9718 7104 9764
rect 7160 9718 7212 9764
rect 7268 9718 7320 9764
rect 7376 9718 7428 9764
rect 7484 9718 7536 9764
rect 7592 9718 7644 9764
rect 7700 9718 7752 9764
rect 7808 9718 7860 9764
rect 7916 9718 7968 9764
rect 8024 9718 8076 9764
rect 8132 9718 8184 9764
rect 8240 9718 8292 9764
rect 8348 9718 8400 9764
rect 8456 9718 8508 9764
rect 8564 9718 8616 9764
rect 8672 9718 8724 9764
rect 8780 9718 8832 9764
rect 9206 9718 9258 9764
rect 9314 9718 9366 9764
rect 9422 9718 9474 9764
rect 9530 9718 9582 9764
rect 9638 9718 9690 9764
rect 9746 9718 9798 9764
rect 9854 9718 9906 9764
rect 9962 9718 10014 9764
rect 10070 9718 10122 9764
rect 10178 9718 10230 9764
rect 10286 9718 10338 9764
rect 10394 9718 10446 9764
rect 10502 9718 10554 9764
rect 10610 9718 10662 9764
rect 10718 9718 10770 9764
rect 10826 9718 10878 9764
rect 10934 9718 10986 9764
rect 11042 9718 11094 9764
rect 11150 9718 11202 9764
rect 1760 9715 1812 9718
rect 1868 9715 1920 9718
rect 1976 9715 2028 9718
rect 2084 9715 2136 9718
rect 2192 9715 2244 9718
rect 2300 9715 2352 9718
rect 2408 9715 2460 9718
rect 2516 9715 2568 9718
rect 2624 9715 2676 9718
rect 2732 9715 2784 9718
rect 2840 9715 2892 9718
rect 2948 9715 3000 9718
rect 3056 9715 3108 9718
rect 3164 9715 3216 9718
rect 3272 9715 3324 9718
rect 3380 9715 3432 9718
rect 3488 9715 3540 9718
rect 3596 9715 3648 9718
rect 3704 9715 3756 9718
rect 4130 9715 4182 9718
rect 4238 9715 4290 9718
rect 4346 9715 4398 9718
rect 4454 9715 4506 9718
rect 4562 9715 4614 9718
rect 4670 9715 4722 9718
rect 4778 9715 4830 9718
rect 4886 9715 4938 9718
rect 4994 9715 5046 9718
rect 5102 9715 5154 9718
rect 5210 9715 5262 9718
rect 5318 9715 5370 9718
rect 5426 9715 5478 9718
rect 5534 9715 5586 9718
rect 5642 9715 5694 9718
rect 5750 9715 5802 9718
rect 5858 9715 5910 9718
rect 5966 9715 6018 9718
rect 6074 9715 6126 9718
rect 6836 9715 6888 9718
rect 6944 9715 6996 9718
rect 7052 9715 7104 9718
rect 7160 9715 7212 9718
rect 7268 9715 7320 9718
rect 7376 9715 7428 9718
rect 7484 9715 7536 9718
rect 7592 9715 7644 9718
rect 7700 9715 7752 9718
rect 7808 9715 7860 9718
rect 7916 9715 7968 9718
rect 8024 9715 8076 9718
rect 8132 9715 8184 9718
rect 8240 9715 8292 9718
rect 8348 9715 8400 9718
rect 8456 9715 8508 9718
rect 8564 9715 8616 9718
rect 8672 9715 8724 9718
rect 8780 9715 8832 9718
rect 9206 9715 9258 9718
rect 9314 9715 9366 9718
rect 9422 9715 9474 9718
rect 9530 9715 9582 9718
rect 9638 9715 9690 9718
rect 9746 9715 9798 9718
rect 9854 9715 9906 9718
rect 9962 9715 10014 9718
rect 10070 9715 10122 9718
rect 10178 9715 10230 9718
rect 10286 9715 10338 9718
rect 10394 9715 10446 9718
rect 10502 9715 10554 9718
rect 10610 9715 10662 9718
rect 10718 9715 10770 9718
rect 10826 9715 10878 9718
rect 10934 9715 10986 9718
rect 11042 9715 11094 9718
rect 11150 9715 11202 9718
rect 1493 9520 1545 9523
rect 1601 9520 1653 9523
rect 3863 9520 3915 9523
rect 3971 9520 4023 9523
rect 6239 9520 6291 9523
rect 6347 9520 6399 9523
rect 6455 9520 6507 9523
rect 6563 9520 6615 9523
rect 6671 9520 6723 9523
rect 8939 9520 8991 9523
rect 9047 9520 9099 9523
rect 11309 9520 11361 9523
rect 11417 9520 11469 9523
rect 1493 9474 1494 9520
rect 1494 9474 1545 9520
rect 1601 9474 1653 9520
rect 3863 9474 3915 9520
rect 3971 9474 4023 9520
rect 6239 9474 6291 9520
rect 6347 9474 6399 9520
rect 6455 9474 6507 9520
rect 6563 9474 6615 9520
rect 6671 9474 6723 9520
rect 8939 9474 8991 9520
rect 9047 9474 9099 9520
rect 11309 9474 11361 9520
rect 11417 9474 11468 9520
rect 11468 9474 11469 9520
rect 1493 9471 1545 9474
rect 1601 9471 1653 9474
rect 3863 9471 3915 9474
rect 3971 9471 4023 9474
rect 6239 9471 6291 9474
rect 6347 9471 6399 9474
rect 6455 9471 6507 9474
rect 6563 9471 6615 9474
rect 6671 9471 6723 9474
rect 8939 9471 8991 9474
rect 9047 9471 9099 9474
rect 11309 9471 11361 9474
rect 11417 9471 11469 9474
rect 1760 9276 1812 9279
rect 1868 9276 1920 9279
rect 1976 9276 2028 9279
rect 2084 9276 2136 9279
rect 2192 9276 2244 9279
rect 2300 9276 2352 9279
rect 2408 9276 2460 9279
rect 2516 9276 2568 9279
rect 2624 9276 2676 9279
rect 2732 9276 2784 9279
rect 2840 9276 2892 9279
rect 2948 9276 3000 9279
rect 3056 9276 3108 9279
rect 3164 9276 3216 9279
rect 3272 9276 3324 9279
rect 3380 9276 3432 9279
rect 3488 9276 3540 9279
rect 3596 9276 3648 9279
rect 3704 9276 3756 9279
rect 4130 9276 4182 9279
rect 4238 9276 4290 9279
rect 4346 9276 4398 9279
rect 4454 9276 4506 9279
rect 4562 9276 4614 9279
rect 4670 9276 4722 9279
rect 4778 9276 4830 9279
rect 4886 9276 4938 9279
rect 4994 9276 5046 9279
rect 5102 9276 5154 9279
rect 5210 9276 5262 9279
rect 5318 9276 5370 9279
rect 5426 9276 5478 9279
rect 5534 9276 5586 9279
rect 5642 9276 5694 9279
rect 5750 9276 5802 9279
rect 5858 9276 5910 9279
rect 5966 9276 6018 9279
rect 6074 9276 6126 9279
rect 6836 9276 6888 9279
rect 6944 9276 6996 9279
rect 7052 9276 7104 9279
rect 7160 9276 7212 9279
rect 7268 9276 7320 9279
rect 7376 9276 7428 9279
rect 7484 9276 7536 9279
rect 7592 9276 7644 9279
rect 7700 9276 7752 9279
rect 7808 9276 7860 9279
rect 7916 9276 7968 9279
rect 8024 9276 8076 9279
rect 8132 9276 8184 9279
rect 8240 9276 8292 9279
rect 8348 9276 8400 9279
rect 8456 9276 8508 9279
rect 8564 9276 8616 9279
rect 8672 9276 8724 9279
rect 8780 9276 8832 9279
rect 9206 9276 9258 9279
rect 9314 9276 9366 9279
rect 9422 9276 9474 9279
rect 9530 9276 9582 9279
rect 9638 9276 9690 9279
rect 9746 9276 9798 9279
rect 9854 9276 9906 9279
rect 9962 9276 10014 9279
rect 10070 9276 10122 9279
rect 10178 9276 10230 9279
rect 10286 9276 10338 9279
rect 10394 9276 10446 9279
rect 10502 9276 10554 9279
rect 10610 9276 10662 9279
rect 10718 9276 10770 9279
rect 10826 9276 10878 9279
rect 10934 9276 10986 9279
rect 11042 9276 11094 9279
rect 11150 9276 11202 9279
rect 1760 9230 1812 9276
rect 1868 9230 1920 9276
rect 1976 9230 2028 9276
rect 2084 9230 2136 9276
rect 2192 9230 2244 9276
rect 2300 9230 2352 9276
rect 2408 9230 2460 9276
rect 2516 9230 2568 9276
rect 2624 9230 2676 9276
rect 2732 9230 2784 9276
rect 2840 9230 2892 9276
rect 2948 9230 3000 9276
rect 3056 9230 3108 9276
rect 3164 9230 3216 9276
rect 3272 9230 3324 9276
rect 3380 9230 3432 9276
rect 3488 9230 3540 9276
rect 3596 9230 3648 9276
rect 3704 9230 3756 9276
rect 4130 9230 4182 9276
rect 4238 9230 4290 9276
rect 4346 9230 4398 9276
rect 4454 9230 4506 9276
rect 4562 9230 4614 9276
rect 4670 9230 4722 9276
rect 4778 9230 4830 9276
rect 4886 9230 4938 9276
rect 4994 9230 5046 9276
rect 5102 9230 5154 9276
rect 5210 9230 5262 9276
rect 5318 9230 5370 9276
rect 5426 9230 5478 9276
rect 5534 9230 5586 9276
rect 5642 9230 5694 9276
rect 5750 9230 5802 9276
rect 5858 9230 5910 9276
rect 5966 9230 6018 9276
rect 6074 9230 6126 9276
rect 6836 9230 6888 9276
rect 6944 9230 6996 9276
rect 7052 9230 7104 9276
rect 7160 9230 7212 9276
rect 7268 9230 7320 9276
rect 7376 9230 7428 9276
rect 7484 9230 7536 9276
rect 7592 9230 7644 9276
rect 7700 9230 7752 9276
rect 7808 9230 7860 9276
rect 7916 9230 7968 9276
rect 8024 9230 8076 9276
rect 8132 9230 8184 9276
rect 8240 9230 8292 9276
rect 8348 9230 8400 9276
rect 8456 9230 8508 9276
rect 8564 9230 8616 9276
rect 8672 9230 8724 9276
rect 8780 9230 8832 9276
rect 9206 9230 9258 9276
rect 9314 9230 9366 9276
rect 9422 9230 9474 9276
rect 9530 9230 9582 9276
rect 9638 9230 9690 9276
rect 9746 9230 9798 9276
rect 9854 9230 9906 9276
rect 9962 9230 10014 9276
rect 10070 9230 10122 9276
rect 10178 9230 10230 9276
rect 10286 9230 10338 9276
rect 10394 9230 10446 9276
rect 10502 9230 10554 9276
rect 10610 9230 10662 9276
rect 10718 9230 10770 9276
rect 10826 9230 10878 9276
rect 10934 9230 10986 9276
rect 11042 9230 11094 9276
rect 11150 9230 11202 9276
rect 1760 9227 1812 9230
rect 1868 9227 1920 9230
rect 1976 9227 2028 9230
rect 2084 9227 2136 9230
rect 2192 9227 2244 9230
rect 2300 9227 2352 9230
rect 2408 9227 2460 9230
rect 2516 9227 2568 9230
rect 2624 9227 2676 9230
rect 2732 9227 2784 9230
rect 2840 9227 2892 9230
rect 2948 9227 3000 9230
rect 3056 9227 3108 9230
rect 3164 9227 3216 9230
rect 3272 9227 3324 9230
rect 3380 9227 3432 9230
rect 3488 9227 3540 9230
rect 3596 9227 3648 9230
rect 3704 9227 3756 9230
rect 4130 9227 4182 9230
rect 4238 9227 4290 9230
rect 4346 9227 4398 9230
rect 4454 9227 4506 9230
rect 4562 9227 4614 9230
rect 4670 9227 4722 9230
rect 4778 9227 4830 9230
rect 4886 9227 4938 9230
rect 4994 9227 5046 9230
rect 5102 9227 5154 9230
rect 5210 9227 5262 9230
rect 5318 9227 5370 9230
rect 5426 9227 5478 9230
rect 5534 9227 5586 9230
rect 5642 9227 5694 9230
rect 5750 9227 5802 9230
rect 5858 9227 5910 9230
rect 5966 9227 6018 9230
rect 6074 9227 6126 9230
rect 6836 9227 6888 9230
rect 6944 9227 6996 9230
rect 7052 9227 7104 9230
rect 7160 9227 7212 9230
rect 7268 9227 7320 9230
rect 7376 9227 7428 9230
rect 7484 9227 7536 9230
rect 7592 9227 7644 9230
rect 7700 9227 7752 9230
rect 7808 9227 7860 9230
rect 7916 9227 7968 9230
rect 8024 9227 8076 9230
rect 8132 9227 8184 9230
rect 8240 9227 8292 9230
rect 8348 9227 8400 9230
rect 8456 9227 8508 9230
rect 8564 9227 8616 9230
rect 8672 9227 8724 9230
rect 8780 9227 8832 9230
rect 9206 9227 9258 9230
rect 9314 9227 9366 9230
rect 9422 9227 9474 9230
rect 9530 9227 9582 9230
rect 9638 9227 9690 9230
rect 9746 9227 9798 9230
rect 9854 9227 9906 9230
rect 9962 9227 10014 9230
rect 10070 9227 10122 9230
rect 10178 9227 10230 9230
rect 10286 9227 10338 9230
rect 10394 9227 10446 9230
rect 10502 9227 10554 9230
rect 10610 9227 10662 9230
rect 10718 9227 10770 9230
rect 10826 9227 10878 9230
rect 10934 9227 10986 9230
rect 11042 9227 11094 9230
rect 11150 9227 11202 9230
rect 1493 9032 1545 9035
rect 1601 9032 1653 9035
rect 3863 9032 3915 9035
rect 3971 9032 4023 9035
rect 6239 9032 6291 9035
rect 6347 9032 6399 9035
rect 6455 9032 6507 9035
rect 6563 9032 6615 9035
rect 6671 9032 6723 9035
rect 8939 9032 8991 9035
rect 9047 9032 9099 9035
rect 11309 9032 11361 9035
rect 11417 9032 11469 9035
rect 1493 8986 1494 9032
rect 1494 8986 1545 9032
rect 1601 8986 1653 9032
rect 3863 8986 3915 9032
rect 3971 8986 4023 9032
rect 6239 8986 6291 9032
rect 6347 8986 6399 9032
rect 6455 8986 6507 9032
rect 6563 8986 6615 9032
rect 6671 8986 6723 9032
rect 8939 8986 8991 9032
rect 9047 8986 9099 9032
rect 11309 8986 11361 9032
rect 11417 8986 11468 9032
rect 11468 8986 11469 9032
rect 1493 8983 1545 8986
rect 1601 8983 1653 8986
rect 3863 8983 3915 8986
rect 3971 8983 4023 8986
rect 6239 8983 6291 8986
rect 6347 8983 6399 8986
rect 6455 8983 6507 8986
rect 6563 8983 6615 8986
rect 6671 8983 6723 8986
rect 8939 8983 8991 8986
rect 9047 8983 9099 8986
rect 11309 8983 11361 8986
rect 11417 8983 11469 8986
rect 1760 8788 1812 8791
rect 1868 8788 1920 8791
rect 1976 8788 2028 8791
rect 2084 8788 2136 8791
rect 2192 8788 2244 8791
rect 2300 8788 2352 8791
rect 2408 8788 2460 8791
rect 2516 8788 2568 8791
rect 2624 8788 2676 8791
rect 2732 8788 2784 8791
rect 2840 8788 2892 8791
rect 2948 8788 3000 8791
rect 3056 8788 3108 8791
rect 3164 8788 3216 8791
rect 3272 8788 3324 8791
rect 3380 8788 3432 8791
rect 3488 8788 3540 8791
rect 3596 8788 3648 8791
rect 3704 8788 3756 8791
rect 4130 8788 4182 8791
rect 4238 8788 4290 8791
rect 4346 8788 4398 8791
rect 4454 8788 4506 8791
rect 4562 8788 4614 8791
rect 4670 8788 4722 8791
rect 4778 8788 4830 8791
rect 4886 8788 4938 8791
rect 4994 8788 5046 8791
rect 5102 8788 5154 8791
rect 5210 8788 5262 8791
rect 5318 8788 5370 8791
rect 5426 8788 5478 8791
rect 5534 8788 5586 8791
rect 5642 8788 5694 8791
rect 5750 8788 5802 8791
rect 5858 8788 5910 8791
rect 5966 8788 6018 8791
rect 6074 8788 6126 8791
rect 6836 8788 6888 8791
rect 6944 8788 6996 8791
rect 7052 8788 7104 8791
rect 7160 8788 7212 8791
rect 7268 8788 7320 8791
rect 7376 8788 7428 8791
rect 7484 8788 7536 8791
rect 7592 8788 7644 8791
rect 7700 8788 7752 8791
rect 7808 8788 7860 8791
rect 7916 8788 7968 8791
rect 8024 8788 8076 8791
rect 8132 8788 8184 8791
rect 8240 8788 8292 8791
rect 8348 8788 8400 8791
rect 8456 8788 8508 8791
rect 8564 8788 8616 8791
rect 8672 8788 8724 8791
rect 8780 8788 8832 8791
rect 9206 8788 9258 8791
rect 9314 8788 9366 8791
rect 9422 8788 9474 8791
rect 9530 8788 9582 8791
rect 9638 8788 9690 8791
rect 9746 8788 9798 8791
rect 9854 8788 9906 8791
rect 9962 8788 10014 8791
rect 10070 8788 10122 8791
rect 10178 8788 10230 8791
rect 10286 8788 10338 8791
rect 10394 8788 10446 8791
rect 10502 8788 10554 8791
rect 10610 8788 10662 8791
rect 10718 8788 10770 8791
rect 10826 8788 10878 8791
rect 10934 8788 10986 8791
rect 11042 8788 11094 8791
rect 11150 8788 11202 8791
rect 1760 8742 1812 8788
rect 1868 8742 1920 8788
rect 1976 8742 2028 8788
rect 2084 8742 2136 8788
rect 2192 8742 2244 8788
rect 2300 8742 2352 8788
rect 2408 8742 2460 8788
rect 2516 8742 2568 8788
rect 2624 8742 2676 8788
rect 2732 8742 2784 8788
rect 2840 8742 2892 8788
rect 2948 8742 3000 8788
rect 3056 8742 3108 8788
rect 3164 8742 3216 8788
rect 3272 8742 3324 8788
rect 3380 8742 3432 8788
rect 3488 8742 3540 8788
rect 3596 8742 3648 8788
rect 3704 8742 3756 8788
rect 4130 8742 4182 8788
rect 4238 8742 4290 8788
rect 4346 8742 4398 8788
rect 4454 8742 4506 8788
rect 4562 8742 4614 8788
rect 4670 8742 4722 8788
rect 4778 8742 4830 8788
rect 4886 8742 4938 8788
rect 4994 8742 5046 8788
rect 5102 8742 5154 8788
rect 5210 8742 5262 8788
rect 5318 8742 5370 8788
rect 5426 8742 5478 8788
rect 5534 8742 5586 8788
rect 5642 8742 5694 8788
rect 5750 8742 5802 8788
rect 5858 8742 5910 8788
rect 5966 8742 6018 8788
rect 6074 8742 6126 8788
rect 6836 8742 6888 8788
rect 6944 8742 6996 8788
rect 7052 8742 7104 8788
rect 7160 8742 7212 8788
rect 7268 8742 7320 8788
rect 7376 8742 7428 8788
rect 7484 8742 7536 8788
rect 7592 8742 7644 8788
rect 7700 8742 7752 8788
rect 7808 8742 7860 8788
rect 7916 8742 7968 8788
rect 8024 8742 8076 8788
rect 8132 8742 8184 8788
rect 8240 8742 8292 8788
rect 8348 8742 8400 8788
rect 8456 8742 8508 8788
rect 8564 8742 8616 8788
rect 8672 8742 8724 8788
rect 8780 8742 8832 8788
rect 9206 8742 9258 8788
rect 9314 8742 9366 8788
rect 9422 8742 9474 8788
rect 9530 8742 9582 8788
rect 9638 8742 9690 8788
rect 9746 8742 9798 8788
rect 9854 8742 9906 8788
rect 9962 8742 10014 8788
rect 10070 8742 10122 8788
rect 10178 8742 10230 8788
rect 10286 8742 10338 8788
rect 10394 8742 10446 8788
rect 10502 8742 10554 8788
rect 10610 8742 10662 8788
rect 10718 8742 10770 8788
rect 10826 8742 10878 8788
rect 10934 8742 10986 8788
rect 11042 8742 11094 8788
rect 11150 8742 11202 8788
rect 1760 8739 1812 8742
rect 1868 8739 1920 8742
rect 1976 8739 2028 8742
rect 2084 8739 2136 8742
rect 2192 8739 2244 8742
rect 2300 8739 2352 8742
rect 2408 8739 2460 8742
rect 2516 8739 2568 8742
rect 2624 8739 2676 8742
rect 2732 8739 2784 8742
rect 2840 8739 2892 8742
rect 2948 8739 3000 8742
rect 3056 8739 3108 8742
rect 3164 8739 3216 8742
rect 3272 8739 3324 8742
rect 3380 8739 3432 8742
rect 3488 8739 3540 8742
rect 3596 8739 3648 8742
rect 3704 8739 3756 8742
rect 4130 8739 4182 8742
rect 4238 8739 4290 8742
rect 4346 8739 4398 8742
rect 4454 8739 4506 8742
rect 4562 8739 4614 8742
rect 4670 8739 4722 8742
rect 4778 8739 4830 8742
rect 4886 8739 4938 8742
rect 4994 8739 5046 8742
rect 5102 8739 5154 8742
rect 5210 8739 5262 8742
rect 5318 8739 5370 8742
rect 5426 8739 5478 8742
rect 5534 8739 5586 8742
rect 5642 8739 5694 8742
rect 5750 8739 5802 8742
rect 5858 8739 5910 8742
rect 5966 8739 6018 8742
rect 6074 8739 6126 8742
rect 6836 8739 6888 8742
rect 6944 8739 6996 8742
rect 7052 8739 7104 8742
rect 7160 8739 7212 8742
rect 7268 8739 7320 8742
rect 7376 8739 7428 8742
rect 7484 8739 7536 8742
rect 7592 8739 7644 8742
rect 7700 8739 7752 8742
rect 7808 8739 7860 8742
rect 7916 8739 7968 8742
rect 8024 8739 8076 8742
rect 8132 8739 8184 8742
rect 8240 8739 8292 8742
rect 8348 8739 8400 8742
rect 8456 8739 8508 8742
rect 8564 8739 8616 8742
rect 8672 8739 8724 8742
rect 8780 8739 8832 8742
rect 9206 8739 9258 8742
rect 9314 8739 9366 8742
rect 9422 8739 9474 8742
rect 9530 8739 9582 8742
rect 9638 8739 9690 8742
rect 9746 8739 9798 8742
rect 9854 8739 9906 8742
rect 9962 8739 10014 8742
rect 10070 8739 10122 8742
rect 10178 8739 10230 8742
rect 10286 8739 10338 8742
rect 10394 8739 10446 8742
rect 10502 8739 10554 8742
rect 10610 8739 10662 8742
rect 10718 8739 10770 8742
rect 10826 8739 10878 8742
rect 10934 8739 10986 8742
rect 11042 8739 11094 8742
rect 11150 8739 11202 8742
rect 1493 8544 1545 8547
rect 1601 8544 1653 8547
rect 3863 8544 3915 8547
rect 3971 8544 4023 8547
rect 6239 8544 6291 8547
rect 6347 8544 6399 8547
rect 6455 8544 6507 8547
rect 6563 8544 6615 8547
rect 6671 8544 6723 8547
rect 8939 8544 8991 8547
rect 9047 8544 9099 8547
rect 11309 8544 11361 8547
rect 11417 8544 11469 8547
rect 1493 8498 1494 8544
rect 1494 8498 1545 8544
rect 1601 8498 1653 8544
rect 3863 8498 3915 8544
rect 3971 8498 4023 8544
rect 6239 8498 6291 8544
rect 6347 8498 6399 8544
rect 6455 8498 6507 8544
rect 6563 8498 6615 8544
rect 6671 8498 6723 8544
rect 8939 8498 8991 8544
rect 9047 8498 9099 8544
rect 11309 8498 11361 8544
rect 11417 8498 11468 8544
rect 11468 8498 11469 8544
rect 1493 8495 1545 8498
rect 1601 8495 1653 8498
rect 3863 8495 3915 8498
rect 3971 8495 4023 8498
rect 6239 8495 6291 8498
rect 6347 8495 6399 8498
rect 6455 8495 6507 8498
rect 6563 8495 6615 8498
rect 6671 8495 6723 8498
rect 8939 8495 8991 8498
rect 9047 8495 9099 8498
rect 11309 8495 11361 8498
rect 11417 8495 11469 8498
rect 1760 8300 1812 8303
rect 1868 8300 1920 8303
rect 1976 8300 2028 8303
rect 2084 8300 2136 8303
rect 2192 8300 2244 8303
rect 2300 8300 2352 8303
rect 2408 8300 2460 8303
rect 2516 8300 2568 8303
rect 2624 8300 2676 8303
rect 2732 8300 2784 8303
rect 2840 8300 2892 8303
rect 2948 8300 3000 8303
rect 3056 8300 3108 8303
rect 3164 8300 3216 8303
rect 3272 8300 3324 8303
rect 3380 8300 3432 8303
rect 3488 8300 3540 8303
rect 3596 8300 3648 8303
rect 3704 8300 3756 8303
rect 4130 8300 4182 8303
rect 4238 8300 4290 8303
rect 4346 8300 4398 8303
rect 4454 8300 4506 8303
rect 4562 8300 4614 8303
rect 4670 8300 4722 8303
rect 4778 8300 4830 8303
rect 4886 8300 4938 8303
rect 4994 8300 5046 8303
rect 5102 8300 5154 8303
rect 5210 8300 5262 8303
rect 5318 8300 5370 8303
rect 5426 8300 5478 8303
rect 5534 8300 5586 8303
rect 5642 8300 5694 8303
rect 5750 8300 5802 8303
rect 5858 8300 5910 8303
rect 5966 8300 6018 8303
rect 6074 8300 6126 8303
rect 6836 8300 6888 8303
rect 6944 8300 6996 8303
rect 7052 8300 7104 8303
rect 7160 8300 7212 8303
rect 7268 8300 7320 8303
rect 7376 8300 7428 8303
rect 7484 8300 7536 8303
rect 7592 8300 7644 8303
rect 7700 8300 7752 8303
rect 7808 8300 7860 8303
rect 7916 8300 7968 8303
rect 8024 8300 8076 8303
rect 8132 8300 8184 8303
rect 8240 8300 8292 8303
rect 8348 8300 8400 8303
rect 8456 8300 8508 8303
rect 8564 8300 8616 8303
rect 8672 8300 8724 8303
rect 8780 8300 8832 8303
rect 9206 8300 9258 8303
rect 9314 8300 9366 8303
rect 9422 8300 9474 8303
rect 9530 8300 9582 8303
rect 9638 8300 9690 8303
rect 9746 8300 9798 8303
rect 9854 8300 9906 8303
rect 9962 8300 10014 8303
rect 10070 8300 10122 8303
rect 10178 8300 10230 8303
rect 10286 8300 10338 8303
rect 10394 8300 10446 8303
rect 10502 8300 10554 8303
rect 10610 8300 10662 8303
rect 10718 8300 10770 8303
rect 10826 8300 10878 8303
rect 10934 8300 10986 8303
rect 11042 8300 11094 8303
rect 11150 8300 11202 8303
rect 1760 8254 1812 8300
rect 1868 8254 1920 8300
rect 1976 8254 2028 8300
rect 2084 8254 2136 8300
rect 2192 8254 2244 8300
rect 2300 8254 2352 8300
rect 2408 8254 2460 8300
rect 2516 8254 2568 8300
rect 2624 8254 2676 8300
rect 2732 8254 2784 8300
rect 2840 8254 2892 8300
rect 2948 8254 3000 8300
rect 3056 8254 3108 8300
rect 3164 8254 3216 8300
rect 3272 8254 3324 8300
rect 3380 8254 3432 8300
rect 3488 8254 3540 8300
rect 3596 8254 3648 8300
rect 3704 8254 3756 8300
rect 4130 8254 4182 8300
rect 4238 8254 4290 8300
rect 4346 8254 4398 8300
rect 4454 8254 4506 8300
rect 4562 8254 4614 8300
rect 4670 8254 4722 8300
rect 4778 8254 4830 8300
rect 4886 8254 4938 8300
rect 4994 8254 5046 8300
rect 5102 8254 5154 8300
rect 5210 8254 5262 8300
rect 5318 8254 5370 8300
rect 5426 8254 5478 8300
rect 5534 8254 5586 8300
rect 5642 8254 5694 8300
rect 5750 8254 5802 8300
rect 5858 8254 5910 8300
rect 5966 8254 6018 8300
rect 6074 8254 6126 8300
rect 6836 8254 6888 8300
rect 6944 8254 6996 8300
rect 7052 8254 7104 8300
rect 7160 8254 7212 8300
rect 7268 8254 7320 8300
rect 7376 8254 7428 8300
rect 7484 8254 7536 8300
rect 7592 8254 7644 8300
rect 7700 8254 7752 8300
rect 7808 8254 7860 8300
rect 7916 8254 7968 8300
rect 8024 8254 8076 8300
rect 8132 8254 8184 8300
rect 8240 8254 8292 8300
rect 8348 8254 8400 8300
rect 8456 8254 8508 8300
rect 8564 8254 8616 8300
rect 8672 8254 8724 8300
rect 8780 8254 8832 8300
rect 9206 8254 9258 8300
rect 9314 8254 9366 8300
rect 9422 8254 9474 8300
rect 9530 8254 9582 8300
rect 9638 8254 9690 8300
rect 9746 8254 9798 8300
rect 9854 8254 9906 8300
rect 9962 8254 10014 8300
rect 10070 8254 10122 8300
rect 10178 8254 10230 8300
rect 10286 8254 10338 8300
rect 10394 8254 10446 8300
rect 10502 8254 10554 8300
rect 10610 8254 10662 8300
rect 10718 8254 10770 8300
rect 10826 8254 10878 8300
rect 10934 8254 10986 8300
rect 11042 8254 11094 8300
rect 11150 8254 11202 8300
rect 1760 8251 1812 8254
rect 1868 8251 1920 8254
rect 1976 8251 2028 8254
rect 2084 8251 2136 8254
rect 2192 8251 2244 8254
rect 2300 8251 2352 8254
rect 2408 8251 2460 8254
rect 2516 8251 2568 8254
rect 2624 8251 2676 8254
rect 2732 8251 2784 8254
rect 2840 8251 2892 8254
rect 2948 8251 3000 8254
rect 3056 8251 3108 8254
rect 3164 8251 3216 8254
rect 3272 8251 3324 8254
rect 3380 8251 3432 8254
rect 3488 8251 3540 8254
rect 3596 8251 3648 8254
rect 3704 8251 3756 8254
rect 4130 8251 4182 8254
rect 4238 8251 4290 8254
rect 4346 8251 4398 8254
rect 4454 8251 4506 8254
rect 4562 8251 4614 8254
rect 4670 8251 4722 8254
rect 4778 8251 4830 8254
rect 4886 8251 4938 8254
rect 4994 8251 5046 8254
rect 5102 8251 5154 8254
rect 5210 8251 5262 8254
rect 5318 8251 5370 8254
rect 5426 8251 5478 8254
rect 5534 8251 5586 8254
rect 5642 8251 5694 8254
rect 5750 8251 5802 8254
rect 5858 8251 5910 8254
rect 5966 8251 6018 8254
rect 6074 8251 6126 8254
rect 6836 8251 6888 8254
rect 6944 8251 6996 8254
rect 7052 8251 7104 8254
rect 7160 8251 7212 8254
rect 7268 8251 7320 8254
rect 7376 8251 7428 8254
rect 7484 8251 7536 8254
rect 7592 8251 7644 8254
rect 7700 8251 7752 8254
rect 7808 8251 7860 8254
rect 7916 8251 7968 8254
rect 8024 8251 8076 8254
rect 8132 8251 8184 8254
rect 8240 8251 8292 8254
rect 8348 8251 8400 8254
rect 8456 8251 8508 8254
rect 8564 8251 8616 8254
rect 8672 8251 8724 8254
rect 8780 8251 8832 8254
rect 9206 8251 9258 8254
rect 9314 8251 9366 8254
rect 9422 8251 9474 8254
rect 9530 8251 9582 8254
rect 9638 8251 9690 8254
rect 9746 8251 9798 8254
rect 9854 8251 9906 8254
rect 9962 8251 10014 8254
rect 10070 8251 10122 8254
rect 10178 8251 10230 8254
rect 10286 8251 10338 8254
rect 10394 8251 10446 8254
rect 10502 8251 10554 8254
rect 10610 8251 10662 8254
rect 10718 8251 10770 8254
rect 10826 8251 10878 8254
rect 10934 8251 10986 8254
rect 11042 8251 11094 8254
rect 11150 8251 11202 8254
rect 1493 8056 1545 8059
rect 1601 8056 1653 8059
rect 3863 8056 3915 8059
rect 3971 8056 4023 8059
rect 6239 8056 6291 8059
rect 6347 8056 6399 8059
rect 6455 8056 6507 8059
rect 6563 8056 6615 8059
rect 6671 8056 6723 8059
rect 8939 8056 8991 8059
rect 9047 8056 9099 8059
rect 11309 8056 11361 8059
rect 11417 8056 11469 8059
rect 1493 8010 1494 8056
rect 1494 8010 1545 8056
rect 1601 8010 1653 8056
rect 3863 8010 3915 8056
rect 3971 8010 4023 8056
rect 6239 8010 6291 8056
rect 6347 8010 6399 8056
rect 6455 8010 6507 8056
rect 6563 8010 6615 8056
rect 6671 8010 6723 8056
rect 8939 8010 8991 8056
rect 9047 8010 9099 8056
rect 11309 8010 11361 8056
rect 11417 8010 11468 8056
rect 11468 8010 11469 8056
rect 1493 8007 1545 8010
rect 1601 8007 1653 8010
rect 3863 8007 3915 8010
rect 3971 8007 4023 8010
rect 6239 8007 6291 8010
rect 6347 8007 6399 8010
rect 6455 8007 6507 8010
rect 6563 8007 6615 8010
rect 6671 8007 6723 8010
rect 8939 8007 8991 8010
rect 9047 8007 9099 8010
rect 11309 8007 11361 8010
rect 11417 8007 11469 8010
rect 1760 7812 1812 7815
rect 1868 7812 1920 7815
rect 1976 7812 2028 7815
rect 2084 7812 2136 7815
rect 2192 7812 2244 7815
rect 2300 7812 2352 7815
rect 2408 7812 2460 7815
rect 2516 7812 2568 7815
rect 2624 7812 2676 7815
rect 2732 7812 2784 7815
rect 2840 7812 2892 7815
rect 2948 7812 3000 7815
rect 3056 7812 3108 7815
rect 3164 7812 3216 7815
rect 3272 7812 3324 7815
rect 3380 7812 3432 7815
rect 3488 7812 3540 7815
rect 3596 7812 3648 7815
rect 3704 7812 3756 7815
rect 4130 7812 4182 7815
rect 4238 7812 4290 7815
rect 4346 7812 4398 7815
rect 4454 7812 4506 7815
rect 4562 7812 4614 7815
rect 4670 7812 4722 7815
rect 4778 7812 4830 7815
rect 4886 7812 4938 7815
rect 4994 7812 5046 7815
rect 5102 7812 5154 7815
rect 5210 7812 5262 7815
rect 5318 7812 5370 7815
rect 5426 7812 5478 7815
rect 5534 7812 5586 7815
rect 5642 7812 5694 7815
rect 5750 7812 5802 7815
rect 5858 7812 5910 7815
rect 5966 7812 6018 7815
rect 6074 7812 6126 7815
rect 6836 7812 6888 7815
rect 6944 7812 6996 7815
rect 7052 7812 7104 7815
rect 7160 7812 7212 7815
rect 7268 7812 7320 7815
rect 7376 7812 7428 7815
rect 7484 7812 7536 7815
rect 7592 7812 7644 7815
rect 7700 7812 7752 7815
rect 7808 7812 7860 7815
rect 7916 7812 7968 7815
rect 8024 7812 8076 7815
rect 8132 7812 8184 7815
rect 8240 7812 8292 7815
rect 8348 7812 8400 7815
rect 8456 7812 8508 7815
rect 8564 7812 8616 7815
rect 8672 7812 8724 7815
rect 8780 7812 8832 7815
rect 9206 7812 9258 7815
rect 9314 7812 9366 7815
rect 9422 7812 9474 7815
rect 9530 7812 9582 7815
rect 9638 7812 9690 7815
rect 9746 7812 9798 7815
rect 9854 7812 9906 7815
rect 9962 7812 10014 7815
rect 10070 7812 10122 7815
rect 10178 7812 10230 7815
rect 10286 7812 10338 7815
rect 10394 7812 10446 7815
rect 10502 7812 10554 7815
rect 10610 7812 10662 7815
rect 10718 7812 10770 7815
rect 10826 7812 10878 7815
rect 10934 7812 10986 7815
rect 11042 7812 11094 7815
rect 11150 7812 11202 7815
rect 1760 7766 1812 7812
rect 1868 7766 1920 7812
rect 1976 7766 2028 7812
rect 2084 7766 2136 7812
rect 2192 7766 2244 7812
rect 2300 7766 2352 7812
rect 2408 7766 2460 7812
rect 2516 7766 2568 7812
rect 2624 7766 2676 7812
rect 2732 7766 2784 7812
rect 2840 7766 2892 7812
rect 2948 7766 3000 7812
rect 3056 7766 3108 7812
rect 3164 7766 3216 7812
rect 3272 7766 3324 7812
rect 3380 7766 3432 7812
rect 3488 7766 3540 7812
rect 3596 7766 3648 7812
rect 3704 7766 3756 7812
rect 4130 7766 4182 7812
rect 4238 7766 4290 7812
rect 4346 7766 4398 7812
rect 4454 7766 4506 7812
rect 4562 7766 4614 7812
rect 4670 7766 4722 7812
rect 4778 7766 4830 7812
rect 4886 7766 4938 7812
rect 4994 7766 5046 7812
rect 5102 7766 5154 7812
rect 5210 7766 5262 7812
rect 5318 7766 5370 7812
rect 5426 7766 5478 7812
rect 5534 7766 5586 7812
rect 5642 7766 5694 7812
rect 5750 7766 5802 7812
rect 5858 7766 5910 7812
rect 5966 7766 6018 7812
rect 6074 7766 6126 7812
rect 6836 7766 6888 7812
rect 6944 7766 6996 7812
rect 7052 7766 7104 7812
rect 7160 7766 7212 7812
rect 7268 7766 7320 7812
rect 7376 7766 7428 7812
rect 7484 7766 7536 7812
rect 7592 7766 7644 7812
rect 7700 7766 7752 7812
rect 7808 7766 7860 7812
rect 7916 7766 7968 7812
rect 8024 7766 8076 7812
rect 8132 7766 8184 7812
rect 8240 7766 8292 7812
rect 8348 7766 8400 7812
rect 8456 7766 8508 7812
rect 8564 7766 8616 7812
rect 8672 7766 8724 7812
rect 8780 7766 8832 7812
rect 9206 7766 9258 7812
rect 9314 7766 9366 7812
rect 9422 7766 9474 7812
rect 9530 7766 9582 7812
rect 9638 7766 9690 7812
rect 9746 7766 9798 7812
rect 9854 7766 9906 7812
rect 9962 7766 10014 7812
rect 10070 7766 10122 7812
rect 10178 7766 10230 7812
rect 10286 7766 10338 7812
rect 10394 7766 10446 7812
rect 10502 7766 10554 7812
rect 10610 7766 10662 7812
rect 10718 7766 10770 7812
rect 10826 7766 10878 7812
rect 10934 7766 10986 7812
rect 11042 7766 11094 7812
rect 11150 7766 11202 7812
rect 1760 7763 1812 7766
rect 1868 7763 1920 7766
rect 1976 7763 2028 7766
rect 2084 7763 2136 7766
rect 2192 7763 2244 7766
rect 2300 7763 2352 7766
rect 2408 7763 2460 7766
rect 2516 7763 2568 7766
rect 2624 7763 2676 7766
rect 2732 7763 2784 7766
rect 2840 7763 2892 7766
rect 2948 7763 3000 7766
rect 3056 7763 3108 7766
rect 3164 7763 3216 7766
rect 3272 7763 3324 7766
rect 3380 7763 3432 7766
rect 3488 7763 3540 7766
rect 3596 7763 3648 7766
rect 3704 7763 3756 7766
rect 4130 7763 4182 7766
rect 4238 7763 4290 7766
rect 4346 7763 4398 7766
rect 4454 7763 4506 7766
rect 4562 7763 4614 7766
rect 4670 7763 4722 7766
rect 4778 7763 4830 7766
rect 4886 7763 4938 7766
rect 4994 7763 5046 7766
rect 5102 7763 5154 7766
rect 5210 7763 5262 7766
rect 5318 7763 5370 7766
rect 5426 7763 5478 7766
rect 5534 7763 5586 7766
rect 5642 7763 5694 7766
rect 5750 7763 5802 7766
rect 5858 7763 5910 7766
rect 5966 7763 6018 7766
rect 6074 7763 6126 7766
rect 6836 7763 6888 7766
rect 6944 7763 6996 7766
rect 7052 7763 7104 7766
rect 7160 7763 7212 7766
rect 7268 7763 7320 7766
rect 7376 7763 7428 7766
rect 7484 7763 7536 7766
rect 7592 7763 7644 7766
rect 7700 7763 7752 7766
rect 7808 7763 7860 7766
rect 7916 7763 7968 7766
rect 8024 7763 8076 7766
rect 8132 7763 8184 7766
rect 8240 7763 8292 7766
rect 8348 7763 8400 7766
rect 8456 7763 8508 7766
rect 8564 7763 8616 7766
rect 8672 7763 8724 7766
rect 8780 7763 8832 7766
rect 9206 7763 9258 7766
rect 9314 7763 9366 7766
rect 9422 7763 9474 7766
rect 9530 7763 9582 7766
rect 9638 7763 9690 7766
rect 9746 7763 9798 7766
rect 9854 7763 9906 7766
rect 9962 7763 10014 7766
rect 10070 7763 10122 7766
rect 10178 7763 10230 7766
rect 10286 7763 10338 7766
rect 10394 7763 10446 7766
rect 10502 7763 10554 7766
rect 10610 7763 10662 7766
rect 10718 7763 10770 7766
rect 10826 7763 10878 7766
rect 10934 7763 10986 7766
rect 11042 7763 11094 7766
rect 11150 7763 11202 7766
rect 1493 7568 1545 7571
rect 1601 7568 1653 7571
rect 3863 7568 3915 7571
rect 3971 7568 4023 7571
rect 6239 7568 6291 7571
rect 6347 7568 6399 7571
rect 6455 7568 6507 7571
rect 6563 7568 6615 7571
rect 6671 7568 6723 7571
rect 8939 7568 8991 7571
rect 9047 7568 9099 7571
rect 11309 7568 11361 7571
rect 11417 7568 11469 7571
rect 1493 7522 1494 7568
rect 1494 7522 1545 7568
rect 1601 7522 1653 7568
rect 3863 7522 3915 7568
rect 3971 7522 4023 7568
rect 6239 7522 6291 7568
rect 6347 7522 6399 7568
rect 6455 7522 6507 7568
rect 6563 7522 6615 7568
rect 6671 7522 6723 7568
rect 8939 7522 8991 7568
rect 9047 7522 9099 7568
rect 11309 7522 11361 7568
rect 11417 7522 11468 7568
rect 11468 7522 11469 7568
rect 1493 7519 1545 7522
rect 1601 7519 1653 7522
rect 3863 7519 3915 7522
rect 3971 7519 4023 7522
rect 6239 7519 6291 7522
rect 6347 7519 6399 7522
rect 6455 7519 6507 7522
rect 6563 7519 6615 7522
rect 6671 7519 6723 7522
rect 8939 7519 8991 7522
rect 9047 7519 9099 7522
rect 11309 7519 11361 7522
rect 11417 7519 11469 7522
rect 1233 7339 1285 7391
rect 1341 7339 1393 7391
rect 11569 11983 11621 12035
rect 11677 11983 11706 12035
rect 11706 11983 11729 12035
rect 11569 11875 11621 11927
rect 11677 11875 11706 11927
rect 11706 11875 11729 11927
rect 11569 11767 11621 11819
rect 11677 11767 11706 11819
rect 11706 11767 11729 11819
rect 11569 11659 11621 11711
rect 11677 11659 11706 11711
rect 11706 11659 11729 11711
rect 11569 11551 11621 11603
rect 11677 11551 11706 11603
rect 11706 11551 11729 11603
rect 11569 11443 11621 11495
rect 11677 11443 11706 11495
rect 11706 11443 11729 11495
rect 11569 11335 11621 11387
rect 11677 11335 11706 11387
rect 11706 11335 11729 11387
rect 11569 11227 11621 11279
rect 11677 11227 11706 11279
rect 11706 11227 11729 11279
rect 11569 11119 11621 11171
rect 11677 11119 11706 11171
rect 11706 11119 11729 11171
rect 11569 11011 11621 11063
rect 11677 11011 11706 11063
rect 11706 11011 11729 11063
rect 11569 10903 11621 10955
rect 11677 10903 11706 10955
rect 11706 10903 11729 10955
rect 11569 10795 11621 10847
rect 11677 10795 11706 10847
rect 11706 10795 11729 10847
rect 11569 10687 11621 10739
rect 11677 10687 11706 10739
rect 11706 10687 11729 10739
rect 11569 10579 11621 10631
rect 11677 10579 11706 10631
rect 11706 10579 11729 10631
rect 11569 10471 11621 10523
rect 11677 10471 11706 10523
rect 11706 10471 11729 10523
rect 11569 10363 11621 10415
rect 11677 10363 11706 10415
rect 11706 10363 11729 10415
rect 11569 10255 11621 10307
rect 11677 10255 11706 10307
rect 11706 10255 11729 10307
rect 11569 10147 11621 10199
rect 11677 10147 11706 10199
rect 11706 10147 11729 10199
rect 11569 10039 11621 10091
rect 11677 10039 11706 10091
rect 11706 10039 11729 10091
rect 11569 9931 11621 9983
rect 11677 9931 11706 9983
rect 11706 9931 11729 9983
rect 11569 9823 11621 9875
rect 11677 9823 11706 9875
rect 11706 9823 11729 9875
rect 11569 9715 11621 9767
rect 11677 9715 11706 9767
rect 11706 9715 11729 9767
rect 11569 9607 11621 9659
rect 11677 9607 11706 9659
rect 11706 9607 11729 9659
rect 11569 9499 11621 9551
rect 11677 9499 11706 9551
rect 11706 9499 11729 9551
rect 11569 9391 11621 9443
rect 11677 9391 11706 9443
rect 11706 9391 11729 9443
rect 11569 9283 11621 9335
rect 11677 9283 11706 9335
rect 11706 9283 11729 9335
rect 11569 9175 11621 9227
rect 11677 9175 11706 9227
rect 11706 9175 11729 9227
rect 11569 9067 11621 9119
rect 11677 9067 11706 9119
rect 11706 9067 11729 9119
rect 11569 8959 11621 9011
rect 11677 8959 11706 9011
rect 11706 8959 11729 9011
rect 11569 8851 11621 8903
rect 11677 8851 11706 8903
rect 11706 8851 11729 8903
rect 11569 8743 11621 8795
rect 11677 8743 11706 8795
rect 11706 8743 11729 8795
rect 11569 8635 11621 8687
rect 11677 8635 11706 8687
rect 11706 8635 11729 8687
rect 11569 8527 11621 8579
rect 11677 8527 11706 8579
rect 11706 8527 11729 8579
rect 11569 8419 11621 8471
rect 11677 8419 11706 8471
rect 11706 8419 11729 8471
rect 11569 8311 11621 8363
rect 11677 8311 11706 8363
rect 11706 8311 11729 8363
rect 11569 8203 11621 8255
rect 11677 8203 11706 8255
rect 11706 8203 11729 8255
rect 11569 8095 11621 8147
rect 11677 8095 11706 8147
rect 11706 8095 11729 8147
rect 11569 7987 11621 8039
rect 11677 7987 11706 8039
rect 11706 7987 11729 8039
rect 11569 7879 11621 7931
rect 11677 7879 11706 7931
rect 11706 7879 11729 7931
rect 11569 7771 11621 7823
rect 11677 7771 11706 7823
rect 11706 7771 11729 7823
rect 11569 7663 11621 7715
rect 11677 7663 11706 7715
rect 11706 7663 11729 7715
rect 11569 7555 11621 7607
rect 11677 7555 11706 7607
rect 11706 7555 11729 7607
rect 11569 7447 11621 7499
rect 11677 7447 11706 7499
rect 11706 7447 11729 7499
rect 11569 7339 11621 7391
rect 11677 7339 11729 7391
rect 1760 7324 1812 7327
rect 1868 7324 1920 7327
rect 1976 7324 2028 7327
rect 2084 7324 2136 7327
rect 2192 7324 2244 7327
rect 2300 7324 2352 7327
rect 2408 7324 2460 7327
rect 2516 7324 2568 7327
rect 2624 7324 2676 7327
rect 2732 7324 2784 7327
rect 2840 7324 2892 7327
rect 2948 7324 3000 7327
rect 3056 7324 3108 7327
rect 3164 7324 3216 7327
rect 3272 7324 3324 7327
rect 3380 7324 3432 7327
rect 3488 7324 3540 7327
rect 3596 7324 3648 7327
rect 3704 7324 3756 7327
rect 4130 7324 4182 7327
rect 4238 7324 4290 7327
rect 4346 7324 4398 7327
rect 4454 7324 4506 7327
rect 4562 7324 4614 7327
rect 4670 7324 4722 7327
rect 4778 7324 4830 7327
rect 4886 7324 4938 7327
rect 4994 7324 5046 7327
rect 5102 7324 5154 7327
rect 5210 7324 5262 7327
rect 5318 7324 5370 7327
rect 5426 7324 5478 7327
rect 5534 7324 5586 7327
rect 5642 7324 5694 7327
rect 5750 7324 5802 7327
rect 5858 7324 5910 7327
rect 5966 7324 6018 7327
rect 6074 7324 6126 7327
rect 6836 7324 6888 7327
rect 6944 7324 6996 7327
rect 7052 7324 7104 7327
rect 7160 7324 7212 7327
rect 7268 7324 7320 7327
rect 7376 7324 7428 7327
rect 7484 7324 7536 7327
rect 7592 7324 7644 7327
rect 7700 7324 7752 7327
rect 7808 7324 7860 7327
rect 7916 7324 7968 7327
rect 8024 7324 8076 7327
rect 8132 7324 8184 7327
rect 8240 7324 8292 7327
rect 8348 7324 8400 7327
rect 8456 7324 8508 7327
rect 8564 7324 8616 7327
rect 8672 7324 8724 7327
rect 8780 7324 8832 7327
rect 9206 7324 9258 7327
rect 9314 7324 9366 7327
rect 9422 7324 9474 7327
rect 9530 7324 9582 7327
rect 9638 7324 9690 7327
rect 9746 7324 9798 7327
rect 9854 7324 9906 7327
rect 9962 7324 10014 7327
rect 10070 7324 10122 7327
rect 10178 7324 10230 7327
rect 10286 7324 10338 7327
rect 10394 7324 10446 7327
rect 10502 7324 10554 7327
rect 10610 7324 10662 7327
rect 10718 7324 10770 7327
rect 10826 7324 10878 7327
rect 10934 7324 10986 7327
rect 11042 7324 11094 7327
rect 11150 7324 11202 7327
rect 1760 7278 1812 7324
rect 1868 7278 1920 7324
rect 1976 7278 2028 7324
rect 2084 7278 2136 7324
rect 2192 7278 2244 7324
rect 2300 7278 2352 7324
rect 2408 7278 2460 7324
rect 2516 7278 2568 7324
rect 2624 7278 2676 7324
rect 2732 7278 2784 7324
rect 2840 7278 2892 7324
rect 2948 7278 3000 7324
rect 3056 7278 3108 7324
rect 3164 7278 3216 7324
rect 3272 7278 3324 7324
rect 3380 7278 3432 7324
rect 3488 7278 3540 7324
rect 3596 7278 3648 7324
rect 3704 7278 3756 7324
rect 4130 7278 4182 7324
rect 4238 7278 4290 7324
rect 4346 7278 4398 7324
rect 4454 7278 4506 7324
rect 4562 7278 4614 7324
rect 4670 7278 4722 7324
rect 4778 7278 4830 7324
rect 4886 7278 4938 7324
rect 4994 7278 5046 7324
rect 5102 7278 5154 7324
rect 5210 7278 5262 7324
rect 5318 7278 5370 7324
rect 5426 7278 5478 7324
rect 5534 7278 5586 7324
rect 5642 7278 5694 7324
rect 5750 7278 5802 7324
rect 5858 7278 5910 7324
rect 5966 7278 6018 7324
rect 6074 7278 6126 7324
rect 6836 7278 6888 7324
rect 6944 7278 6996 7324
rect 7052 7278 7104 7324
rect 7160 7278 7212 7324
rect 7268 7278 7320 7324
rect 7376 7278 7428 7324
rect 7484 7278 7536 7324
rect 7592 7278 7644 7324
rect 7700 7278 7752 7324
rect 7808 7278 7860 7324
rect 7916 7278 7968 7324
rect 8024 7278 8076 7324
rect 8132 7278 8184 7324
rect 8240 7278 8292 7324
rect 8348 7278 8400 7324
rect 8456 7278 8508 7324
rect 8564 7278 8616 7324
rect 8672 7278 8724 7324
rect 8780 7278 8832 7324
rect 9206 7278 9258 7324
rect 9314 7278 9366 7324
rect 9422 7278 9474 7324
rect 9530 7278 9582 7324
rect 9638 7278 9690 7324
rect 9746 7278 9798 7324
rect 9854 7278 9906 7324
rect 9962 7278 10014 7324
rect 10070 7278 10122 7324
rect 10178 7278 10230 7324
rect 10286 7278 10338 7324
rect 10394 7278 10446 7324
rect 10502 7278 10554 7324
rect 10610 7278 10662 7324
rect 10718 7278 10770 7324
rect 10826 7278 10878 7324
rect 10934 7278 10986 7324
rect 11042 7278 11094 7324
rect 11150 7278 11202 7324
rect 1760 7275 1812 7278
rect 1868 7275 1920 7278
rect 1976 7275 2028 7278
rect 2084 7275 2136 7278
rect 2192 7275 2244 7278
rect 2300 7275 2352 7278
rect 2408 7275 2460 7278
rect 2516 7275 2568 7278
rect 2624 7275 2676 7278
rect 2732 7275 2784 7278
rect 2840 7275 2892 7278
rect 2948 7275 3000 7278
rect 3056 7275 3108 7278
rect 3164 7275 3216 7278
rect 3272 7275 3324 7278
rect 3380 7275 3432 7278
rect 3488 7275 3540 7278
rect 3596 7275 3648 7278
rect 3704 7275 3756 7278
rect 4130 7275 4182 7278
rect 4238 7275 4290 7278
rect 4346 7275 4398 7278
rect 4454 7275 4506 7278
rect 4562 7275 4614 7278
rect 4670 7275 4722 7278
rect 4778 7275 4830 7278
rect 4886 7275 4938 7278
rect 4994 7275 5046 7278
rect 5102 7275 5154 7278
rect 5210 7275 5262 7278
rect 5318 7275 5370 7278
rect 5426 7275 5478 7278
rect 5534 7275 5586 7278
rect 5642 7275 5694 7278
rect 5750 7275 5802 7278
rect 5858 7275 5910 7278
rect 5966 7275 6018 7278
rect 6074 7275 6126 7278
rect 6836 7275 6888 7278
rect 6944 7275 6996 7278
rect 7052 7275 7104 7278
rect 7160 7275 7212 7278
rect 7268 7275 7320 7278
rect 7376 7275 7428 7278
rect 7484 7275 7536 7278
rect 7592 7275 7644 7278
rect 7700 7275 7752 7278
rect 7808 7275 7860 7278
rect 7916 7275 7968 7278
rect 8024 7275 8076 7278
rect 8132 7275 8184 7278
rect 8240 7275 8292 7278
rect 8348 7275 8400 7278
rect 8456 7275 8508 7278
rect 8564 7275 8616 7278
rect 8672 7275 8724 7278
rect 8780 7275 8832 7278
rect 9206 7275 9258 7278
rect 9314 7275 9366 7278
rect 9422 7275 9474 7278
rect 9530 7275 9582 7278
rect 9638 7275 9690 7278
rect 9746 7275 9798 7278
rect 9854 7275 9906 7278
rect 9962 7275 10014 7278
rect 10070 7275 10122 7278
rect 10178 7275 10230 7278
rect 10286 7275 10338 7278
rect 10394 7275 10446 7278
rect 10502 7275 10554 7278
rect 10610 7275 10662 7278
rect 10718 7275 10770 7278
rect 10826 7275 10878 7278
rect 10934 7275 10986 7278
rect 11042 7275 11094 7278
rect 11150 7275 11202 7278
rect 12051 12543 12103 12595
rect 12159 12543 12211 12595
rect 12267 12543 12319 12595
rect 12051 12435 12103 12487
rect 12159 12435 12211 12487
rect 12267 12435 12319 12487
rect 12051 12327 12103 12379
rect 12159 12327 12211 12379
rect 12267 12327 12319 12379
rect 12051 12219 12103 12271
rect 12159 12219 12211 12271
rect 12267 12219 12319 12271
rect 12051 12111 12103 12163
rect 12159 12111 12211 12163
rect 12267 12111 12319 12163
rect 12051 12003 12103 12055
rect 12159 12003 12211 12055
rect 12267 12003 12319 12055
rect 12051 11895 12103 11947
rect 12159 11895 12211 11947
rect 12267 11895 12319 11947
rect 12051 11787 12103 11839
rect 12159 11787 12211 11839
rect 12267 11787 12319 11839
rect 12051 11679 12103 11731
rect 12159 11679 12211 11731
rect 12267 11679 12319 11731
rect 12051 11571 12103 11623
rect 12159 11571 12211 11623
rect 12267 11571 12319 11623
rect 12051 11463 12103 11515
rect 12159 11463 12211 11515
rect 12267 11463 12319 11515
rect 12051 11355 12103 11407
rect 12159 11355 12211 11407
rect 12267 11355 12319 11407
rect 12051 11247 12103 11299
rect 12159 11247 12211 11299
rect 12267 11247 12319 11299
rect 12051 11139 12103 11191
rect 12159 11139 12211 11191
rect 12267 11139 12319 11191
rect 12051 11031 12103 11083
rect 12159 11031 12211 11083
rect 12267 11031 12319 11083
rect 12051 10923 12103 10975
rect 12159 10923 12211 10975
rect 12267 10923 12319 10975
rect 12051 10815 12103 10867
rect 12159 10815 12211 10867
rect 12267 10815 12319 10867
rect 12051 10707 12103 10759
rect 12159 10707 12211 10759
rect 12267 10707 12319 10759
rect 12051 10599 12103 10651
rect 12159 10599 12211 10651
rect 12267 10599 12319 10651
rect 12051 10491 12103 10543
rect 12159 10491 12211 10543
rect 12267 10491 12319 10543
rect 12051 10383 12103 10435
rect 12159 10383 12211 10435
rect 12267 10383 12319 10435
rect 12051 10275 12103 10327
rect 12159 10275 12211 10327
rect 12267 10275 12319 10327
rect 12051 10167 12103 10219
rect 12159 10167 12211 10219
rect 12267 10167 12319 10219
rect 12051 10059 12103 10111
rect 12159 10059 12211 10111
rect 12267 10059 12319 10111
rect 12051 9951 12103 10003
rect 12159 9951 12211 10003
rect 12267 9951 12319 10003
rect 12051 9843 12103 9895
rect 12159 9843 12211 9895
rect 12267 9843 12319 9895
rect 12051 9735 12103 9787
rect 12159 9735 12211 9787
rect 12267 9735 12319 9787
rect 12051 9627 12103 9679
rect 12159 9627 12211 9679
rect 12267 9627 12319 9679
rect 12051 9519 12103 9571
rect 12159 9519 12211 9571
rect 12267 9519 12319 9571
rect 12051 9411 12103 9463
rect 12159 9411 12211 9463
rect 12267 9411 12319 9463
rect 12051 9303 12103 9355
rect 12159 9303 12211 9355
rect 12267 9303 12319 9355
rect 12051 9195 12103 9247
rect 12159 9195 12211 9247
rect 12267 9195 12319 9247
rect 12051 9087 12103 9139
rect 12159 9087 12211 9139
rect 12267 9087 12319 9139
rect 12051 8979 12103 9031
rect 12159 8979 12211 9031
rect 12267 8979 12319 9031
rect 12051 8871 12103 8923
rect 12159 8871 12211 8923
rect 12267 8871 12319 8923
rect 12051 8763 12103 8815
rect 12159 8763 12211 8815
rect 12267 8763 12319 8815
rect 12051 8655 12103 8707
rect 12159 8655 12211 8707
rect 12267 8655 12319 8707
rect 12051 8547 12103 8599
rect 12159 8547 12211 8599
rect 12267 8547 12319 8599
rect 12051 8439 12103 8491
rect 12159 8439 12211 8491
rect 12267 8439 12319 8491
rect 12051 8331 12103 8383
rect 12159 8331 12211 8383
rect 12267 8331 12319 8383
rect 12051 8223 12103 8275
rect 12159 8223 12211 8275
rect 12267 8223 12319 8275
rect 12051 8115 12103 8167
rect 12159 8115 12211 8167
rect 12267 8115 12319 8167
rect 12051 8007 12103 8059
rect 12159 8007 12211 8059
rect 12267 8007 12319 8059
rect 12051 7899 12103 7951
rect 12159 7899 12211 7951
rect 12267 7899 12319 7951
rect 12051 7791 12103 7843
rect 12159 7791 12211 7843
rect 12267 7791 12319 7843
rect 12051 7683 12103 7735
rect 12159 7683 12211 7735
rect 12267 7683 12319 7735
rect 12051 7575 12103 7627
rect 12159 7575 12211 7627
rect 12267 7575 12319 7627
rect 12051 7467 12103 7519
rect 12159 7467 12211 7519
rect 12267 7467 12319 7519
rect 12051 7359 12103 7411
rect 12159 7359 12211 7411
rect 12267 7359 12319 7411
rect 12051 7251 12103 7303
rect 12159 7251 12211 7303
rect 12267 7251 12319 7303
rect 12051 7143 12103 7195
rect 12159 7143 12211 7195
rect 12267 7143 12319 7195
rect 12051 7035 12103 7087
rect 12159 7035 12211 7087
rect 12267 7035 12319 7087
rect 12051 6927 12103 6979
rect 12159 6927 12211 6979
rect 12267 6927 12319 6979
rect 1760 6878 1812 6885
rect 1868 6878 1920 6885
rect 1976 6878 2028 6885
rect 2084 6878 2136 6885
rect 2192 6878 2244 6885
rect 2300 6878 2352 6885
rect 2408 6878 2460 6885
rect 2516 6878 2568 6885
rect 2624 6878 2676 6885
rect 2732 6878 2784 6885
rect 2840 6878 2892 6885
rect 2948 6878 3000 6885
rect 3056 6878 3108 6885
rect 3164 6878 3216 6885
rect 3272 6878 3324 6885
rect 3380 6878 3432 6885
rect 3488 6878 3540 6885
rect 3596 6878 3648 6885
rect 3704 6878 3756 6885
rect 4130 6878 4182 6885
rect 4238 6878 4290 6885
rect 4346 6878 4398 6885
rect 4454 6878 4506 6885
rect 4562 6878 4614 6885
rect 4670 6878 4722 6885
rect 4778 6878 4830 6885
rect 4886 6878 4938 6885
rect 4994 6878 5046 6885
rect 5102 6878 5154 6885
rect 5210 6878 5262 6885
rect 5318 6878 5370 6885
rect 5426 6878 5478 6885
rect 5534 6878 5586 6885
rect 5642 6878 5694 6885
rect 5750 6878 5802 6885
rect 5858 6878 5910 6885
rect 5966 6878 6018 6885
rect 6074 6878 6126 6885
rect 6836 6878 6888 6885
rect 6944 6878 6996 6885
rect 7052 6878 7104 6885
rect 7160 6878 7212 6885
rect 7268 6878 7320 6885
rect 7376 6878 7428 6885
rect 7484 6878 7536 6885
rect 7592 6878 7644 6885
rect 7700 6878 7752 6885
rect 7808 6878 7860 6885
rect 7916 6878 7968 6885
rect 8024 6878 8076 6885
rect 8132 6878 8184 6885
rect 8240 6878 8292 6885
rect 8348 6878 8400 6885
rect 8456 6878 8508 6885
rect 8564 6878 8616 6885
rect 8672 6878 8724 6885
rect 8780 6878 8832 6885
rect 9206 6878 9258 6885
rect 9314 6878 9366 6885
rect 9422 6878 9474 6885
rect 9530 6878 9582 6885
rect 9638 6878 9690 6885
rect 9746 6878 9798 6885
rect 9854 6878 9906 6885
rect 9962 6878 10014 6885
rect 10070 6878 10122 6885
rect 10178 6878 10230 6885
rect 10286 6878 10338 6885
rect 10394 6878 10446 6885
rect 10502 6878 10554 6885
rect 10610 6878 10662 6885
rect 10718 6878 10770 6885
rect 10826 6878 10878 6885
rect 10934 6878 10986 6885
rect 11042 6878 11094 6885
rect 11150 6878 11202 6885
rect 643 6819 695 6871
rect 751 6819 803 6871
rect 859 6819 911 6871
rect 643 6711 695 6763
rect 751 6711 803 6763
rect 859 6711 911 6763
rect 1760 6833 1812 6878
rect 1868 6833 1920 6878
rect 1976 6833 2028 6878
rect 2084 6833 2136 6878
rect 2192 6833 2244 6878
rect 2300 6833 2352 6878
rect 2408 6833 2460 6878
rect 2516 6833 2568 6878
rect 2624 6833 2676 6878
rect 2732 6833 2784 6878
rect 2840 6833 2892 6878
rect 2948 6833 3000 6878
rect 3056 6833 3108 6878
rect 3164 6833 3216 6878
rect 3272 6833 3324 6878
rect 3380 6833 3432 6878
rect 3488 6833 3540 6878
rect 3596 6833 3648 6878
rect 3704 6833 3756 6878
rect 4130 6833 4182 6878
rect 4238 6833 4290 6878
rect 4346 6833 4398 6878
rect 4454 6833 4506 6878
rect 4562 6833 4614 6878
rect 4670 6833 4722 6878
rect 4778 6833 4830 6878
rect 4886 6833 4938 6878
rect 4994 6833 5046 6878
rect 5102 6833 5154 6878
rect 5210 6833 5262 6878
rect 5318 6833 5370 6878
rect 5426 6833 5478 6878
rect 5534 6833 5586 6878
rect 5642 6833 5694 6878
rect 5750 6833 5802 6878
rect 5858 6833 5910 6878
rect 5966 6833 6018 6878
rect 6074 6833 6126 6878
rect 6836 6833 6888 6878
rect 6944 6833 6996 6878
rect 7052 6833 7104 6878
rect 7160 6833 7212 6878
rect 7268 6833 7320 6878
rect 7376 6833 7428 6878
rect 7484 6833 7536 6878
rect 7592 6833 7644 6878
rect 7700 6833 7752 6878
rect 7808 6833 7860 6878
rect 7916 6833 7968 6878
rect 8024 6833 8076 6878
rect 8132 6833 8184 6878
rect 8240 6833 8292 6878
rect 8348 6833 8400 6878
rect 8456 6833 8508 6878
rect 8564 6833 8616 6878
rect 8672 6833 8724 6878
rect 8780 6833 8832 6878
rect 9206 6833 9258 6878
rect 9314 6833 9366 6878
rect 9422 6833 9474 6878
rect 9530 6833 9582 6878
rect 9638 6833 9690 6878
rect 9746 6833 9798 6878
rect 9854 6833 9906 6878
rect 9962 6833 10014 6878
rect 10070 6833 10122 6878
rect 10178 6833 10230 6878
rect 10286 6833 10338 6878
rect 10394 6833 10446 6878
rect 10502 6833 10554 6878
rect 10610 6833 10662 6878
rect 10718 6833 10770 6878
rect 10826 6833 10878 6878
rect 10934 6833 10986 6878
rect 11042 6833 11094 6878
rect 11150 6833 11202 6878
rect 1760 6732 1812 6777
rect 1868 6732 1920 6777
rect 1976 6732 2028 6777
rect 2084 6732 2136 6777
rect 2192 6732 2244 6777
rect 2300 6732 2352 6777
rect 2408 6732 2460 6777
rect 2516 6732 2568 6777
rect 2624 6732 2676 6777
rect 2732 6732 2784 6777
rect 2840 6732 2892 6777
rect 2948 6732 3000 6777
rect 3056 6732 3108 6777
rect 3164 6732 3216 6777
rect 3272 6732 3324 6777
rect 3380 6732 3432 6777
rect 3488 6732 3540 6777
rect 3596 6732 3648 6777
rect 3704 6732 3756 6777
rect 4130 6732 4182 6777
rect 4238 6732 4290 6777
rect 4346 6732 4398 6777
rect 4454 6732 4506 6777
rect 4562 6732 4614 6777
rect 4670 6732 4722 6777
rect 4778 6732 4830 6777
rect 4886 6732 4938 6777
rect 4994 6732 5046 6777
rect 5102 6732 5154 6777
rect 5210 6732 5262 6777
rect 5318 6732 5370 6777
rect 5426 6732 5478 6777
rect 5534 6732 5586 6777
rect 5642 6732 5694 6777
rect 5750 6732 5802 6777
rect 5858 6732 5910 6777
rect 5966 6732 6018 6777
rect 6074 6732 6126 6777
rect 6836 6732 6888 6777
rect 6944 6732 6996 6777
rect 7052 6732 7104 6777
rect 7160 6732 7212 6777
rect 7268 6732 7320 6777
rect 7376 6732 7428 6777
rect 7484 6732 7536 6777
rect 7592 6732 7644 6777
rect 7700 6732 7752 6777
rect 7808 6732 7860 6777
rect 7916 6732 7968 6777
rect 8024 6732 8076 6777
rect 8132 6732 8184 6777
rect 8240 6732 8292 6777
rect 8348 6732 8400 6777
rect 8456 6732 8508 6777
rect 8564 6732 8616 6777
rect 8672 6732 8724 6777
rect 8780 6732 8832 6777
rect 9206 6732 9258 6777
rect 9314 6732 9366 6777
rect 9422 6732 9474 6777
rect 9530 6732 9582 6777
rect 9638 6732 9690 6777
rect 9746 6732 9798 6777
rect 9854 6732 9906 6777
rect 9962 6732 10014 6777
rect 10070 6732 10122 6777
rect 10178 6732 10230 6777
rect 10286 6732 10338 6777
rect 10394 6732 10446 6777
rect 10502 6732 10554 6777
rect 10610 6732 10662 6777
rect 10718 6732 10770 6777
rect 10826 6732 10878 6777
rect 10934 6732 10986 6777
rect 11042 6732 11094 6777
rect 11150 6732 11202 6777
rect 12051 6819 12103 6871
rect 12159 6819 12211 6871
rect 12267 6819 12319 6871
rect 1760 6725 1812 6732
rect 1868 6725 1920 6732
rect 1976 6725 2028 6732
rect 2084 6725 2136 6732
rect 2192 6725 2244 6732
rect 2300 6725 2352 6732
rect 2408 6725 2460 6732
rect 2516 6725 2568 6732
rect 2624 6725 2676 6732
rect 2732 6725 2784 6732
rect 2840 6725 2892 6732
rect 2948 6725 3000 6732
rect 3056 6725 3108 6732
rect 3164 6725 3216 6732
rect 3272 6725 3324 6732
rect 3380 6725 3432 6732
rect 3488 6725 3540 6732
rect 3596 6725 3648 6732
rect 3704 6725 3756 6732
rect 4130 6725 4182 6732
rect 4238 6725 4290 6732
rect 4346 6725 4398 6732
rect 4454 6725 4506 6732
rect 4562 6725 4614 6732
rect 4670 6725 4722 6732
rect 4778 6725 4830 6732
rect 4886 6725 4938 6732
rect 4994 6725 5046 6732
rect 5102 6725 5154 6732
rect 5210 6725 5262 6732
rect 5318 6725 5370 6732
rect 5426 6725 5478 6732
rect 5534 6725 5586 6732
rect 5642 6725 5694 6732
rect 5750 6725 5802 6732
rect 5858 6725 5910 6732
rect 5966 6725 6018 6732
rect 6074 6725 6126 6732
rect 6836 6725 6888 6732
rect 6944 6725 6996 6732
rect 7052 6725 7104 6732
rect 7160 6725 7212 6732
rect 7268 6725 7320 6732
rect 7376 6725 7428 6732
rect 7484 6725 7536 6732
rect 7592 6725 7644 6732
rect 7700 6725 7752 6732
rect 7808 6725 7860 6732
rect 7916 6725 7968 6732
rect 8024 6725 8076 6732
rect 8132 6725 8184 6732
rect 8240 6725 8292 6732
rect 8348 6725 8400 6732
rect 8456 6725 8508 6732
rect 8564 6725 8616 6732
rect 8672 6725 8724 6732
rect 8780 6725 8832 6732
rect 9206 6725 9258 6732
rect 9314 6725 9366 6732
rect 9422 6725 9474 6732
rect 9530 6725 9582 6732
rect 9638 6725 9690 6732
rect 9746 6725 9798 6732
rect 9854 6725 9906 6732
rect 9962 6725 10014 6732
rect 10070 6725 10122 6732
rect 10178 6725 10230 6732
rect 10286 6725 10338 6732
rect 10394 6725 10446 6732
rect 10502 6725 10554 6732
rect 10610 6725 10662 6732
rect 10718 6725 10770 6732
rect 10826 6725 10878 6732
rect 10934 6725 10986 6732
rect 11042 6725 11094 6732
rect 11150 6725 11202 6732
rect 643 6603 695 6655
rect 751 6603 803 6655
rect 859 6603 911 6655
rect 643 6495 695 6547
rect 751 6495 803 6547
rect 859 6495 911 6547
rect 643 6387 695 6439
rect 751 6387 803 6439
rect 859 6387 911 6439
rect 643 6279 695 6331
rect 751 6279 803 6331
rect 859 6279 911 6331
rect 643 6171 695 6223
rect 751 6171 803 6223
rect 859 6171 911 6223
rect 643 6063 695 6115
rect 751 6063 803 6115
rect 859 6063 911 6115
rect 643 5955 695 6007
rect 751 5955 803 6007
rect 859 5955 911 6007
rect 643 5847 695 5899
rect 751 5847 803 5899
rect 859 5847 911 5899
rect 643 5739 695 5791
rect 751 5739 803 5791
rect 859 5739 911 5791
rect 643 5631 695 5683
rect 751 5631 803 5683
rect 859 5631 911 5683
rect 643 5523 695 5575
rect 751 5523 803 5575
rect 859 5523 911 5575
rect 643 5415 695 5467
rect 751 5415 803 5467
rect 859 5415 911 5467
rect 643 5307 695 5359
rect 751 5307 803 5359
rect 859 5307 911 5359
rect 643 5199 695 5251
rect 751 5199 803 5251
rect 859 5199 911 5251
rect 643 5091 695 5143
rect 751 5091 803 5143
rect 859 5091 911 5143
rect 643 4983 695 5035
rect 751 4983 803 5035
rect 859 4983 911 5035
rect 643 4875 695 4927
rect 751 4875 803 4927
rect 859 4875 911 4927
rect 643 4767 695 4819
rect 751 4767 803 4819
rect 859 4767 911 4819
rect 643 4659 695 4711
rect 751 4659 803 4711
rect 859 4659 911 4711
rect 643 4551 695 4603
rect 751 4551 803 4603
rect 859 4551 911 4603
rect 643 4443 695 4495
rect 751 4443 803 4495
rect 859 4443 911 4495
rect 643 4335 695 4387
rect 751 4335 803 4387
rect 859 4335 911 4387
rect 643 4227 695 4279
rect 751 4227 803 4279
rect 859 4227 911 4279
rect 643 4119 695 4171
rect 751 4119 803 4171
rect 859 4119 911 4171
rect 643 4011 695 4063
rect 751 4011 803 4063
rect 859 4011 911 4063
rect 643 3903 695 3955
rect 751 3903 803 3955
rect 859 3903 911 3955
rect 643 3795 695 3847
rect 751 3795 803 3847
rect 859 3795 911 3847
rect 643 3687 695 3739
rect 751 3687 803 3739
rect 859 3687 911 3739
rect 643 3579 695 3631
rect 751 3579 803 3631
rect 859 3579 911 3631
rect 643 3471 695 3523
rect 751 3471 803 3523
rect 859 3471 911 3523
rect 643 3363 695 3415
rect 751 3363 803 3415
rect 859 3363 911 3415
rect 643 3255 695 3307
rect 751 3255 803 3307
rect 859 3255 911 3307
rect 643 3147 695 3199
rect 751 3147 803 3199
rect 859 3147 911 3199
rect 643 3039 695 3091
rect 751 3039 803 3091
rect 859 3039 911 3091
rect 643 2931 695 2983
rect 751 2931 803 2983
rect 859 2931 911 2983
rect 643 2823 695 2875
rect 751 2823 803 2875
rect 859 2823 911 2875
rect 643 2715 695 2767
rect 751 2715 803 2767
rect 859 2715 911 2767
rect 643 2607 695 2659
rect 751 2607 803 2659
rect 859 2607 911 2659
rect 643 2499 695 2551
rect 751 2499 803 2551
rect 859 2499 911 2551
rect 643 2391 695 2443
rect 751 2391 803 2443
rect 859 2391 911 2443
rect 643 2283 695 2335
rect 751 2283 803 2335
rect 859 2283 911 2335
rect 643 2175 695 2227
rect 751 2175 803 2227
rect 859 2175 911 2227
rect 643 2067 695 2119
rect 751 2067 803 2119
rect 859 2067 911 2119
rect 643 1959 695 2011
rect 751 1959 803 2011
rect 859 1959 911 2011
rect 643 1851 695 1903
rect 751 1851 803 1903
rect 859 1851 911 1903
rect 643 1743 695 1795
rect 751 1743 803 1795
rect 859 1743 911 1795
rect 643 1635 695 1687
rect 751 1635 803 1687
rect 859 1635 911 1687
rect 643 1527 695 1579
rect 751 1527 803 1579
rect 859 1527 911 1579
rect 643 1419 695 1471
rect 751 1419 803 1471
rect 859 1419 911 1471
rect 643 1311 695 1363
rect 751 1311 803 1363
rect 859 1311 911 1363
rect 643 1203 695 1255
rect 751 1203 803 1255
rect 859 1203 911 1255
rect 643 1095 695 1147
rect 751 1095 803 1147
rect 859 1095 911 1147
rect 643 987 695 1039
rect 751 987 803 1039
rect 859 987 911 1039
rect 1760 6332 1812 6335
rect 1868 6332 1920 6335
rect 1976 6332 2028 6335
rect 2084 6332 2136 6335
rect 2192 6332 2244 6335
rect 2300 6332 2352 6335
rect 2408 6332 2460 6335
rect 2516 6332 2568 6335
rect 2624 6332 2676 6335
rect 2732 6332 2784 6335
rect 2840 6332 2892 6335
rect 2948 6332 3000 6335
rect 3056 6332 3108 6335
rect 3164 6332 3216 6335
rect 3272 6332 3324 6335
rect 3380 6332 3432 6335
rect 3488 6332 3540 6335
rect 3596 6332 3648 6335
rect 3704 6332 3756 6335
rect 4130 6332 4182 6335
rect 4238 6332 4290 6335
rect 4346 6332 4398 6335
rect 4454 6332 4506 6335
rect 4562 6332 4614 6335
rect 4670 6332 4722 6335
rect 4778 6332 4830 6335
rect 4886 6332 4938 6335
rect 4994 6332 5046 6335
rect 5102 6332 5154 6335
rect 5210 6332 5262 6335
rect 5318 6332 5370 6335
rect 5426 6332 5478 6335
rect 5534 6332 5586 6335
rect 5642 6332 5694 6335
rect 5750 6332 5802 6335
rect 5858 6332 5910 6335
rect 5966 6332 6018 6335
rect 6074 6332 6126 6335
rect 6836 6332 6888 6335
rect 6944 6332 6996 6335
rect 7052 6332 7104 6335
rect 7160 6332 7212 6335
rect 7268 6332 7320 6335
rect 7376 6332 7428 6335
rect 7484 6332 7536 6335
rect 7592 6332 7644 6335
rect 7700 6332 7752 6335
rect 7808 6332 7860 6335
rect 7916 6332 7968 6335
rect 8024 6332 8076 6335
rect 8132 6332 8184 6335
rect 8240 6332 8292 6335
rect 8348 6332 8400 6335
rect 8456 6332 8508 6335
rect 8564 6332 8616 6335
rect 8672 6332 8724 6335
rect 8780 6332 8832 6335
rect 9206 6332 9258 6335
rect 9314 6332 9366 6335
rect 9422 6332 9474 6335
rect 9530 6332 9582 6335
rect 9638 6332 9690 6335
rect 9746 6332 9798 6335
rect 9854 6332 9906 6335
rect 9962 6332 10014 6335
rect 10070 6332 10122 6335
rect 10178 6332 10230 6335
rect 10286 6332 10338 6335
rect 10394 6332 10446 6335
rect 10502 6332 10554 6335
rect 10610 6332 10662 6335
rect 10718 6332 10770 6335
rect 10826 6332 10878 6335
rect 10934 6332 10986 6335
rect 11042 6332 11094 6335
rect 11150 6332 11202 6335
rect 1760 6286 1812 6332
rect 1868 6286 1920 6332
rect 1976 6286 2028 6332
rect 2084 6286 2136 6332
rect 2192 6286 2244 6332
rect 2300 6286 2352 6332
rect 2408 6286 2460 6332
rect 2516 6286 2568 6332
rect 2624 6286 2676 6332
rect 2732 6286 2784 6332
rect 2840 6286 2892 6332
rect 2948 6286 3000 6332
rect 3056 6286 3108 6332
rect 3164 6286 3216 6332
rect 3272 6286 3324 6332
rect 3380 6286 3432 6332
rect 3488 6286 3540 6332
rect 3596 6286 3648 6332
rect 3704 6286 3756 6332
rect 4130 6286 4182 6332
rect 4238 6286 4290 6332
rect 4346 6286 4398 6332
rect 4454 6286 4506 6332
rect 4562 6286 4614 6332
rect 4670 6286 4722 6332
rect 4778 6286 4830 6332
rect 4886 6286 4938 6332
rect 4994 6286 5046 6332
rect 5102 6286 5154 6332
rect 5210 6286 5262 6332
rect 5318 6286 5370 6332
rect 5426 6286 5478 6332
rect 5534 6286 5586 6332
rect 5642 6286 5694 6332
rect 5750 6286 5802 6332
rect 5858 6286 5910 6332
rect 5966 6286 6018 6332
rect 6074 6286 6126 6332
rect 6836 6286 6888 6332
rect 6944 6286 6996 6332
rect 7052 6286 7104 6332
rect 7160 6286 7212 6332
rect 7268 6286 7320 6332
rect 7376 6286 7428 6332
rect 7484 6286 7536 6332
rect 7592 6286 7644 6332
rect 7700 6286 7752 6332
rect 7808 6286 7860 6332
rect 7916 6286 7968 6332
rect 8024 6286 8076 6332
rect 8132 6286 8184 6332
rect 8240 6286 8292 6332
rect 8348 6286 8400 6332
rect 8456 6286 8508 6332
rect 8564 6286 8616 6332
rect 8672 6286 8724 6332
rect 8780 6286 8832 6332
rect 9206 6286 9258 6332
rect 9314 6286 9366 6332
rect 9422 6286 9474 6332
rect 9530 6286 9582 6332
rect 9638 6286 9690 6332
rect 9746 6286 9798 6332
rect 9854 6286 9906 6332
rect 9962 6286 10014 6332
rect 10070 6286 10122 6332
rect 10178 6286 10230 6332
rect 10286 6286 10338 6332
rect 10394 6286 10446 6332
rect 10502 6286 10554 6332
rect 10610 6286 10662 6332
rect 10718 6286 10770 6332
rect 10826 6286 10878 6332
rect 10934 6286 10986 6332
rect 11042 6286 11094 6332
rect 11150 6286 11202 6332
rect 1760 6283 1812 6286
rect 1868 6283 1920 6286
rect 1976 6283 2028 6286
rect 2084 6283 2136 6286
rect 2192 6283 2244 6286
rect 2300 6283 2352 6286
rect 2408 6283 2460 6286
rect 2516 6283 2568 6286
rect 2624 6283 2676 6286
rect 2732 6283 2784 6286
rect 2840 6283 2892 6286
rect 2948 6283 3000 6286
rect 3056 6283 3108 6286
rect 3164 6283 3216 6286
rect 3272 6283 3324 6286
rect 3380 6283 3432 6286
rect 3488 6283 3540 6286
rect 3596 6283 3648 6286
rect 3704 6283 3756 6286
rect 4130 6283 4182 6286
rect 4238 6283 4290 6286
rect 4346 6283 4398 6286
rect 4454 6283 4506 6286
rect 4562 6283 4614 6286
rect 4670 6283 4722 6286
rect 4778 6283 4830 6286
rect 4886 6283 4938 6286
rect 4994 6283 5046 6286
rect 5102 6283 5154 6286
rect 5210 6283 5262 6286
rect 5318 6283 5370 6286
rect 5426 6283 5478 6286
rect 5534 6283 5586 6286
rect 5642 6283 5694 6286
rect 5750 6283 5802 6286
rect 5858 6283 5910 6286
rect 5966 6283 6018 6286
rect 6074 6283 6126 6286
rect 6836 6283 6888 6286
rect 6944 6283 6996 6286
rect 7052 6283 7104 6286
rect 7160 6283 7212 6286
rect 7268 6283 7320 6286
rect 7376 6283 7428 6286
rect 7484 6283 7536 6286
rect 7592 6283 7644 6286
rect 7700 6283 7752 6286
rect 7808 6283 7860 6286
rect 7916 6283 7968 6286
rect 8024 6283 8076 6286
rect 8132 6283 8184 6286
rect 8240 6283 8292 6286
rect 8348 6283 8400 6286
rect 8456 6283 8508 6286
rect 8564 6283 8616 6286
rect 8672 6283 8724 6286
rect 8780 6283 8832 6286
rect 9206 6283 9258 6286
rect 9314 6283 9366 6286
rect 9422 6283 9474 6286
rect 9530 6283 9582 6286
rect 9638 6283 9690 6286
rect 9746 6283 9798 6286
rect 9854 6283 9906 6286
rect 9962 6283 10014 6286
rect 10070 6283 10122 6286
rect 10178 6283 10230 6286
rect 10286 6283 10338 6286
rect 10394 6283 10446 6286
rect 10502 6283 10554 6286
rect 10610 6283 10662 6286
rect 10718 6283 10770 6286
rect 10826 6283 10878 6286
rect 10934 6283 10986 6286
rect 11042 6283 11094 6286
rect 11150 6283 11202 6286
rect 1233 6219 1285 6271
rect 1341 6219 1393 6271
rect 1233 6111 1256 6163
rect 1256 6111 1285 6163
rect 1341 6111 1393 6163
rect 1233 6003 1256 6055
rect 1256 6003 1285 6055
rect 1341 6003 1393 6055
rect 1233 5895 1256 5947
rect 1256 5895 1285 5947
rect 1341 5895 1393 5947
rect 1233 5787 1256 5839
rect 1256 5787 1285 5839
rect 1341 5787 1393 5839
rect 1233 5679 1256 5731
rect 1256 5679 1285 5731
rect 1341 5679 1393 5731
rect 1233 5571 1256 5623
rect 1256 5571 1285 5623
rect 1341 5571 1393 5623
rect 1233 5463 1256 5515
rect 1256 5463 1285 5515
rect 1341 5463 1393 5515
rect 1233 5355 1256 5407
rect 1256 5355 1285 5407
rect 1341 5355 1393 5407
rect 1233 5247 1256 5299
rect 1256 5247 1285 5299
rect 1341 5247 1393 5299
rect 1233 5139 1256 5191
rect 1256 5139 1285 5191
rect 1341 5139 1393 5191
rect 1233 5031 1256 5083
rect 1256 5031 1285 5083
rect 1341 5031 1393 5083
rect 1233 4923 1256 4975
rect 1256 4923 1285 4975
rect 1341 4923 1393 4975
rect 1233 4815 1256 4867
rect 1256 4815 1285 4867
rect 1341 4815 1393 4867
rect 1233 4707 1256 4759
rect 1256 4707 1285 4759
rect 1341 4707 1393 4759
rect 1233 4599 1256 4651
rect 1256 4599 1285 4651
rect 1341 4599 1393 4651
rect 1233 4491 1256 4543
rect 1256 4491 1285 4543
rect 1341 4491 1393 4543
rect 1233 4383 1256 4435
rect 1256 4383 1285 4435
rect 1341 4383 1393 4435
rect 1233 4275 1256 4327
rect 1256 4275 1285 4327
rect 1341 4275 1393 4327
rect 1233 4167 1256 4219
rect 1256 4167 1285 4219
rect 1341 4167 1393 4219
rect 1233 4059 1256 4111
rect 1256 4059 1285 4111
rect 1341 4059 1393 4111
rect 1233 3951 1256 4003
rect 1256 3951 1285 4003
rect 1341 3951 1393 4003
rect 1233 3843 1256 3895
rect 1256 3843 1285 3895
rect 1341 3843 1393 3895
rect 1233 3735 1256 3787
rect 1256 3735 1285 3787
rect 1341 3735 1393 3787
rect 1233 3627 1256 3679
rect 1256 3627 1285 3679
rect 1341 3627 1393 3679
rect 1233 3519 1256 3571
rect 1256 3519 1285 3571
rect 1341 3519 1393 3571
rect 1233 3411 1256 3463
rect 1256 3411 1285 3463
rect 1341 3411 1393 3463
rect 1233 3303 1256 3355
rect 1256 3303 1285 3355
rect 1341 3303 1393 3355
rect 1233 3195 1256 3247
rect 1256 3195 1285 3247
rect 1341 3195 1393 3247
rect 1233 3087 1256 3139
rect 1256 3087 1285 3139
rect 1341 3087 1393 3139
rect 1233 2979 1256 3031
rect 1256 2979 1285 3031
rect 1341 2979 1393 3031
rect 1233 2871 1256 2923
rect 1256 2871 1285 2923
rect 1341 2871 1393 2923
rect 1233 2763 1256 2815
rect 1256 2763 1285 2815
rect 1341 2763 1393 2815
rect 1233 2655 1256 2707
rect 1256 2655 1285 2707
rect 1341 2655 1393 2707
rect 1233 2547 1256 2599
rect 1256 2547 1285 2599
rect 1341 2547 1393 2599
rect 1233 2439 1256 2491
rect 1256 2439 1285 2491
rect 1341 2439 1393 2491
rect 1233 2331 1256 2383
rect 1256 2331 1285 2383
rect 1341 2331 1393 2383
rect 1233 2223 1256 2275
rect 1256 2223 1285 2275
rect 1341 2223 1393 2275
rect 1233 2115 1256 2167
rect 1256 2115 1285 2167
rect 1341 2115 1393 2167
rect 1233 2007 1256 2059
rect 1256 2007 1285 2059
rect 1341 2007 1393 2059
rect 1233 1899 1256 1951
rect 1256 1899 1285 1951
rect 1341 1899 1393 1951
rect 1233 1791 1256 1843
rect 1256 1791 1285 1843
rect 1341 1791 1393 1843
rect 1233 1683 1256 1735
rect 1256 1683 1285 1735
rect 1341 1683 1393 1735
rect 1233 1575 1256 1627
rect 1256 1575 1285 1627
rect 1341 1575 1393 1627
rect 11569 6219 11621 6271
rect 11677 6219 11729 6271
rect 1493 6088 1545 6091
rect 1601 6088 1653 6091
rect 3863 6088 3915 6091
rect 3971 6088 4023 6091
rect 6239 6088 6291 6091
rect 6347 6088 6399 6091
rect 6455 6088 6507 6091
rect 6563 6088 6615 6091
rect 6671 6088 6723 6091
rect 8939 6088 8991 6091
rect 9047 6088 9099 6091
rect 11309 6088 11361 6091
rect 11417 6088 11469 6091
rect 1493 6042 1494 6088
rect 1494 6042 1545 6088
rect 1601 6042 1653 6088
rect 3863 6042 3915 6088
rect 3971 6042 4023 6088
rect 6239 6042 6291 6088
rect 6347 6042 6399 6088
rect 6455 6042 6507 6088
rect 6563 6042 6615 6088
rect 6671 6042 6723 6088
rect 8939 6042 8991 6088
rect 9047 6042 9099 6088
rect 11309 6042 11361 6088
rect 11417 6042 11468 6088
rect 11468 6042 11469 6088
rect 1493 6039 1545 6042
rect 1601 6039 1653 6042
rect 3863 6039 3915 6042
rect 3971 6039 4023 6042
rect 6239 6039 6291 6042
rect 6347 6039 6399 6042
rect 6455 6039 6507 6042
rect 6563 6039 6615 6042
rect 6671 6039 6723 6042
rect 8939 6039 8991 6042
rect 9047 6039 9099 6042
rect 11309 6039 11361 6042
rect 11417 6039 11469 6042
rect 1760 5844 1812 5847
rect 1868 5844 1920 5847
rect 1976 5844 2028 5847
rect 2084 5844 2136 5847
rect 2192 5844 2244 5847
rect 2300 5844 2352 5847
rect 2408 5844 2460 5847
rect 2516 5844 2568 5847
rect 2624 5844 2676 5847
rect 2732 5844 2784 5847
rect 2840 5844 2892 5847
rect 2948 5844 3000 5847
rect 3056 5844 3108 5847
rect 3164 5844 3216 5847
rect 3272 5844 3324 5847
rect 3380 5844 3432 5847
rect 3488 5844 3540 5847
rect 3596 5844 3648 5847
rect 3704 5844 3756 5847
rect 4130 5844 4182 5847
rect 4238 5844 4290 5847
rect 4346 5844 4398 5847
rect 4454 5844 4506 5847
rect 4562 5844 4614 5847
rect 4670 5844 4722 5847
rect 4778 5844 4830 5847
rect 4886 5844 4938 5847
rect 4994 5844 5046 5847
rect 5102 5844 5154 5847
rect 5210 5844 5262 5847
rect 5318 5844 5370 5847
rect 5426 5844 5478 5847
rect 5534 5844 5586 5847
rect 5642 5844 5694 5847
rect 5750 5844 5802 5847
rect 5858 5844 5910 5847
rect 5966 5844 6018 5847
rect 6074 5844 6126 5847
rect 6836 5844 6888 5847
rect 6944 5844 6996 5847
rect 7052 5844 7104 5847
rect 7160 5844 7212 5847
rect 7268 5844 7320 5847
rect 7376 5844 7428 5847
rect 7484 5844 7536 5847
rect 7592 5844 7644 5847
rect 7700 5844 7752 5847
rect 7808 5844 7860 5847
rect 7916 5844 7968 5847
rect 8024 5844 8076 5847
rect 8132 5844 8184 5847
rect 8240 5844 8292 5847
rect 8348 5844 8400 5847
rect 8456 5844 8508 5847
rect 8564 5844 8616 5847
rect 8672 5844 8724 5847
rect 8780 5844 8832 5847
rect 9206 5844 9258 5847
rect 9314 5844 9366 5847
rect 9422 5844 9474 5847
rect 9530 5844 9582 5847
rect 9638 5844 9690 5847
rect 9746 5844 9798 5847
rect 9854 5844 9906 5847
rect 9962 5844 10014 5847
rect 10070 5844 10122 5847
rect 10178 5844 10230 5847
rect 10286 5844 10338 5847
rect 10394 5844 10446 5847
rect 10502 5844 10554 5847
rect 10610 5844 10662 5847
rect 10718 5844 10770 5847
rect 10826 5844 10878 5847
rect 10934 5844 10986 5847
rect 11042 5844 11094 5847
rect 11150 5844 11202 5847
rect 1760 5798 1812 5844
rect 1868 5798 1920 5844
rect 1976 5798 2028 5844
rect 2084 5798 2136 5844
rect 2192 5798 2244 5844
rect 2300 5798 2352 5844
rect 2408 5798 2460 5844
rect 2516 5798 2568 5844
rect 2624 5798 2676 5844
rect 2732 5798 2784 5844
rect 2840 5798 2892 5844
rect 2948 5798 3000 5844
rect 3056 5798 3108 5844
rect 3164 5798 3216 5844
rect 3272 5798 3324 5844
rect 3380 5798 3432 5844
rect 3488 5798 3540 5844
rect 3596 5798 3648 5844
rect 3704 5798 3756 5844
rect 4130 5798 4182 5844
rect 4238 5798 4290 5844
rect 4346 5798 4398 5844
rect 4454 5798 4506 5844
rect 4562 5798 4614 5844
rect 4670 5798 4722 5844
rect 4778 5798 4830 5844
rect 4886 5798 4938 5844
rect 4994 5798 5046 5844
rect 5102 5798 5154 5844
rect 5210 5798 5262 5844
rect 5318 5798 5370 5844
rect 5426 5798 5478 5844
rect 5534 5798 5586 5844
rect 5642 5798 5694 5844
rect 5750 5798 5802 5844
rect 5858 5798 5910 5844
rect 5966 5798 6018 5844
rect 6074 5798 6126 5844
rect 6836 5798 6888 5844
rect 6944 5798 6996 5844
rect 7052 5798 7104 5844
rect 7160 5798 7212 5844
rect 7268 5798 7320 5844
rect 7376 5798 7428 5844
rect 7484 5798 7536 5844
rect 7592 5798 7644 5844
rect 7700 5798 7752 5844
rect 7808 5798 7860 5844
rect 7916 5798 7968 5844
rect 8024 5798 8076 5844
rect 8132 5798 8184 5844
rect 8240 5798 8292 5844
rect 8348 5798 8400 5844
rect 8456 5798 8508 5844
rect 8564 5798 8616 5844
rect 8672 5798 8724 5844
rect 8780 5798 8832 5844
rect 9206 5798 9258 5844
rect 9314 5798 9366 5844
rect 9422 5798 9474 5844
rect 9530 5798 9582 5844
rect 9638 5798 9690 5844
rect 9746 5798 9798 5844
rect 9854 5798 9906 5844
rect 9962 5798 10014 5844
rect 10070 5798 10122 5844
rect 10178 5798 10230 5844
rect 10286 5798 10338 5844
rect 10394 5798 10446 5844
rect 10502 5798 10554 5844
rect 10610 5798 10662 5844
rect 10718 5798 10770 5844
rect 10826 5798 10878 5844
rect 10934 5798 10986 5844
rect 11042 5798 11094 5844
rect 11150 5798 11202 5844
rect 1760 5795 1812 5798
rect 1868 5795 1920 5798
rect 1976 5795 2028 5798
rect 2084 5795 2136 5798
rect 2192 5795 2244 5798
rect 2300 5795 2352 5798
rect 2408 5795 2460 5798
rect 2516 5795 2568 5798
rect 2624 5795 2676 5798
rect 2732 5795 2784 5798
rect 2840 5795 2892 5798
rect 2948 5795 3000 5798
rect 3056 5795 3108 5798
rect 3164 5795 3216 5798
rect 3272 5795 3324 5798
rect 3380 5795 3432 5798
rect 3488 5795 3540 5798
rect 3596 5795 3648 5798
rect 3704 5795 3756 5798
rect 4130 5795 4182 5798
rect 4238 5795 4290 5798
rect 4346 5795 4398 5798
rect 4454 5795 4506 5798
rect 4562 5795 4614 5798
rect 4670 5795 4722 5798
rect 4778 5795 4830 5798
rect 4886 5795 4938 5798
rect 4994 5795 5046 5798
rect 5102 5795 5154 5798
rect 5210 5795 5262 5798
rect 5318 5795 5370 5798
rect 5426 5795 5478 5798
rect 5534 5795 5586 5798
rect 5642 5795 5694 5798
rect 5750 5795 5802 5798
rect 5858 5795 5910 5798
rect 5966 5795 6018 5798
rect 6074 5795 6126 5798
rect 6836 5795 6888 5798
rect 6944 5795 6996 5798
rect 7052 5795 7104 5798
rect 7160 5795 7212 5798
rect 7268 5795 7320 5798
rect 7376 5795 7428 5798
rect 7484 5795 7536 5798
rect 7592 5795 7644 5798
rect 7700 5795 7752 5798
rect 7808 5795 7860 5798
rect 7916 5795 7968 5798
rect 8024 5795 8076 5798
rect 8132 5795 8184 5798
rect 8240 5795 8292 5798
rect 8348 5795 8400 5798
rect 8456 5795 8508 5798
rect 8564 5795 8616 5798
rect 8672 5795 8724 5798
rect 8780 5795 8832 5798
rect 9206 5795 9258 5798
rect 9314 5795 9366 5798
rect 9422 5795 9474 5798
rect 9530 5795 9582 5798
rect 9638 5795 9690 5798
rect 9746 5795 9798 5798
rect 9854 5795 9906 5798
rect 9962 5795 10014 5798
rect 10070 5795 10122 5798
rect 10178 5795 10230 5798
rect 10286 5795 10338 5798
rect 10394 5795 10446 5798
rect 10502 5795 10554 5798
rect 10610 5795 10662 5798
rect 10718 5795 10770 5798
rect 10826 5795 10878 5798
rect 10934 5795 10986 5798
rect 11042 5795 11094 5798
rect 11150 5795 11202 5798
rect 1493 5600 1545 5603
rect 1601 5600 1653 5603
rect 3863 5600 3915 5603
rect 3971 5600 4023 5603
rect 6239 5600 6291 5603
rect 6347 5600 6399 5603
rect 6455 5600 6507 5603
rect 6563 5600 6615 5603
rect 6671 5600 6723 5603
rect 8939 5600 8991 5603
rect 9047 5600 9099 5603
rect 11309 5600 11361 5603
rect 11417 5600 11469 5603
rect 1493 5554 1494 5600
rect 1494 5554 1545 5600
rect 1601 5554 1653 5600
rect 3863 5554 3915 5600
rect 3971 5554 4023 5600
rect 6239 5554 6291 5600
rect 6347 5554 6399 5600
rect 6455 5554 6507 5600
rect 6563 5554 6615 5600
rect 6671 5554 6723 5600
rect 8939 5554 8991 5600
rect 9047 5554 9099 5600
rect 11309 5554 11361 5600
rect 11417 5554 11468 5600
rect 11468 5554 11469 5600
rect 1493 5551 1545 5554
rect 1601 5551 1653 5554
rect 3863 5551 3915 5554
rect 3971 5551 4023 5554
rect 6239 5551 6291 5554
rect 6347 5551 6399 5554
rect 6455 5551 6507 5554
rect 6563 5551 6615 5554
rect 6671 5551 6723 5554
rect 8939 5551 8991 5554
rect 9047 5551 9099 5554
rect 11309 5551 11361 5554
rect 11417 5551 11469 5554
rect 1760 5356 1812 5359
rect 1868 5356 1920 5359
rect 1976 5356 2028 5359
rect 2084 5356 2136 5359
rect 2192 5356 2244 5359
rect 2300 5356 2352 5359
rect 2408 5356 2460 5359
rect 2516 5356 2568 5359
rect 2624 5356 2676 5359
rect 2732 5356 2784 5359
rect 2840 5356 2892 5359
rect 2948 5356 3000 5359
rect 3056 5356 3108 5359
rect 3164 5356 3216 5359
rect 3272 5356 3324 5359
rect 3380 5356 3432 5359
rect 3488 5356 3540 5359
rect 3596 5356 3648 5359
rect 3704 5356 3756 5359
rect 4130 5356 4182 5359
rect 4238 5356 4290 5359
rect 4346 5356 4398 5359
rect 4454 5356 4506 5359
rect 4562 5356 4614 5359
rect 4670 5356 4722 5359
rect 4778 5356 4830 5359
rect 4886 5356 4938 5359
rect 4994 5356 5046 5359
rect 5102 5356 5154 5359
rect 5210 5356 5262 5359
rect 5318 5356 5370 5359
rect 5426 5356 5478 5359
rect 5534 5356 5586 5359
rect 5642 5356 5694 5359
rect 5750 5356 5802 5359
rect 5858 5356 5910 5359
rect 5966 5356 6018 5359
rect 6074 5356 6126 5359
rect 6836 5356 6888 5359
rect 6944 5356 6996 5359
rect 7052 5356 7104 5359
rect 7160 5356 7212 5359
rect 7268 5356 7320 5359
rect 7376 5356 7428 5359
rect 7484 5356 7536 5359
rect 7592 5356 7644 5359
rect 7700 5356 7752 5359
rect 7808 5356 7860 5359
rect 7916 5356 7968 5359
rect 8024 5356 8076 5359
rect 8132 5356 8184 5359
rect 8240 5356 8292 5359
rect 8348 5356 8400 5359
rect 8456 5356 8508 5359
rect 8564 5356 8616 5359
rect 8672 5356 8724 5359
rect 8780 5356 8832 5359
rect 9206 5356 9258 5359
rect 9314 5356 9366 5359
rect 9422 5356 9474 5359
rect 9530 5356 9582 5359
rect 9638 5356 9690 5359
rect 9746 5356 9798 5359
rect 9854 5356 9906 5359
rect 9962 5356 10014 5359
rect 10070 5356 10122 5359
rect 10178 5356 10230 5359
rect 10286 5356 10338 5359
rect 10394 5356 10446 5359
rect 10502 5356 10554 5359
rect 10610 5356 10662 5359
rect 10718 5356 10770 5359
rect 10826 5356 10878 5359
rect 10934 5356 10986 5359
rect 11042 5356 11094 5359
rect 11150 5356 11202 5359
rect 1760 5310 1812 5356
rect 1868 5310 1920 5356
rect 1976 5310 2028 5356
rect 2084 5310 2136 5356
rect 2192 5310 2244 5356
rect 2300 5310 2352 5356
rect 2408 5310 2460 5356
rect 2516 5310 2568 5356
rect 2624 5310 2676 5356
rect 2732 5310 2784 5356
rect 2840 5310 2892 5356
rect 2948 5310 3000 5356
rect 3056 5310 3108 5356
rect 3164 5310 3216 5356
rect 3272 5310 3324 5356
rect 3380 5310 3432 5356
rect 3488 5310 3540 5356
rect 3596 5310 3648 5356
rect 3704 5310 3756 5356
rect 4130 5310 4182 5356
rect 4238 5310 4290 5356
rect 4346 5310 4398 5356
rect 4454 5310 4506 5356
rect 4562 5310 4614 5356
rect 4670 5310 4722 5356
rect 4778 5310 4830 5356
rect 4886 5310 4938 5356
rect 4994 5310 5046 5356
rect 5102 5310 5154 5356
rect 5210 5310 5262 5356
rect 5318 5310 5370 5356
rect 5426 5310 5478 5356
rect 5534 5310 5586 5356
rect 5642 5310 5694 5356
rect 5750 5310 5802 5356
rect 5858 5310 5910 5356
rect 5966 5310 6018 5356
rect 6074 5310 6126 5356
rect 6836 5310 6888 5356
rect 6944 5310 6996 5356
rect 7052 5310 7104 5356
rect 7160 5310 7212 5356
rect 7268 5310 7320 5356
rect 7376 5310 7428 5356
rect 7484 5310 7536 5356
rect 7592 5310 7644 5356
rect 7700 5310 7752 5356
rect 7808 5310 7860 5356
rect 7916 5310 7968 5356
rect 8024 5310 8076 5356
rect 8132 5310 8184 5356
rect 8240 5310 8292 5356
rect 8348 5310 8400 5356
rect 8456 5310 8508 5356
rect 8564 5310 8616 5356
rect 8672 5310 8724 5356
rect 8780 5310 8832 5356
rect 9206 5310 9258 5356
rect 9314 5310 9366 5356
rect 9422 5310 9474 5356
rect 9530 5310 9582 5356
rect 9638 5310 9690 5356
rect 9746 5310 9798 5356
rect 9854 5310 9906 5356
rect 9962 5310 10014 5356
rect 10070 5310 10122 5356
rect 10178 5310 10230 5356
rect 10286 5310 10338 5356
rect 10394 5310 10446 5356
rect 10502 5310 10554 5356
rect 10610 5310 10662 5356
rect 10718 5310 10770 5356
rect 10826 5310 10878 5356
rect 10934 5310 10986 5356
rect 11042 5310 11094 5356
rect 11150 5310 11202 5356
rect 1760 5307 1812 5310
rect 1868 5307 1920 5310
rect 1976 5307 2028 5310
rect 2084 5307 2136 5310
rect 2192 5307 2244 5310
rect 2300 5307 2352 5310
rect 2408 5307 2460 5310
rect 2516 5307 2568 5310
rect 2624 5307 2676 5310
rect 2732 5307 2784 5310
rect 2840 5307 2892 5310
rect 2948 5307 3000 5310
rect 3056 5307 3108 5310
rect 3164 5307 3216 5310
rect 3272 5307 3324 5310
rect 3380 5307 3432 5310
rect 3488 5307 3540 5310
rect 3596 5307 3648 5310
rect 3704 5307 3756 5310
rect 4130 5307 4182 5310
rect 4238 5307 4290 5310
rect 4346 5307 4398 5310
rect 4454 5307 4506 5310
rect 4562 5307 4614 5310
rect 4670 5307 4722 5310
rect 4778 5307 4830 5310
rect 4886 5307 4938 5310
rect 4994 5307 5046 5310
rect 5102 5307 5154 5310
rect 5210 5307 5262 5310
rect 5318 5307 5370 5310
rect 5426 5307 5478 5310
rect 5534 5307 5586 5310
rect 5642 5307 5694 5310
rect 5750 5307 5802 5310
rect 5858 5307 5910 5310
rect 5966 5307 6018 5310
rect 6074 5307 6126 5310
rect 6836 5307 6888 5310
rect 6944 5307 6996 5310
rect 7052 5307 7104 5310
rect 7160 5307 7212 5310
rect 7268 5307 7320 5310
rect 7376 5307 7428 5310
rect 7484 5307 7536 5310
rect 7592 5307 7644 5310
rect 7700 5307 7752 5310
rect 7808 5307 7860 5310
rect 7916 5307 7968 5310
rect 8024 5307 8076 5310
rect 8132 5307 8184 5310
rect 8240 5307 8292 5310
rect 8348 5307 8400 5310
rect 8456 5307 8508 5310
rect 8564 5307 8616 5310
rect 8672 5307 8724 5310
rect 8780 5307 8832 5310
rect 9206 5307 9258 5310
rect 9314 5307 9366 5310
rect 9422 5307 9474 5310
rect 9530 5307 9582 5310
rect 9638 5307 9690 5310
rect 9746 5307 9798 5310
rect 9854 5307 9906 5310
rect 9962 5307 10014 5310
rect 10070 5307 10122 5310
rect 10178 5307 10230 5310
rect 10286 5307 10338 5310
rect 10394 5307 10446 5310
rect 10502 5307 10554 5310
rect 10610 5307 10662 5310
rect 10718 5307 10770 5310
rect 10826 5307 10878 5310
rect 10934 5307 10986 5310
rect 11042 5307 11094 5310
rect 11150 5307 11202 5310
rect 1493 5112 1545 5115
rect 1601 5112 1653 5115
rect 3863 5112 3915 5115
rect 3971 5112 4023 5115
rect 6239 5112 6291 5115
rect 6347 5112 6399 5115
rect 6455 5112 6507 5115
rect 6563 5112 6615 5115
rect 6671 5112 6723 5115
rect 8939 5112 8991 5115
rect 9047 5112 9099 5115
rect 11309 5112 11361 5115
rect 11417 5112 11469 5115
rect 1493 5066 1494 5112
rect 1494 5066 1545 5112
rect 1601 5066 1653 5112
rect 3863 5066 3915 5112
rect 3971 5066 4023 5112
rect 6239 5066 6291 5112
rect 6347 5066 6399 5112
rect 6455 5066 6507 5112
rect 6563 5066 6615 5112
rect 6671 5066 6723 5112
rect 8939 5066 8991 5112
rect 9047 5066 9099 5112
rect 11309 5066 11361 5112
rect 11417 5066 11468 5112
rect 11468 5066 11469 5112
rect 1493 5063 1545 5066
rect 1601 5063 1653 5066
rect 3863 5063 3915 5066
rect 3971 5063 4023 5066
rect 6239 5063 6291 5066
rect 6347 5063 6399 5066
rect 6455 5063 6507 5066
rect 6563 5063 6615 5066
rect 6671 5063 6723 5066
rect 8939 5063 8991 5066
rect 9047 5063 9099 5066
rect 11309 5063 11361 5066
rect 11417 5063 11469 5066
rect 1760 4868 1812 4871
rect 1868 4868 1920 4871
rect 1976 4868 2028 4871
rect 2084 4868 2136 4871
rect 2192 4868 2244 4871
rect 2300 4868 2352 4871
rect 2408 4868 2460 4871
rect 2516 4868 2568 4871
rect 2624 4868 2676 4871
rect 2732 4868 2784 4871
rect 2840 4868 2892 4871
rect 2948 4868 3000 4871
rect 3056 4868 3108 4871
rect 3164 4868 3216 4871
rect 3272 4868 3324 4871
rect 3380 4868 3432 4871
rect 3488 4868 3540 4871
rect 3596 4868 3648 4871
rect 3704 4868 3756 4871
rect 4130 4868 4182 4871
rect 4238 4868 4290 4871
rect 4346 4868 4398 4871
rect 4454 4868 4506 4871
rect 4562 4868 4614 4871
rect 4670 4868 4722 4871
rect 4778 4868 4830 4871
rect 4886 4868 4938 4871
rect 4994 4868 5046 4871
rect 5102 4868 5154 4871
rect 5210 4868 5262 4871
rect 5318 4868 5370 4871
rect 5426 4868 5478 4871
rect 5534 4868 5586 4871
rect 5642 4868 5694 4871
rect 5750 4868 5802 4871
rect 5858 4868 5910 4871
rect 5966 4868 6018 4871
rect 6074 4868 6126 4871
rect 6836 4868 6888 4871
rect 6944 4868 6996 4871
rect 7052 4868 7104 4871
rect 7160 4868 7212 4871
rect 7268 4868 7320 4871
rect 7376 4868 7428 4871
rect 7484 4868 7536 4871
rect 7592 4868 7644 4871
rect 7700 4868 7752 4871
rect 7808 4868 7860 4871
rect 7916 4868 7968 4871
rect 8024 4868 8076 4871
rect 8132 4868 8184 4871
rect 8240 4868 8292 4871
rect 8348 4868 8400 4871
rect 8456 4868 8508 4871
rect 8564 4868 8616 4871
rect 8672 4868 8724 4871
rect 8780 4868 8832 4871
rect 9206 4868 9258 4871
rect 9314 4868 9366 4871
rect 9422 4868 9474 4871
rect 9530 4868 9582 4871
rect 9638 4868 9690 4871
rect 9746 4868 9798 4871
rect 9854 4868 9906 4871
rect 9962 4868 10014 4871
rect 10070 4868 10122 4871
rect 10178 4868 10230 4871
rect 10286 4868 10338 4871
rect 10394 4868 10446 4871
rect 10502 4868 10554 4871
rect 10610 4868 10662 4871
rect 10718 4868 10770 4871
rect 10826 4868 10878 4871
rect 10934 4868 10986 4871
rect 11042 4868 11094 4871
rect 11150 4868 11202 4871
rect 1760 4822 1812 4868
rect 1868 4822 1920 4868
rect 1976 4822 2028 4868
rect 2084 4822 2136 4868
rect 2192 4822 2244 4868
rect 2300 4822 2352 4868
rect 2408 4822 2460 4868
rect 2516 4822 2568 4868
rect 2624 4822 2676 4868
rect 2732 4822 2784 4868
rect 2840 4822 2892 4868
rect 2948 4822 3000 4868
rect 3056 4822 3108 4868
rect 3164 4822 3216 4868
rect 3272 4822 3324 4868
rect 3380 4822 3432 4868
rect 3488 4822 3540 4868
rect 3596 4822 3648 4868
rect 3704 4822 3756 4868
rect 4130 4822 4182 4868
rect 4238 4822 4290 4868
rect 4346 4822 4398 4868
rect 4454 4822 4506 4868
rect 4562 4822 4614 4868
rect 4670 4822 4722 4868
rect 4778 4822 4830 4868
rect 4886 4822 4938 4868
rect 4994 4822 5046 4868
rect 5102 4822 5154 4868
rect 5210 4822 5262 4868
rect 5318 4822 5370 4868
rect 5426 4822 5478 4868
rect 5534 4822 5586 4868
rect 5642 4822 5694 4868
rect 5750 4822 5802 4868
rect 5858 4822 5910 4868
rect 5966 4822 6018 4868
rect 6074 4822 6126 4868
rect 6836 4822 6888 4868
rect 6944 4822 6996 4868
rect 7052 4822 7104 4868
rect 7160 4822 7212 4868
rect 7268 4822 7320 4868
rect 7376 4822 7428 4868
rect 7484 4822 7536 4868
rect 7592 4822 7644 4868
rect 7700 4822 7752 4868
rect 7808 4822 7860 4868
rect 7916 4822 7968 4868
rect 8024 4822 8076 4868
rect 8132 4822 8184 4868
rect 8240 4822 8292 4868
rect 8348 4822 8400 4868
rect 8456 4822 8508 4868
rect 8564 4822 8616 4868
rect 8672 4822 8724 4868
rect 8780 4822 8832 4868
rect 9206 4822 9258 4868
rect 9314 4822 9366 4868
rect 9422 4822 9474 4868
rect 9530 4822 9582 4868
rect 9638 4822 9690 4868
rect 9746 4822 9798 4868
rect 9854 4822 9906 4868
rect 9962 4822 10014 4868
rect 10070 4822 10122 4868
rect 10178 4822 10230 4868
rect 10286 4822 10338 4868
rect 10394 4822 10446 4868
rect 10502 4822 10554 4868
rect 10610 4822 10662 4868
rect 10718 4822 10770 4868
rect 10826 4822 10878 4868
rect 10934 4822 10986 4868
rect 11042 4822 11094 4868
rect 11150 4822 11202 4868
rect 1760 4819 1812 4822
rect 1868 4819 1920 4822
rect 1976 4819 2028 4822
rect 2084 4819 2136 4822
rect 2192 4819 2244 4822
rect 2300 4819 2352 4822
rect 2408 4819 2460 4822
rect 2516 4819 2568 4822
rect 2624 4819 2676 4822
rect 2732 4819 2784 4822
rect 2840 4819 2892 4822
rect 2948 4819 3000 4822
rect 3056 4819 3108 4822
rect 3164 4819 3216 4822
rect 3272 4819 3324 4822
rect 3380 4819 3432 4822
rect 3488 4819 3540 4822
rect 3596 4819 3648 4822
rect 3704 4819 3756 4822
rect 4130 4819 4182 4822
rect 4238 4819 4290 4822
rect 4346 4819 4398 4822
rect 4454 4819 4506 4822
rect 4562 4819 4614 4822
rect 4670 4819 4722 4822
rect 4778 4819 4830 4822
rect 4886 4819 4938 4822
rect 4994 4819 5046 4822
rect 5102 4819 5154 4822
rect 5210 4819 5262 4822
rect 5318 4819 5370 4822
rect 5426 4819 5478 4822
rect 5534 4819 5586 4822
rect 5642 4819 5694 4822
rect 5750 4819 5802 4822
rect 5858 4819 5910 4822
rect 5966 4819 6018 4822
rect 6074 4819 6126 4822
rect 6836 4819 6888 4822
rect 6944 4819 6996 4822
rect 7052 4819 7104 4822
rect 7160 4819 7212 4822
rect 7268 4819 7320 4822
rect 7376 4819 7428 4822
rect 7484 4819 7536 4822
rect 7592 4819 7644 4822
rect 7700 4819 7752 4822
rect 7808 4819 7860 4822
rect 7916 4819 7968 4822
rect 8024 4819 8076 4822
rect 8132 4819 8184 4822
rect 8240 4819 8292 4822
rect 8348 4819 8400 4822
rect 8456 4819 8508 4822
rect 8564 4819 8616 4822
rect 8672 4819 8724 4822
rect 8780 4819 8832 4822
rect 9206 4819 9258 4822
rect 9314 4819 9366 4822
rect 9422 4819 9474 4822
rect 9530 4819 9582 4822
rect 9638 4819 9690 4822
rect 9746 4819 9798 4822
rect 9854 4819 9906 4822
rect 9962 4819 10014 4822
rect 10070 4819 10122 4822
rect 10178 4819 10230 4822
rect 10286 4819 10338 4822
rect 10394 4819 10446 4822
rect 10502 4819 10554 4822
rect 10610 4819 10662 4822
rect 10718 4819 10770 4822
rect 10826 4819 10878 4822
rect 10934 4819 10986 4822
rect 11042 4819 11094 4822
rect 11150 4819 11202 4822
rect 1493 4624 1545 4627
rect 1601 4624 1653 4627
rect 3863 4624 3915 4627
rect 3971 4624 4023 4627
rect 6239 4624 6291 4627
rect 6347 4624 6399 4627
rect 6455 4624 6507 4627
rect 6563 4624 6615 4627
rect 6671 4624 6723 4627
rect 8939 4624 8991 4627
rect 9047 4624 9099 4627
rect 11309 4624 11361 4627
rect 11417 4624 11469 4627
rect 1493 4578 1494 4624
rect 1494 4578 1545 4624
rect 1601 4578 1653 4624
rect 3863 4578 3915 4624
rect 3971 4578 4023 4624
rect 6239 4578 6291 4624
rect 6347 4578 6399 4624
rect 6455 4578 6507 4624
rect 6563 4578 6615 4624
rect 6671 4578 6723 4624
rect 8939 4578 8991 4624
rect 9047 4578 9099 4624
rect 11309 4578 11361 4624
rect 11417 4578 11468 4624
rect 11468 4578 11469 4624
rect 1493 4575 1545 4578
rect 1601 4575 1653 4578
rect 3863 4575 3915 4578
rect 3971 4575 4023 4578
rect 6239 4575 6291 4578
rect 6347 4575 6399 4578
rect 6455 4575 6507 4578
rect 6563 4575 6615 4578
rect 6671 4575 6723 4578
rect 8939 4575 8991 4578
rect 9047 4575 9099 4578
rect 11309 4575 11361 4578
rect 11417 4575 11469 4578
rect 1760 4380 1812 4383
rect 1868 4380 1920 4383
rect 1976 4380 2028 4383
rect 2084 4380 2136 4383
rect 2192 4380 2244 4383
rect 2300 4380 2352 4383
rect 2408 4380 2460 4383
rect 2516 4380 2568 4383
rect 2624 4380 2676 4383
rect 2732 4380 2784 4383
rect 2840 4380 2892 4383
rect 2948 4380 3000 4383
rect 3056 4380 3108 4383
rect 3164 4380 3216 4383
rect 3272 4380 3324 4383
rect 3380 4380 3432 4383
rect 3488 4380 3540 4383
rect 3596 4380 3648 4383
rect 3704 4380 3756 4383
rect 4130 4380 4182 4383
rect 4238 4380 4290 4383
rect 4346 4380 4398 4383
rect 4454 4380 4506 4383
rect 4562 4380 4614 4383
rect 4670 4380 4722 4383
rect 4778 4380 4830 4383
rect 4886 4380 4938 4383
rect 4994 4380 5046 4383
rect 5102 4380 5154 4383
rect 5210 4380 5262 4383
rect 5318 4380 5370 4383
rect 5426 4380 5478 4383
rect 5534 4380 5586 4383
rect 5642 4380 5694 4383
rect 5750 4380 5802 4383
rect 5858 4380 5910 4383
rect 5966 4380 6018 4383
rect 6074 4380 6126 4383
rect 6836 4380 6888 4383
rect 6944 4380 6996 4383
rect 7052 4380 7104 4383
rect 7160 4380 7212 4383
rect 7268 4380 7320 4383
rect 7376 4380 7428 4383
rect 7484 4380 7536 4383
rect 7592 4380 7644 4383
rect 7700 4380 7752 4383
rect 7808 4380 7860 4383
rect 7916 4380 7968 4383
rect 8024 4380 8076 4383
rect 8132 4380 8184 4383
rect 8240 4380 8292 4383
rect 8348 4380 8400 4383
rect 8456 4380 8508 4383
rect 8564 4380 8616 4383
rect 8672 4380 8724 4383
rect 8780 4380 8832 4383
rect 9206 4380 9258 4383
rect 9314 4380 9366 4383
rect 9422 4380 9474 4383
rect 9530 4380 9582 4383
rect 9638 4380 9690 4383
rect 9746 4380 9798 4383
rect 9854 4380 9906 4383
rect 9962 4380 10014 4383
rect 10070 4380 10122 4383
rect 10178 4380 10230 4383
rect 10286 4380 10338 4383
rect 10394 4380 10446 4383
rect 10502 4380 10554 4383
rect 10610 4380 10662 4383
rect 10718 4380 10770 4383
rect 10826 4380 10878 4383
rect 10934 4380 10986 4383
rect 11042 4380 11094 4383
rect 11150 4380 11202 4383
rect 1760 4334 1812 4380
rect 1868 4334 1920 4380
rect 1976 4334 2028 4380
rect 2084 4334 2136 4380
rect 2192 4334 2244 4380
rect 2300 4334 2352 4380
rect 2408 4334 2460 4380
rect 2516 4334 2568 4380
rect 2624 4334 2676 4380
rect 2732 4334 2784 4380
rect 2840 4334 2892 4380
rect 2948 4334 3000 4380
rect 3056 4334 3108 4380
rect 3164 4334 3216 4380
rect 3272 4334 3324 4380
rect 3380 4334 3432 4380
rect 3488 4334 3540 4380
rect 3596 4334 3648 4380
rect 3704 4334 3756 4380
rect 4130 4334 4182 4380
rect 4238 4334 4290 4380
rect 4346 4334 4398 4380
rect 4454 4334 4506 4380
rect 4562 4334 4614 4380
rect 4670 4334 4722 4380
rect 4778 4334 4830 4380
rect 4886 4334 4938 4380
rect 4994 4334 5046 4380
rect 5102 4334 5154 4380
rect 5210 4334 5262 4380
rect 5318 4334 5370 4380
rect 5426 4334 5478 4380
rect 5534 4334 5586 4380
rect 5642 4334 5694 4380
rect 5750 4334 5802 4380
rect 5858 4334 5910 4380
rect 5966 4334 6018 4380
rect 6074 4334 6126 4380
rect 6836 4334 6888 4380
rect 6944 4334 6996 4380
rect 7052 4334 7104 4380
rect 7160 4334 7212 4380
rect 7268 4334 7320 4380
rect 7376 4334 7428 4380
rect 7484 4334 7536 4380
rect 7592 4334 7644 4380
rect 7700 4334 7752 4380
rect 7808 4334 7860 4380
rect 7916 4334 7968 4380
rect 8024 4334 8076 4380
rect 8132 4334 8184 4380
rect 8240 4334 8292 4380
rect 8348 4334 8400 4380
rect 8456 4334 8508 4380
rect 8564 4334 8616 4380
rect 8672 4334 8724 4380
rect 8780 4334 8832 4380
rect 9206 4334 9258 4380
rect 9314 4334 9366 4380
rect 9422 4334 9474 4380
rect 9530 4334 9582 4380
rect 9638 4334 9690 4380
rect 9746 4334 9798 4380
rect 9854 4334 9906 4380
rect 9962 4334 10014 4380
rect 10070 4334 10122 4380
rect 10178 4334 10230 4380
rect 10286 4334 10338 4380
rect 10394 4334 10446 4380
rect 10502 4334 10554 4380
rect 10610 4334 10662 4380
rect 10718 4334 10770 4380
rect 10826 4334 10878 4380
rect 10934 4334 10986 4380
rect 11042 4334 11094 4380
rect 11150 4334 11202 4380
rect 1760 4331 1812 4334
rect 1868 4331 1920 4334
rect 1976 4331 2028 4334
rect 2084 4331 2136 4334
rect 2192 4331 2244 4334
rect 2300 4331 2352 4334
rect 2408 4331 2460 4334
rect 2516 4331 2568 4334
rect 2624 4331 2676 4334
rect 2732 4331 2784 4334
rect 2840 4331 2892 4334
rect 2948 4331 3000 4334
rect 3056 4331 3108 4334
rect 3164 4331 3216 4334
rect 3272 4331 3324 4334
rect 3380 4331 3432 4334
rect 3488 4331 3540 4334
rect 3596 4331 3648 4334
rect 3704 4331 3756 4334
rect 4130 4331 4182 4334
rect 4238 4331 4290 4334
rect 4346 4331 4398 4334
rect 4454 4331 4506 4334
rect 4562 4331 4614 4334
rect 4670 4331 4722 4334
rect 4778 4331 4830 4334
rect 4886 4331 4938 4334
rect 4994 4331 5046 4334
rect 5102 4331 5154 4334
rect 5210 4331 5262 4334
rect 5318 4331 5370 4334
rect 5426 4331 5478 4334
rect 5534 4331 5586 4334
rect 5642 4331 5694 4334
rect 5750 4331 5802 4334
rect 5858 4331 5910 4334
rect 5966 4331 6018 4334
rect 6074 4331 6126 4334
rect 6836 4331 6888 4334
rect 6944 4331 6996 4334
rect 7052 4331 7104 4334
rect 7160 4331 7212 4334
rect 7268 4331 7320 4334
rect 7376 4331 7428 4334
rect 7484 4331 7536 4334
rect 7592 4331 7644 4334
rect 7700 4331 7752 4334
rect 7808 4331 7860 4334
rect 7916 4331 7968 4334
rect 8024 4331 8076 4334
rect 8132 4331 8184 4334
rect 8240 4331 8292 4334
rect 8348 4331 8400 4334
rect 8456 4331 8508 4334
rect 8564 4331 8616 4334
rect 8672 4331 8724 4334
rect 8780 4331 8832 4334
rect 9206 4331 9258 4334
rect 9314 4331 9366 4334
rect 9422 4331 9474 4334
rect 9530 4331 9582 4334
rect 9638 4331 9690 4334
rect 9746 4331 9798 4334
rect 9854 4331 9906 4334
rect 9962 4331 10014 4334
rect 10070 4331 10122 4334
rect 10178 4331 10230 4334
rect 10286 4331 10338 4334
rect 10394 4331 10446 4334
rect 10502 4331 10554 4334
rect 10610 4331 10662 4334
rect 10718 4331 10770 4334
rect 10826 4331 10878 4334
rect 10934 4331 10986 4334
rect 11042 4331 11094 4334
rect 11150 4331 11202 4334
rect 1493 4136 1545 4139
rect 1601 4136 1653 4139
rect 3863 4136 3915 4139
rect 3971 4136 4023 4139
rect 6239 4136 6291 4139
rect 6347 4136 6399 4139
rect 6455 4136 6507 4139
rect 6563 4136 6615 4139
rect 6671 4136 6723 4139
rect 8939 4136 8991 4139
rect 9047 4136 9099 4139
rect 11309 4136 11361 4139
rect 11417 4136 11469 4139
rect 1493 4090 1494 4136
rect 1494 4090 1545 4136
rect 1601 4090 1653 4136
rect 3863 4090 3915 4136
rect 3971 4090 4023 4136
rect 6239 4090 6291 4136
rect 6347 4090 6399 4136
rect 6455 4090 6507 4136
rect 6563 4090 6615 4136
rect 6671 4090 6723 4136
rect 8939 4090 8991 4136
rect 9047 4090 9099 4136
rect 11309 4090 11361 4136
rect 11417 4090 11468 4136
rect 11468 4090 11469 4136
rect 1493 4087 1545 4090
rect 1601 4087 1653 4090
rect 3863 4087 3915 4090
rect 3971 4087 4023 4090
rect 6239 4087 6291 4090
rect 6347 4087 6399 4090
rect 6455 4087 6507 4090
rect 6563 4087 6615 4090
rect 6671 4087 6723 4090
rect 8939 4087 8991 4090
rect 9047 4087 9099 4090
rect 11309 4087 11361 4090
rect 11417 4087 11469 4090
rect 1760 3892 1812 3895
rect 1868 3892 1920 3895
rect 1976 3892 2028 3895
rect 2084 3892 2136 3895
rect 2192 3892 2244 3895
rect 2300 3892 2352 3895
rect 2408 3892 2460 3895
rect 2516 3892 2568 3895
rect 2624 3892 2676 3895
rect 2732 3892 2784 3895
rect 2840 3892 2892 3895
rect 2948 3892 3000 3895
rect 3056 3892 3108 3895
rect 3164 3892 3216 3895
rect 3272 3892 3324 3895
rect 3380 3892 3432 3895
rect 3488 3892 3540 3895
rect 3596 3892 3648 3895
rect 3704 3892 3756 3895
rect 4130 3892 4182 3895
rect 4238 3892 4290 3895
rect 4346 3892 4398 3895
rect 4454 3892 4506 3895
rect 4562 3892 4614 3895
rect 4670 3892 4722 3895
rect 4778 3892 4830 3895
rect 4886 3892 4938 3895
rect 4994 3892 5046 3895
rect 5102 3892 5154 3895
rect 5210 3892 5262 3895
rect 5318 3892 5370 3895
rect 5426 3892 5478 3895
rect 5534 3892 5586 3895
rect 5642 3892 5694 3895
rect 5750 3892 5802 3895
rect 5858 3892 5910 3895
rect 5966 3892 6018 3895
rect 6074 3892 6126 3895
rect 6836 3892 6888 3895
rect 6944 3892 6996 3895
rect 7052 3892 7104 3895
rect 7160 3892 7212 3895
rect 7268 3892 7320 3895
rect 7376 3892 7428 3895
rect 7484 3892 7536 3895
rect 7592 3892 7644 3895
rect 7700 3892 7752 3895
rect 7808 3892 7860 3895
rect 7916 3892 7968 3895
rect 8024 3892 8076 3895
rect 8132 3892 8184 3895
rect 8240 3892 8292 3895
rect 8348 3892 8400 3895
rect 8456 3892 8508 3895
rect 8564 3892 8616 3895
rect 8672 3892 8724 3895
rect 8780 3892 8832 3895
rect 9206 3892 9258 3895
rect 9314 3892 9366 3895
rect 9422 3892 9474 3895
rect 9530 3892 9582 3895
rect 9638 3892 9690 3895
rect 9746 3892 9798 3895
rect 9854 3892 9906 3895
rect 9962 3892 10014 3895
rect 10070 3892 10122 3895
rect 10178 3892 10230 3895
rect 10286 3892 10338 3895
rect 10394 3892 10446 3895
rect 10502 3892 10554 3895
rect 10610 3892 10662 3895
rect 10718 3892 10770 3895
rect 10826 3892 10878 3895
rect 10934 3892 10986 3895
rect 11042 3892 11094 3895
rect 11150 3892 11202 3895
rect 1760 3846 1812 3892
rect 1868 3846 1920 3892
rect 1976 3846 2028 3892
rect 2084 3846 2136 3892
rect 2192 3846 2244 3892
rect 2300 3846 2352 3892
rect 2408 3846 2460 3892
rect 2516 3846 2568 3892
rect 2624 3846 2676 3892
rect 2732 3846 2784 3892
rect 2840 3846 2892 3892
rect 2948 3846 3000 3892
rect 3056 3846 3108 3892
rect 3164 3846 3216 3892
rect 3272 3846 3324 3892
rect 3380 3846 3432 3892
rect 3488 3846 3540 3892
rect 3596 3846 3648 3892
rect 3704 3846 3756 3892
rect 4130 3846 4182 3892
rect 4238 3846 4290 3892
rect 4346 3846 4398 3892
rect 4454 3846 4506 3892
rect 4562 3846 4614 3892
rect 4670 3846 4722 3892
rect 4778 3846 4830 3892
rect 4886 3846 4938 3892
rect 4994 3846 5046 3892
rect 5102 3846 5154 3892
rect 5210 3846 5262 3892
rect 5318 3846 5370 3892
rect 5426 3846 5478 3892
rect 5534 3846 5586 3892
rect 5642 3846 5694 3892
rect 5750 3846 5802 3892
rect 5858 3846 5910 3892
rect 5966 3846 6018 3892
rect 6074 3846 6126 3892
rect 6836 3846 6888 3892
rect 6944 3846 6996 3892
rect 7052 3846 7104 3892
rect 7160 3846 7212 3892
rect 7268 3846 7320 3892
rect 7376 3846 7428 3892
rect 7484 3846 7536 3892
rect 7592 3846 7644 3892
rect 7700 3846 7752 3892
rect 7808 3846 7860 3892
rect 7916 3846 7968 3892
rect 8024 3846 8076 3892
rect 8132 3846 8184 3892
rect 8240 3846 8292 3892
rect 8348 3846 8400 3892
rect 8456 3846 8508 3892
rect 8564 3846 8616 3892
rect 8672 3846 8724 3892
rect 8780 3846 8832 3892
rect 9206 3846 9258 3892
rect 9314 3846 9366 3892
rect 9422 3846 9474 3892
rect 9530 3846 9582 3892
rect 9638 3846 9690 3892
rect 9746 3846 9798 3892
rect 9854 3846 9906 3892
rect 9962 3846 10014 3892
rect 10070 3846 10122 3892
rect 10178 3846 10230 3892
rect 10286 3846 10338 3892
rect 10394 3846 10446 3892
rect 10502 3846 10554 3892
rect 10610 3846 10662 3892
rect 10718 3846 10770 3892
rect 10826 3846 10878 3892
rect 10934 3846 10986 3892
rect 11042 3846 11094 3892
rect 11150 3846 11202 3892
rect 1760 3843 1812 3846
rect 1868 3843 1920 3846
rect 1976 3843 2028 3846
rect 2084 3843 2136 3846
rect 2192 3843 2244 3846
rect 2300 3843 2352 3846
rect 2408 3843 2460 3846
rect 2516 3843 2568 3846
rect 2624 3843 2676 3846
rect 2732 3843 2784 3846
rect 2840 3843 2892 3846
rect 2948 3843 3000 3846
rect 3056 3843 3108 3846
rect 3164 3843 3216 3846
rect 3272 3843 3324 3846
rect 3380 3843 3432 3846
rect 3488 3843 3540 3846
rect 3596 3843 3648 3846
rect 3704 3843 3756 3846
rect 4130 3843 4182 3846
rect 4238 3843 4290 3846
rect 4346 3843 4398 3846
rect 4454 3843 4506 3846
rect 4562 3843 4614 3846
rect 4670 3843 4722 3846
rect 4778 3843 4830 3846
rect 4886 3843 4938 3846
rect 4994 3843 5046 3846
rect 5102 3843 5154 3846
rect 5210 3843 5262 3846
rect 5318 3843 5370 3846
rect 5426 3843 5478 3846
rect 5534 3843 5586 3846
rect 5642 3843 5694 3846
rect 5750 3843 5802 3846
rect 5858 3843 5910 3846
rect 5966 3843 6018 3846
rect 6074 3843 6126 3846
rect 6836 3843 6888 3846
rect 6944 3843 6996 3846
rect 7052 3843 7104 3846
rect 7160 3843 7212 3846
rect 7268 3843 7320 3846
rect 7376 3843 7428 3846
rect 7484 3843 7536 3846
rect 7592 3843 7644 3846
rect 7700 3843 7752 3846
rect 7808 3843 7860 3846
rect 7916 3843 7968 3846
rect 8024 3843 8076 3846
rect 8132 3843 8184 3846
rect 8240 3843 8292 3846
rect 8348 3843 8400 3846
rect 8456 3843 8508 3846
rect 8564 3843 8616 3846
rect 8672 3843 8724 3846
rect 8780 3843 8832 3846
rect 9206 3843 9258 3846
rect 9314 3843 9366 3846
rect 9422 3843 9474 3846
rect 9530 3843 9582 3846
rect 9638 3843 9690 3846
rect 9746 3843 9798 3846
rect 9854 3843 9906 3846
rect 9962 3843 10014 3846
rect 10070 3843 10122 3846
rect 10178 3843 10230 3846
rect 10286 3843 10338 3846
rect 10394 3843 10446 3846
rect 10502 3843 10554 3846
rect 10610 3843 10662 3846
rect 10718 3843 10770 3846
rect 10826 3843 10878 3846
rect 10934 3843 10986 3846
rect 11042 3843 11094 3846
rect 11150 3843 11202 3846
rect 1493 3648 1545 3651
rect 1601 3648 1653 3651
rect 3863 3648 3915 3651
rect 3971 3648 4023 3651
rect 6239 3648 6291 3651
rect 6347 3648 6399 3651
rect 6455 3648 6507 3651
rect 6563 3648 6615 3651
rect 6671 3648 6723 3651
rect 8939 3648 8991 3651
rect 9047 3648 9099 3651
rect 11309 3648 11361 3651
rect 11417 3648 11469 3651
rect 1493 3602 1494 3648
rect 1494 3602 1545 3648
rect 1601 3602 1653 3648
rect 3863 3602 3915 3648
rect 3971 3602 4023 3648
rect 6239 3602 6291 3648
rect 6347 3602 6399 3648
rect 6455 3602 6507 3648
rect 6563 3602 6615 3648
rect 6671 3602 6723 3648
rect 8939 3602 8991 3648
rect 9047 3602 9099 3648
rect 11309 3602 11361 3648
rect 11417 3602 11468 3648
rect 11468 3602 11469 3648
rect 1493 3599 1545 3602
rect 1601 3599 1653 3602
rect 3863 3599 3915 3602
rect 3971 3599 4023 3602
rect 6239 3599 6291 3602
rect 6347 3599 6399 3602
rect 6455 3599 6507 3602
rect 6563 3599 6615 3602
rect 6671 3599 6723 3602
rect 8939 3599 8991 3602
rect 9047 3599 9099 3602
rect 11309 3599 11361 3602
rect 11417 3599 11469 3602
rect 1760 3404 1812 3407
rect 1868 3404 1920 3407
rect 1976 3404 2028 3407
rect 2084 3404 2136 3407
rect 2192 3404 2244 3407
rect 2300 3404 2352 3407
rect 2408 3404 2460 3407
rect 2516 3404 2568 3407
rect 2624 3404 2676 3407
rect 2732 3404 2784 3407
rect 2840 3404 2892 3407
rect 2948 3404 3000 3407
rect 3056 3404 3108 3407
rect 3164 3404 3216 3407
rect 3272 3404 3324 3407
rect 3380 3404 3432 3407
rect 3488 3404 3540 3407
rect 3596 3404 3648 3407
rect 3704 3404 3756 3407
rect 4130 3404 4182 3407
rect 4238 3404 4290 3407
rect 4346 3404 4398 3407
rect 4454 3404 4506 3407
rect 4562 3404 4614 3407
rect 4670 3404 4722 3407
rect 4778 3404 4830 3407
rect 4886 3404 4938 3407
rect 4994 3404 5046 3407
rect 5102 3404 5154 3407
rect 5210 3404 5262 3407
rect 5318 3404 5370 3407
rect 5426 3404 5478 3407
rect 5534 3404 5586 3407
rect 5642 3404 5694 3407
rect 5750 3404 5802 3407
rect 5858 3404 5910 3407
rect 5966 3404 6018 3407
rect 6074 3404 6126 3407
rect 6836 3404 6888 3407
rect 6944 3404 6996 3407
rect 7052 3404 7104 3407
rect 7160 3404 7212 3407
rect 7268 3404 7320 3407
rect 7376 3404 7428 3407
rect 7484 3404 7536 3407
rect 7592 3404 7644 3407
rect 7700 3404 7752 3407
rect 7808 3404 7860 3407
rect 7916 3404 7968 3407
rect 8024 3404 8076 3407
rect 8132 3404 8184 3407
rect 8240 3404 8292 3407
rect 8348 3404 8400 3407
rect 8456 3404 8508 3407
rect 8564 3404 8616 3407
rect 8672 3404 8724 3407
rect 8780 3404 8832 3407
rect 9206 3404 9258 3407
rect 9314 3404 9366 3407
rect 9422 3404 9474 3407
rect 9530 3404 9582 3407
rect 9638 3404 9690 3407
rect 9746 3404 9798 3407
rect 9854 3404 9906 3407
rect 9962 3404 10014 3407
rect 10070 3404 10122 3407
rect 10178 3404 10230 3407
rect 10286 3404 10338 3407
rect 10394 3404 10446 3407
rect 10502 3404 10554 3407
rect 10610 3404 10662 3407
rect 10718 3404 10770 3407
rect 10826 3404 10878 3407
rect 10934 3404 10986 3407
rect 11042 3404 11094 3407
rect 11150 3404 11202 3407
rect 1760 3358 1812 3404
rect 1868 3358 1920 3404
rect 1976 3358 2028 3404
rect 2084 3358 2136 3404
rect 2192 3358 2244 3404
rect 2300 3358 2352 3404
rect 2408 3358 2460 3404
rect 2516 3358 2568 3404
rect 2624 3358 2676 3404
rect 2732 3358 2784 3404
rect 2840 3358 2892 3404
rect 2948 3358 3000 3404
rect 3056 3358 3108 3404
rect 3164 3358 3216 3404
rect 3272 3358 3324 3404
rect 3380 3358 3432 3404
rect 3488 3358 3540 3404
rect 3596 3358 3648 3404
rect 3704 3358 3756 3404
rect 4130 3358 4182 3404
rect 4238 3358 4290 3404
rect 4346 3358 4398 3404
rect 4454 3358 4506 3404
rect 4562 3358 4614 3404
rect 4670 3358 4722 3404
rect 4778 3358 4830 3404
rect 4886 3358 4938 3404
rect 4994 3358 5046 3404
rect 5102 3358 5154 3404
rect 5210 3358 5262 3404
rect 5318 3358 5370 3404
rect 5426 3358 5478 3404
rect 5534 3358 5586 3404
rect 5642 3358 5694 3404
rect 5750 3358 5802 3404
rect 5858 3358 5910 3404
rect 5966 3358 6018 3404
rect 6074 3358 6126 3404
rect 6836 3358 6888 3404
rect 6944 3358 6996 3404
rect 7052 3358 7104 3404
rect 7160 3358 7212 3404
rect 7268 3358 7320 3404
rect 7376 3358 7428 3404
rect 7484 3358 7536 3404
rect 7592 3358 7644 3404
rect 7700 3358 7752 3404
rect 7808 3358 7860 3404
rect 7916 3358 7968 3404
rect 8024 3358 8076 3404
rect 8132 3358 8184 3404
rect 8240 3358 8292 3404
rect 8348 3358 8400 3404
rect 8456 3358 8508 3404
rect 8564 3358 8616 3404
rect 8672 3358 8724 3404
rect 8780 3358 8832 3404
rect 9206 3358 9258 3404
rect 9314 3358 9366 3404
rect 9422 3358 9474 3404
rect 9530 3358 9582 3404
rect 9638 3358 9690 3404
rect 9746 3358 9798 3404
rect 9854 3358 9906 3404
rect 9962 3358 10014 3404
rect 10070 3358 10122 3404
rect 10178 3358 10230 3404
rect 10286 3358 10338 3404
rect 10394 3358 10446 3404
rect 10502 3358 10554 3404
rect 10610 3358 10662 3404
rect 10718 3358 10770 3404
rect 10826 3358 10878 3404
rect 10934 3358 10986 3404
rect 11042 3358 11094 3404
rect 11150 3358 11202 3404
rect 1760 3355 1812 3358
rect 1868 3355 1920 3358
rect 1976 3355 2028 3358
rect 2084 3355 2136 3358
rect 2192 3355 2244 3358
rect 2300 3355 2352 3358
rect 2408 3355 2460 3358
rect 2516 3355 2568 3358
rect 2624 3355 2676 3358
rect 2732 3355 2784 3358
rect 2840 3355 2892 3358
rect 2948 3355 3000 3358
rect 3056 3355 3108 3358
rect 3164 3355 3216 3358
rect 3272 3355 3324 3358
rect 3380 3355 3432 3358
rect 3488 3355 3540 3358
rect 3596 3355 3648 3358
rect 3704 3355 3756 3358
rect 4130 3355 4182 3358
rect 4238 3355 4290 3358
rect 4346 3355 4398 3358
rect 4454 3355 4506 3358
rect 4562 3355 4614 3358
rect 4670 3355 4722 3358
rect 4778 3355 4830 3358
rect 4886 3355 4938 3358
rect 4994 3355 5046 3358
rect 5102 3355 5154 3358
rect 5210 3355 5262 3358
rect 5318 3355 5370 3358
rect 5426 3355 5478 3358
rect 5534 3355 5586 3358
rect 5642 3355 5694 3358
rect 5750 3355 5802 3358
rect 5858 3355 5910 3358
rect 5966 3355 6018 3358
rect 6074 3355 6126 3358
rect 6836 3355 6888 3358
rect 6944 3355 6996 3358
rect 7052 3355 7104 3358
rect 7160 3355 7212 3358
rect 7268 3355 7320 3358
rect 7376 3355 7428 3358
rect 7484 3355 7536 3358
rect 7592 3355 7644 3358
rect 7700 3355 7752 3358
rect 7808 3355 7860 3358
rect 7916 3355 7968 3358
rect 8024 3355 8076 3358
rect 8132 3355 8184 3358
rect 8240 3355 8292 3358
rect 8348 3355 8400 3358
rect 8456 3355 8508 3358
rect 8564 3355 8616 3358
rect 8672 3355 8724 3358
rect 8780 3355 8832 3358
rect 9206 3355 9258 3358
rect 9314 3355 9366 3358
rect 9422 3355 9474 3358
rect 9530 3355 9582 3358
rect 9638 3355 9690 3358
rect 9746 3355 9798 3358
rect 9854 3355 9906 3358
rect 9962 3355 10014 3358
rect 10070 3355 10122 3358
rect 10178 3355 10230 3358
rect 10286 3355 10338 3358
rect 10394 3355 10446 3358
rect 10502 3355 10554 3358
rect 10610 3355 10662 3358
rect 10718 3355 10770 3358
rect 10826 3355 10878 3358
rect 10934 3355 10986 3358
rect 11042 3355 11094 3358
rect 11150 3355 11202 3358
rect 1493 3160 1545 3163
rect 1601 3160 1653 3163
rect 3863 3160 3915 3163
rect 3971 3160 4023 3163
rect 6239 3160 6291 3163
rect 6347 3160 6399 3163
rect 6455 3160 6507 3163
rect 6563 3160 6615 3163
rect 6671 3160 6723 3163
rect 8939 3160 8991 3163
rect 9047 3160 9099 3163
rect 11309 3160 11361 3163
rect 11417 3160 11469 3163
rect 1493 3114 1494 3160
rect 1494 3114 1545 3160
rect 1601 3114 1653 3160
rect 3863 3114 3915 3160
rect 3971 3114 4023 3160
rect 6239 3114 6291 3160
rect 6347 3114 6399 3160
rect 6455 3114 6507 3160
rect 6563 3114 6615 3160
rect 6671 3114 6723 3160
rect 8939 3114 8991 3160
rect 9047 3114 9099 3160
rect 11309 3114 11361 3160
rect 11417 3114 11468 3160
rect 11468 3114 11469 3160
rect 1493 3111 1545 3114
rect 1601 3111 1653 3114
rect 3863 3111 3915 3114
rect 3971 3111 4023 3114
rect 6239 3111 6291 3114
rect 6347 3111 6399 3114
rect 6455 3111 6507 3114
rect 6563 3111 6615 3114
rect 6671 3111 6723 3114
rect 8939 3111 8991 3114
rect 9047 3111 9099 3114
rect 11309 3111 11361 3114
rect 11417 3111 11469 3114
rect 1760 2916 1812 2919
rect 1868 2916 1920 2919
rect 1976 2916 2028 2919
rect 2084 2916 2136 2919
rect 2192 2916 2244 2919
rect 2300 2916 2352 2919
rect 2408 2916 2460 2919
rect 2516 2916 2568 2919
rect 2624 2916 2676 2919
rect 2732 2916 2784 2919
rect 2840 2916 2892 2919
rect 2948 2916 3000 2919
rect 3056 2916 3108 2919
rect 3164 2916 3216 2919
rect 3272 2916 3324 2919
rect 3380 2916 3432 2919
rect 3488 2916 3540 2919
rect 3596 2916 3648 2919
rect 3704 2916 3756 2919
rect 4130 2916 4182 2919
rect 4238 2916 4290 2919
rect 4346 2916 4398 2919
rect 4454 2916 4506 2919
rect 4562 2916 4614 2919
rect 4670 2916 4722 2919
rect 4778 2916 4830 2919
rect 4886 2916 4938 2919
rect 4994 2916 5046 2919
rect 5102 2916 5154 2919
rect 5210 2916 5262 2919
rect 5318 2916 5370 2919
rect 5426 2916 5478 2919
rect 5534 2916 5586 2919
rect 5642 2916 5694 2919
rect 5750 2916 5802 2919
rect 5858 2916 5910 2919
rect 5966 2916 6018 2919
rect 6074 2916 6126 2919
rect 6836 2916 6888 2919
rect 6944 2916 6996 2919
rect 7052 2916 7104 2919
rect 7160 2916 7212 2919
rect 7268 2916 7320 2919
rect 7376 2916 7428 2919
rect 7484 2916 7536 2919
rect 7592 2916 7644 2919
rect 7700 2916 7752 2919
rect 7808 2916 7860 2919
rect 7916 2916 7968 2919
rect 8024 2916 8076 2919
rect 8132 2916 8184 2919
rect 8240 2916 8292 2919
rect 8348 2916 8400 2919
rect 8456 2916 8508 2919
rect 8564 2916 8616 2919
rect 8672 2916 8724 2919
rect 8780 2916 8832 2919
rect 9206 2916 9258 2919
rect 9314 2916 9366 2919
rect 9422 2916 9474 2919
rect 9530 2916 9582 2919
rect 9638 2916 9690 2919
rect 9746 2916 9798 2919
rect 9854 2916 9906 2919
rect 9962 2916 10014 2919
rect 10070 2916 10122 2919
rect 10178 2916 10230 2919
rect 10286 2916 10338 2919
rect 10394 2916 10446 2919
rect 10502 2916 10554 2919
rect 10610 2916 10662 2919
rect 10718 2916 10770 2919
rect 10826 2916 10878 2919
rect 10934 2916 10986 2919
rect 11042 2916 11094 2919
rect 11150 2916 11202 2919
rect 1760 2870 1812 2916
rect 1868 2870 1920 2916
rect 1976 2870 2028 2916
rect 2084 2870 2136 2916
rect 2192 2870 2244 2916
rect 2300 2870 2352 2916
rect 2408 2870 2460 2916
rect 2516 2870 2568 2916
rect 2624 2870 2676 2916
rect 2732 2870 2784 2916
rect 2840 2870 2892 2916
rect 2948 2870 3000 2916
rect 3056 2870 3108 2916
rect 3164 2870 3216 2916
rect 3272 2870 3324 2916
rect 3380 2870 3432 2916
rect 3488 2870 3540 2916
rect 3596 2870 3648 2916
rect 3704 2870 3756 2916
rect 4130 2870 4182 2916
rect 4238 2870 4290 2916
rect 4346 2870 4398 2916
rect 4454 2870 4506 2916
rect 4562 2870 4614 2916
rect 4670 2870 4722 2916
rect 4778 2870 4830 2916
rect 4886 2870 4938 2916
rect 4994 2870 5046 2916
rect 5102 2870 5154 2916
rect 5210 2870 5262 2916
rect 5318 2870 5370 2916
rect 5426 2870 5478 2916
rect 5534 2870 5586 2916
rect 5642 2870 5694 2916
rect 5750 2870 5802 2916
rect 5858 2870 5910 2916
rect 5966 2870 6018 2916
rect 6074 2870 6126 2916
rect 6836 2870 6888 2916
rect 6944 2870 6996 2916
rect 7052 2870 7104 2916
rect 7160 2870 7212 2916
rect 7268 2870 7320 2916
rect 7376 2870 7428 2916
rect 7484 2870 7536 2916
rect 7592 2870 7644 2916
rect 7700 2870 7752 2916
rect 7808 2870 7860 2916
rect 7916 2870 7968 2916
rect 8024 2870 8076 2916
rect 8132 2870 8184 2916
rect 8240 2870 8292 2916
rect 8348 2870 8400 2916
rect 8456 2870 8508 2916
rect 8564 2870 8616 2916
rect 8672 2870 8724 2916
rect 8780 2870 8832 2916
rect 9206 2870 9258 2916
rect 9314 2870 9366 2916
rect 9422 2870 9474 2916
rect 9530 2870 9582 2916
rect 9638 2870 9690 2916
rect 9746 2870 9798 2916
rect 9854 2870 9906 2916
rect 9962 2870 10014 2916
rect 10070 2870 10122 2916
rect 10178 2870 10230 2916
rect 10286 2870 10338 2916
rect 10394 2870 10446 2916
rect 10502 2870 10554 2916
rect 10610 2870 10662 2916
rect 10718 2870 10770 2916
rect 10826 2870 10878 2916
rect 10934 2870 10986 2916
rect 11042 2870 11094 2916
rect 11150 2870 11202 2916
rect 1760 2867 1812 2870
rect 1868 2867 1920 2870
rect 1976 2867 2028 2870
rect 2084 2867 2136 2870
rect 2192 2867 2244 2870
rect 2300 2867 2352 2870
rect 2408 2867 2460 2870
rect 2516 2867 2568 2870
rect 2624 2867 2676 2870
rect 2732 2867 2784 2870
rect 2840 2867 2892 2870
rect 2948 2867 3000 2870
rect 3056 2867 3108 2870
rect 3164 2867 3216 2870
rect 3272 2867 3324 2870
rect 3380 2867 3432 2870
rect 3488 2867 3540 2870
rect 3596 2867 3648 2870
rect 3704 2867 3756 2870
rect 4130 2867 4182 2870
rect 4238 2867 4290 2870
rect 4346 2867 4398 2870
rect 4454 2867 4506 2870
rect 4562 2867 4614 2870
rect 4670 2867 4722 2870
rect 4778 2867 4830 2870
rect 4886 2867 4938 2870
rect 4994 2867 5046 2870
rect 5102 2867 5154 2870
rect 5210 2867 5262 2870
rect 5318 2867 5370 2870
rect 5426 2867 5478 2870
rect 5534 2867 5586 2870
rect 5642 2867 5694 2870
rect 5750 2867 5802 2870
rect 5858 2867 5910 2870
rect 5966 2867 6018 2870
rect 6074 2867 6126 2870
rect 6836 2867 6888 2870
rect 6944 2867 6996 2870
rect 7052 2867 7104 2870
rect 7160 2867 7212 2870
rect 7268 2867 7320 2870
rect 7376 2867 7428 2870
rect 7484 2867 7536 2870
rect 7592 2867 7644 2870
rect 7700 2867 7752 2870
rect 7808 2867 7860 2870
rect 7916 2867 7968 2870
rect 8024 2867 8076 2870
rect 8132 2867 8184 2870
rect 8240 2867 8292 2870
rect 8348 2867 8400 2870
rect 8456 2867 8508 2870
rect 8564 2867 8616 2870
rect 8672 2867 8724 2870
rect 8780 2867 8832 2870
rect 9206 2867 9258 2870
rect 9314 2867 9366 2870
rect 9422 2867 9474 2870
rect 9530 2867 9582 2870
rect 9638 2867 9690 2870
rect 9746 2867 9798 2870
rect 9854 2867 9906 2870
rect 9962 2867 10014 2870
rect 10070 2867 10122 2870
rect 10178 2867 10230 2870
rect 10286 2867 10338 2870
rect 10394 2867 10446 2870
rect 10502 2867 10554 2870
rect 10610 2867 10662 2870
rect 10718 2867 10770 2870
rect 10826 2867 10878 2870
rect 10934 2867 10986 2870
rect 11042 2867 11094 2870
rect 11150 2867 11202 2870
rect 1493 2672 1545 2675
rect 1601 2672 1653 2675
rect 3863 2672 3915 2675
rect 3971 2672 4023 2675
rect 6239 2672 6291 2675
rect 6347 2672 6399 2675
rect 6455 2672 6507 2675
rect 6563 2672 6615 2675
rect 6671 2672 6723 2675
rect 8939 2672 8991 2675
rect 9047 2672 9099 2675
rect 11309 2672 11361 2675
rect 11417 2672 11469 2675
rect 1493 2626 1494 2672
rect 1494 2626 1545 2672
rect 1601 2626 1653 2672
rect 3863 2626 3915 2672
rect 3971 2626 4023 2672
rect 6239 2626 6291 2672
rect 6347 2626 6399 2672
rect 6455 2626 6507 2672
rect 6563 2626 6615 2672
rect 6671 2626 6723 2672
rect 8939 2626 8991 2672
rect 9047 2626 9099 2672
rect 11309 2626 11361 2672
rect 11417 2626 11468 2672
rect 11468 2626 11469 2672
rect 1493 2623 1545 2626
rect 1601 2623 1653 2626
rect 3863 2623 3915 2626
rect 3971 2623 4023 2626
rect 6239 2623 6291 2626
rect 6347 2623 6399 2626
rect 6455 2623 6507 2626
rect 6563 2623 6615 2626
rect 6671 2623 6723 2626
rect 8939 2623 8991 2626
rect 9047 2623 9099 2626
rect 11309 2623 11361 2626
rect 11417 2623 11469 2626
rect 1760 2428 1812 2431
rect 1868 2428 1920 2431
rect 1976 2428 2028 2431
rect 2084 2428 2136 2431
rect 2192 2428 2244 2431
rect 2300 2428 2352 2431
rect 2408 2428 2460 2431
rect 2516 2428 2568 2431
rect 2624 2428 2676 2431
rect 2732 2428 2784 2431
rect 2840 2428 2892 2431
rect 2948 2428 3000 2431
rect 3056 2428 3108 2431
rect 3164 2428 3216 2431
rect 3272 2428 3324 2431
rect 3380 2428 3432 2431
rect 3488 2428 3540 2431
rect 3596 2428 3648 2431
rect 3704 2428 3756 2431
rect 4130 2428 4182 2431
rect 4238 2428 4290 2431
rect 4346 2428 4398 2431
rect 4454 2428 4506 2431
rect 4562 2428 4614 2431
rect 4670 2428 4722 2431
rect 4778 2428 4830 2431
rect 4886 2428 4938 2431
rect 4994 2428 5046 2431
rect 5102 2428 5154 2431
rect 5210 2428 5262 2431
rect 5318 2428 5370 2431
rect 5426 2428 5478 2431
rect 5534 2428 5586 2431
rect 5642 2428 5694 2431
rect 5750 2428 5802 2431
rect 5858 2428 5910 2431
rect 5966 2428 6018 2431
rect 6074 2428 6126 2431
rect 6836 2428 6888 2431
rect 6944 2428 6996 2431
rect 7052 2428 7104 2431
rect 7160 2428 7212 2431
rect 7268 2428 7320 2431
rect 7376 2428 7428 2431
rect 7484 2428 7536 2431
rect 7592 2428 7644 2431
rect 7700 2428 7752 2431
rect 7808 2428 7860 2431
rect 7916 2428 7968 2431
rect 8024 2428 8076 2431
rect 8132 2428 8184 2431
rect 8240 2428 8292 2431
rect 8348 2428 8400 2431
rect 8456 2428 8508 2431
rect 8564 2428 8616 2431
rect 8672 2428 8724 2431
rect 8780 2428 8832 2431
rect 9206 2428 9258 2431
rect 9314 2428 9366 2431
rect 9422 2428 9474 2431
rect 9530 2428 9582 2431
rect 9638 2428 9690 2431
rect 9746 2428 9798 2431
rect 9854 2428 9906 2431
rect 9962 2428 10014 2431
rect 10070 2428 10122 2431
rect 10178 2428 10230 2431
rect 10286 2428 10338 2431
rect 10394 2428 10446 2431
rect 10502 2428 10554 2431
rect 10610 2428 10662 2431
rect 10718 2428 10770 2431
rect 10826 2428 10878 2431
rect 10934 2428 10986 2431
rect 11042 2428 11094 2431
rect 11150 2428 11202 2431
rect 1760 2382 1812 2428
rect 1868 2382 1920 2428
rect 1976 2382 2028 2428
rect 2084 2382 2136 2428
rect 2192 2382 2244 2428
rect 2300 2382 2352 2428
rect 2408 2382 2460 2428
rect 2516 2382 2568 2428
rect 2624 2382 2676 2428
rect 2732 2382 2784 2428
rect 2840 2382 2892 2428
rect 2948 2382 3000 2428
rect 3056 2382 3108 2428
rect 3164 2382 3216 2428
rect 3272 2382 3324 2428
rect 3380 2382 3432 2428
rect 3488 2382 3540 2428
rect 3596 2382 3648 2428
rect 3704 2382 3756 2428
rect 4130 2382 4182 2428
rect 4238 2382 4290 2428
rect 4346 2382 4398 2428
rect 4454 2382 4506 2428
rect 4562 2382 4614 2428
rect 4670 2382 4722 2428
rect 4778 2382 4830 2428
rect 4886 2382 4938 2428
rect 4994 2382 5046 2428
rect 5102 2382 5154 2428
rect 5210 2382 5262 2428
rect 5318 2382 5370 2428
rect 5426 2382 5478 2428
rect 5534 2382 5586 2428
rect 5642 2382 5694 2428
rect 5750 2382 5802 2428
rect 5858 2382 5910 2428
rect 5966 2382 6018 2428
rect 6074 2382 6126 2428
rect 6836 2382 6888 2428
rect 6944 2382 6996 2428
rect 7052 2382 7104 2428
rect 7160 2382 7212 2428
rect 7268 2382 7320 2428
rect 7376 2382 7428 2428
rect 7484 2382 7536 2428
rect 7592 2382 7644 2428
rect 7700 2382 7752 2428
rect 7808 2382 7860 2428
rect 7916 2382 7968 2428
rect 8024 2382 8076 2428
rect 8132 2382 8184 2428
rect 8240 2382 8292 2428
rect 8348 2382 8400 2428
rect 8456 2382 8508 2428
rect 8564 2382 8616 2428
rect 8672 2382 8724 2428
rect 8780 2382 8832 2428
rect 9206 2382 9258 2428
rect 9314 2382 9366 2428
rect 9422 2382 9474 2428
rect 9530 2382 9582 2428
rect 9638 2382 9690 2428
rect 9746 2382 9798 2428
rect 9854 2382 9906 2428
rect 9962 2382 10014 2428
rect 10070 2382 10122 2428
rect 10178 2382 10230 2428
rect 10286 2382 10338 2428
rect 10394 2382 10446 2428
rect 10502 2382 10554 2428
rect 10610 2382 10662 2428
rect 10718 2382 10770 2428
rect 10826 2382 10878 2428
rect 10934 2382 10986 2428
rect 11042 2382 11094 2428
rect 11150 2382 11202 2428
rect 1760 2379 1812 2382
rect 1868 2379 1920 2382
rect 1976 2379 2028 2382
rect 2084 2379 2136 2382
rect 2192 2379 2244 2382
rect 2300 2379 2352 2382
rect 2408 2379 2460 2382
rect 2516 2379 2568 2382
rect 2624 2379 2676 2382
rect 2732 2379 2784 2382
rect 2840 2379 2892 2382
rect 2948 2379 3000 2382
rect 3056 2379 3108 2382
rect 3164 2379 3216 2382
rect 3272 2379 3324 2382
rect 3380 2379 3432 2382
rect 3488 2379 3540 2382
rect 3596 2379 3648 2382
rect 3704 2379 3756 2382
rect 4130 2379 4182 2382
rect 4238 2379 4290 2382
rect 4346 2379 4398 2382
rect 4454 2379 4506 2382
rect 4562 2379 4614 2382
rect 4670 2379 4722 2382
rect 4778 2379 4830 2382
rect 4886 2379 4938 2382
rect 4994 2379 5046 2382
rect 5102 2379 5154 2382
rect 5210 2379 5262 2382
rect 5318 2379 5370 2382
rect 5426 2379 5478 2382
rect 5534 2379 5586 2382
rect 5642 2379 5694 2382
rect 5750 2379 5802 2382
rect 5858 2379 5910 2382
rect 5966 2379 6018 2382
rect 6074 2379 6126 2382
rect 6836 2379 6888 2382
rect 6944 2379 6996 2382
rect 7052 2379 7104 2382
rect 7160 2379 7212 2382
rect 7268 2379 7320 2382
rect 7376 2379 7428 2382
rect 7484 2379 7536 2382
rect 7592 2379 7644 2382
rect 7700 2379 7752 2382
rect 7808 2379 7860 2382
rect 7916 2379 7968 2382
rect 8024 2379 8076 2382
rect 8132 2379 8184 2382
rect 8240 2379 8292 2382
rect 8348 2379 8400 2382
rect 8456 2379 8508 2382
rect 8564 2379 8616 2382
rect 8672 2379 8724 2382
rect 8780 2379 8832 2382
rect 9206 2379 9258 2382
rect 9314 2379 9366 2382
rect 9422 2379 9474 2382
rect 9530 2379 9582 2382
rect 9638 2379 9690 2382
rect 9746 2379 9798 2382
rect 9854 2379 9906 2382
rect 9962 2379 10014 2382
rect 10070 2379 10122 2382
rect 10178 2379 10230 2382
rect 10286 2379 10338 2382
rect 10394 2379 10446 2382
rect 10502 2379 10554 2382
rect 10610 2379 10662 2382
rect 10718 2379 10770 2382
rect 10826 2379 10878 2382
rect 10934 2379 10986 2382
rect 11042 2379 11094 2382
rect 11150 2379 11202 2382
rect 1493 2184 1545 2187
rect 1601 2184 1653 2187
rect 3863 2184 3915 2187
rect 3971 2184 4023 2187
rect 6239 2184 6291 2187
rect 6347 2184 6399 2187
rect 6455 2184 6507 2187
rect 6563 2184 6615 2187
rect 6671 2184 6723 2187
rect 8939 2184 8991 2187
rect 9047 2184 9099 2187
rect 11309 2184 11361 2187
rect 11417 2184 11469 2187
rect 1493 2138 1494 2184
rect 1494 2138 1545 2184
rect 1601 2138 1653 2184
rect 3863 2138 3915 2184
rect 3971 2138 4023 2184
rect 6239 2138 6291 2184
rect 6347 2138 6399 2184
rect 6455 2138 6507 2184
rect 6563 2138 6615 2184
rect 6671 2138 6723 2184
rect 8939 2138 8991 2184
rect 9047 2138 9099 2184
rect 11309 2138 11361 2184
rect 11417 2138 11468 2184
rect 11468 2138 11469 2184
rect 1493 2135 1545 2138
rect 1601 2135 1653 2138
rect 3863 2135 3915 2138
rect 3971 2135 4023 2138
rect 6239 2135 6291 2138
rect 6347 2135 6399 2138
rect 6455 2135 6507 2138
rect 6563 2135 6615 2138
rect 6671 2135 6723 2138
rect 8939 2135 8991 2138
rect 9047 2135 9099 2138
rect 11309 2135 11361 2138
rect 11417 2135 11469 2138
rect 1760 1940 1812 1943
rect 1868 1940 1920 1943
rect 1976 1940 2028 1943
rect 2084 1940 2136 1943
rect 2192 1940 2244 1943
rect 2300 1940 2352 1943
rect 2408 1940 2460 1943
rect 2516 1940 2568 1943
rect 2624 1940 2676 1943
rect 2732 1940 2784 1943
rect 2840 1940 2892 1943
rect 2948 1940 3000 1943
rect 3056 1940 3108 1943
rect 3164 1940 3216 1943
rect 3272 1940 3324 1943
rect 3380 1940 3432 1943
rect 3488 1940 3540 1943
rect 3596 1940 3648 1943
rect 3704 1940 3756 1943
rect 4130 1940 4182 1943
rect 4238 1940 4290 1943
rect 4346 1940 4398 1943
rect 4454 1940 4506 1943
rect 4562 1940 4614 1943
rect 4670 1940 4722 1943
rect 4778 1940 4830 1943
rect 4886 1940 4938 1943
rect 4994 1940 5046 1943
rect 5102 1940 5154 1943
rect 5210 1940 5262 1943
rect 5318 1940 5370 1943
rect 5426 1940 5478 1943
rect 5534 1940 5586 1943
rect 5642 1940 5694 1943
rect 5750 1940 5802 1943
rect 5858 1940 5910 1943
rect 5966 1940 6018 1943
rect 6074 1940 6126 1943
rect 6836 1940 6888 1943
rect 6944 1940 6996 1943
rect 7052 1940 7104 1943
rect 7160 1940 7212 1943
rect 7268 1940 7320 1943
rect 7376 1940 7428 1943
rect 7484 1940 7536 1943
rect 7592 1940 7644 1943
rect 7700 1940 7752 1943
rect 7808 1940 7860 1943
rect 7916 1940 7968 1943
rect 8024 1940 8076 1943
rect 8132 1940 8184 1943
rect 8240 1940 8292 1943
rect 8348 1940 8400 1943
rect 8456 1940 8508 1943
rect 8564 1940 8616 1943
rect 8672 1940 8724 1943
rect 8780 1940 8832 1943
rect 9206 1940 9258 1943
rect 9314 1940 9366 1943
rect 9422 1940 9474 1943
rect 9530 1940 9582 1943
rect 9638 1940 9690 1943
rect 9746 1940 9798 1943
rect 9854 1940 9906 1943
rect 9962 1940 10014 1943
rect 10070 1940 10122 1943
rect 10178 1940 10230 1943
rect 10286 1940 10338 1943
rect 10394 1940 10446 1943
rect 10502 1940 10554 1943
rect 10610 1940 10662 1943
rect 10718 1940 10770 1943
rect 10826 1940 10878 1943
rect 10934 1940 10986 1943
rect 11042 1940 11094 1943
rect 11150 1940 11202 1943
rect 1760 1894 1812 1940
rect 1868 1894 1920 1940
rect 1976 1894 2028 1940
rect 2084 1894 2136 1940
rect 2192 1894 2244 1940
rect 2300 1894 2352 1940
rect 2408 1894 2460 1940
rect 2516 1894 2568 1940
rect 2624 1894 2676 1940
rect 2732 1894 2784 1940
rect 2840 1894 2892 1940
rect 2948 1894 3000 1940
rect 3056 1894 3108 1940
rect 3164 1894 3216 1940
rect 3272 1894 3324 1940
rect 3380 1894 3432 1940
rect 3488 1894 3540 1940
rect 3596 1894 3648 1940
rect 3704 1894 3756 1940
rect 4130 1894 4182 1940
rect 4238 1894 4290 1940
rect 4346 1894 4398 1940
rect 4454 1894 4506 1940
rect 4562 1894 4614 1940
rect 4670 1894 4722 1940
rect 4778 1894 4830 1940
rect 4886 1894 4938 1940
rect 4994 1894 5046 1940
rect 5102 1894 5154 1940
rect 5210 1894 5262 1940
rect 5318 1894 5370 1940
rect 5426 1894 5478 1940
rect 5534 1894 5586 1940
rect 5642 1894 5694 1940
rect 5750 1894 5802 1940
rect 5858 1894 5910 1940
rect 5966 1894 6018 1940
rect 6074 1894 6126 1940
rect 6836 1894 6888 1940
rect 6944 1894 6996 1940
rect 7052 1894 7104 1940
rect 7160 1894 7212 1940
rect 7268 1894 7320 1940
rect 7376 1894 7428 1940
rect 7484 1894 7536 1940
rect 7592 1894 7644 1940
rect 7700 1894 7752 1940
rect 7808 1894 7860 1940
rect 7916 1894 7968 1940
rect 8024 1894 8076 1940
rect 8132 1894 8184 1940
rect 8240 1894 8292 1940
rect 8348 1894 8400 1940
rect 8456 1894 8508 1940
rect 8564 1894 8616 1940
rect 8672 1894 8724 1940
rect 8780 1894 8832 1940
rect 9206 1894 9258 1940
rect 9314 1894 9366 1940
rect 9422 1894 9474 1940
rect 9530 1894 9582 1940
rect 9638 1894 9690 1940
rect 9746 1894 9798 1940
rect 9854 1894 9906 1940
rect 9962 1894 10014 1940
rect 10070 1894 10122 1940
rect 10178 1894 10230 1940
rect 10286 1894 10338 1940
rect 10394 1894 10446 1940
rect 10502 1894 10554 1940
rect 10610 1894 10662 1940
rect 10718 1894 10770 1940
rect 10826 1894 10878 1940
rect 10934 1894 10986 1940
rect 11042 1894 11094 1940
rect 11150 1894 11202 1940
rect 1760 1891 1812 1894
rect 1868 1891 1920 1894
rect 1976 1891 2028 1894
rect 2084 1891 2136 1894
rect 2192 1891 2244 1894
rect 2300 1891 2352 1894
rect 2408 1891 2460 1894
rect 2516 1891 2568 1894
rect 2624 1891 2676 1894
rect 2732 1891 2784 1894
rect 2840 1891 2892 1894
rect 2948 1891 3000 1894
rect 3056 1891 3108 1894
rect 3164 1891 3216 1894
rect 3272 1891 3324 1894
rect 3380 1891 3432 1894
rect 3488 1891 3540 1894
rect 3596 1891 3648 1894
rect 3704 1891 3756 1894
rect 4130 1891 4182 1894
rect 4238 1891 4290 1894
rect 4346 1891 4398 1894
rect 4454 1891 4506 1894
rect 4562 1891 4614 1894
rect 4670 1891 4722 1894
rect 4778 1891 4830 1894
rect 4886 1891 4938 1894
rect 4994 1891 5046 1894
rect 5102 1891 5154 1894
rect 5210 1891 5262 1894
rect 5318 1891 5370 1894
rect 5426 1891 5478 1894
rect 5534 1891 5586 1894
rect 5642 1891 5694 1894
rect 5750 1891 5802 1894
rect 5858 1891 5910 1894
rect 5966 1891 6018 1894
rect 6074 1891 6126 1894
rect 6836 1891 6888 1894
rect 6944 1891 6996 1894
rect 7052 1891 7104 1894
rect 7160 1891 7212 1894
rect 7268 1891 7320 1894
rect 7376 1891 7428 1894
rect 7484 1891 7536 1894
rect 7592 1891 7644 1894
rect 7700 1891 7752 1894
rect 7808 1891 7860 1894
rect 7916 1891 7968 1894
rect 8024 1891 8076 1894
rect 8132 1891 8184 1894
rect 8240 1891 8292 1894
rect 8348 1891 8400 1894
rect 8456 1891 8508 1894
rect 8564 1891 8616 1894
rect 8672 1891 8724 1894
rect 8780 1891 8832 1894
rect 9206 1891 9258 1894
rect 9314 1891 9366 1894
rect 9422 1891 9474 1894
rect 9530 1891 9582 1894
rect 9638 1891 9690 1894
rect 9746 1891 9798 1894
rect 9854 1891 9906 1894
rect 9962 1891 10014 1894
rect 10070 1891 10122 1894
rect 10178 1891 10230 1894
rect 10286 1891 10338 1894
rect 10394 1891 10446 1894
rect 10502 1891 10554 1894
rect 10610 1891 10662 1894
rect 10718 1891 10770 1894
rect 10826 1891 10878 1894
rect 10934 1891 10986 1894
rect 11042 1891 11094 1894
rect 11150 1891 11202 1894
rect 1493 1696 1545 1699
rect 1601 1696 1653 1699
rect 3863 1696 3915 1699
rect 3971 1696 4023 1699
rect 6239 1696 6291 1699
rect 6347 1696 6399 1699
rect 6455 1696 6507 1699
rect 6563 1696 6615 1699
rect 6671 1696 6723 1699
rect 8939 1696 8991 1699
rect 9047 1696 9099 1699
rect 11309 1696 11361 1699
rect 11417 1696 11469 1699
rect 1493 1650 1494 1696
rect 1494 1650 1545 1696
rect 1601 1650 1653 1696
rect 3863 1650 3915 1696
rect 3971 1650 4023 1696
rect 6239 1650 6291 1696
rect 6347 1650 6399 1696
rect 6455 1650 6507 1696
rect 6563 1650 6615 1696
rect 6671 1650 6723 1696
rect 8939 1650 8991 1696
rect 9047 1650 9099 1696
rect 11309 1650 11361 1696
rect 11417 1650 11468 1696
rect 11468 1650 11469 1696
rect 1493 1647 1545 1650
rect 1601 1647 1653 1650
rect 3863 1647 3915 1650
rect 3971 1647 4023 1650
rect 6239 1647 6291 1650
rect 6347 1647 6399 1650
rect 6455 1647 6507 1650
rect 6563 1647 6615 1650
rect 6671 1647 6723 1650
rect 8939 1647 8991 1650
rect 9047 1647 9099 1650
rect 11309 1647 11361 1650
rect 11417 1647 11469 1650
rect 1233 1467 1285 1519
rect 1341 1467 1393 1519
rect 11569 6111 11621 6163
rect 11677 6111 11706 6163
rect 11706 6111 11729 6163
rect 11569 6003 11621 6055
rect 11677 6003 11706 6055
rect 11706 6003 11729 6055
rect 11569 5895 11621 5947
rect 11677 5895 11706 5947
rect 11706 5895 11729 5947
rect 11569 5787 11621 5839
rect 11677 5787 11706 5839
rect 11706 5787 11729 5839
rect 11569 5679 11621 5731
rect 11677 5679 11706 5731
rect 11706 5679 11729 5731
rect 11569 5571 11621 5623
rect 11677 5571 11706 5623
rect 11706 5571 11729 5623
rect 11569 5463 11621 5515
rect 11677 5463 11706 5515
rect 11706 5463 11729 5515
rect 11569 5355 11621 5407
rect 11677 5355 11706 5407
rect 11706 5355 11729 5407
rect 11569 5247 11621 5299
rect 11677 5247 11706 5299
rect 11706 5247 11729 5299
rect 11569 5139 11621 5191
rect 11677 5139 11706 5191
rect 11706 5139 11729 5191
rect 11569 5031 11621 5083
rect 11677 5031 11706 5083
rect 11706 5031 11729 5083
rect 11569 4923 11621 4975
rect 11677 4923 11706 4975
rect 11706 4923 11729 4975
rect 11569 4815 11621 4867
rect 11677 4815 11706 4867
rect 11706 4815 11729 4867
rect 11569 4707 11621 4759
rect 11677 4707 11706 4759
rect 11706 4707 11729 4759
rect 11569 4599 11621 4651
rect 11677 4599 11706 4651
rect 11706 4599 11729 4651
rect 11569 4491 11621 4543
rect 11677 4491 11706 4543
rect 11706 4491 11729 4543
rect 11569 4383 11621 4435
rect 11677 4383 11706 4435
rect 11706 4383 11729 4435
rect 11569 4275 11621 4327
rect 11677 4275 11706 4327
rect 11706 4275 11729 4327
rect 11569 4167 11621 4219
rect 11677 4167 11706 4219
rect 11706 4167 11729 4219
rect 11569 4059 11621 4111
rect 11677 4059 11706 4111
rect 11706 4059 11729 4111
rect 11569 3951 11621 4003
rect 11677 3951 11706 4003
rect 11706 3951 11729 4003
rect 11569 3843 11621 3895
rect 11677 3843 11706 3895
rect 11706 3843 11729 3895
rect 11569 3735 11621 3787
rect 11677 3735 11706 3787
rect 11706 3735 11729 3787
rect 11569 3627 11621 3679
rect 11677 3627 11706 3679
rect 11706 3627 11729 3679
rect 11569 3519 11621 3571
rect 11677 3519 11706 3571
rect 11706 3519 11729 3571
rect 11569 3411 11621 3463
rect 11677 3411 11706 3463
rect 11706 3411 11729 3463
rect 11569 3303 11621 3355
rect 11677 3303 11706 3355
rect 11706 3303 11729 3355
rect 11569 3195 11621 3247
rect 11677 3195 11706 3247
rect 11706 3195 11729 3247
rect 11569 3087 11621 3139
rect 11677 3087 11706 3139
rect 11706 3087 11729 3139
rect 11569 2979 11621 3031
rect 11677 2979 11706 3031
rect 11706 2979 11729 3031
rect 11569 2871 11621 2923
rect 11677 2871 11706 2923
rect 11706 2871 11729 2923
rect 11569 2763 11621 2815
rect 11677 2763 11706 2815
rect 11706 2763 11729 2815
rect 11569 2655 11621 2707
rect 11677 2655 11706 2707
rect 11706 2655 11729 2707
rect 11569 2547 11621 2599
rect 11677 2547 11706 2599
rect 11706 2547 11729 2599
rect 11569 2439 11621 2491
rect 11677 2439 11706 2491
rect 11706 2439 11729 2491
rect 11569 2331 11621 2383
rect 11677 2331 11706 2383
rect 11706 2331 11729 2383
rect 11569 2223 11621 2275
rect 11677 2223 11706 2275
rect 11706 2223 11729 2275
rect 11569 2115 11621 2167
rect 11677 2115 11706 2167
rect 11706 2115 11729 2167
rect 11569 2007 11621 2059
rect 11677 2007 11706 2059
rect 11706 2007 11729 2059
rect 11569 1899 11621 1951
rect 11677 1899 11706 1951
rect 11706 1899 11729 1951
rect 11569 1791 11621 1843
rect 11677 1791 11706 1843
rect 11706 1791 11729 1843
rect 11569 1683 11621 1735
rect 11677 1683 11706 1735
rect 11706 1683 11729 1735
rect 11569 1575 11621 1627
rect 11677 1575 11706 1627
rect 11706 1575 11729 1627
rect 11569 1467 11621 1519
rect 11677 1467 11729 1519
rect 1760 1452 1812 1455
rect 1868 1452 1920 1455
rect 1976 1452 2028 1455
rect 2084 1452 2136 1455
rect 2192 1452 2244 1455
rect 2300 1452 2352 1455
rect 2408 1452 2460 1455
rect 2516 1452 2568 1455
rect 2624 1452 2676 1455
rect 2732 1452 2784 1455
rect 2840 1452 2892 1455
rect 2948 1452 3000 1455
rect 3056 1452 3108 1455
rect 3164 1452 3216 1455
rect 3272 1452 3324 1455
rect 3380 1452 3432 1455
rect 3488 1452 3540 1455
rect 3596 1452 3648 1455
rect 3704 1452 3756 1455
rect 4130 1452 4182 1455
rect 4238 1452 4290 1455
rect 4346 1452 4398 1455
rect 4454 1452 4506 1455
rect 4562 1452 4614 1455
rect 4670 1452 4722 1455
rect 4778 1452 4830 1455
rect 4886 1452 4938 1455
rect 4994 1452 5046 1455
rect 5102 1452 5154 1455
rect 5210 1452 5262 1455
rect 5318 1452 5370 1455
rect 5426 1452 5478 1455
rect 5534 1452 5586 1455
rect 5642 1452 5694 1455
rect 5750 1452 5802 1455
rect 5858 1452 5910 1455
rect 5966 1452 6018 1455
rect 6074 1452 6126 1455
rect 6836 1452 6888 1455
rect 6944 1452 6996 1455
rect 7052 1452 7104 1455
rect 7160 1452 7212 1455
rect 7268 1452 7320 1455
rect 7376 1452 7428 1455
rect 7484 1452 7536 1455
rect 7592 1452 7644 1455
rect 7700 1452 7752 1455
rect 7808 1452 7860 1455
rect 7916 1452 7968 1455
rect 8024 1452 8076 1455
rect 8132 1452 8184 1455
rect 8240 1452 8292 1455
rect 8348 1452 8400 1455
rect 8456 1452 8508 1455
rect 8564 1452 8616 1455
rect 8672 1452 8724 1455
rect 8780 1452 8832 1455
rect 9206 1452 9258 1455
rect 9314 1452 9366 1455
rect 9422 1452 9474 1455
rect 9530 1452 9582 1455
rect 9638 1452 9690 1455
rect 9746 1452 9798 1455
rect 9854 1452 9906 1455
rect 9962 1452 10014 1455
rect 10070 1452 10122 1455
rect 10178 1452 10230 1455
rect 10286 1452 10338 1455
rect 10394 1452 10446 1455
rect 10502 1452 10554 1455
rect 10610 1452 10662 1455
rect 10718 1452 10770 1455
rect 10826 1452 10878 1455
rect 10934 1452 10986 1455
rect 11042 1452 11094 1455
rect 11150 1452 11202 1455
rect 1760 1406 1812 1452
rect 1868 1406 1920 1452
rect 1976 1406 2028 1452
rect 2084 1406 2136 1452
rect 2192 1406 2244 1452
rect 2300 1406 2352 1452
rect 2408 1406 2460 1452
rect 2516 1406 2568 1452
rect 2624 1406 2676 1452
rect 2732 1406 2784 1452
rect 2840 1406 2892 1452
rect 2948 1406 3000 1452
rect 3056 1406 3108 1452
rect 3164 1406 3216 1452
rect 3272 1406 3324 1452
rect 3380 1406 3432 1452
rect 3488 1406 3540 1452
rect 3596 1406 3648 1452
rect 3704 1406 3756 1452
rect 4130 1406 4182 1452
rect 4238 1406 4290 1452
rect 4346 1406 4398 1452
rect 4454 1406 4506 1452
rect 4562 1406 4614 1452
rect 4670 1406 4722 1452
rect 4778 1406 4830 1452
rect 4886 1406 4938 1452
rect 4994 1406 5046 1452
rect 5102 1406 5154 1452
rect 5210 1406 5262 1452
rect 5318 1406 5370 1452
rect 5426 1406 5478 1452
rect 5534 1406 5586 1452
rect 5642 1406 5694 1452
rect 5750 1406 5802 1452
rect 5858 1406 5910 1452
rect 5966 1406 6018 1452
rect 6074 1406 6126 1452
rect 6836 1406 6888 1452
rect 6944 1406 6996 1452
rect 7052 1406 7104 1452
rect 7160 1406 7212 1452
rect 7268 1406 7320 1452
rect 7376 1406 7428 1452
rect 7484 1406 7536 1452
rect 7592 1406 7644 1452
rect 7700 1406 7752 1452
rect 7808 1406 7860 1452
rect 7916 1406 7968 1452
rect 8024 1406 8076 1452
rect 8132 1406 8184 1452
rect 8240 1406 8292 1452
rect 8348 1406 8400 1452
rect 8456 1406 8508 1452
rect 8564 1406 8616 1452
rect 8672 1406 8724 1452
rect 8780 1406 8832 1452
rect 9206 1406 9258 1452
rect 9314 1406 9366 1452
rect 9422 1406 9474 1452
rect 9530 1406 9582 1452
rect 9638 1406 9690 1452
rect 9746 1406 9798 1452
rect 9854 1406 9906 1452
rect 9962 1406 10014 1452
rect 10070 1406 10122 1452
rect 10178 1406 10230 1452
rect 10286 1406 10338 1452
rect 10394 1406 10446 1452
rect 10502 1406 10554 1452
rect 10610 1406 10662 1452
rect 10718 1406 10770 1452
rect 10826 1406 10878 1452
rect 10934 1406 10986 1452
rect 11042 1406 11094 1452
rect 11150 1406 11202 1452
rect 1760 1403 1812 1406
rect 1868 1403 1920 1406
rect 1976 1403 2028 1406
rect 2084 1403 2136 1406
rect 2192 1403 2244 1406
rect 2300 1403 2352 1406
rect 2408 1403 2460 1406
rect 2516 1403 2568 1406
rect 2624 1403 2676 1406
rect 2732 1403 2784 1406
rect 2840 1403 2892 1406
rect 2948 1403 3000 1406
rect 3056 1403 3108 1406
rect 3164 1403 3216 1406
rect 3272 1403 3324 1406
rect 3380 1403 3432 1406
rect 3488 1403 3540 1406
rect 3596 1403 3648 1406
rect 3704 1403 3756 1406
rect 4130 1403 4182 1406
rect 4238 1403 4290 1406
rect 4346 1403 4398 1406
rect 4454 1403 4506 1406
rect 4562 1403 4614 1406
rect 4670 1403 4722 1406
rect 4778 1403 4830 1406
rect 4886 1403 4938 1406
rect 4994 1403 5046 1406
rect 5102 1403 5154 1406
rect 5210 1403 5262 1406
rect 5318 1403 5370 1406
rect 5426 1403 5478 1406
rect 5534 1403 5586 1406
rect 5642 1403 5694 1406
rect 5750 1403 5802 1406
rect 5858 1403 5910 1406
rect 5966 1403 6018 1406
rect 6074 1403 6126 1406
rect 6836 1403 6888 1406
rect 6944 1403 6996 1406
rect 7052 1403 7104 1406
rect 7160 1403 7212 1406
rect 7268 1403 7320 1406
rect 7376 1403 7428 1406
rect 7484 1403 7536 1406
rect 7592 1403 7644 1406
rect 7700 1403 7752 1406
rect 7808 1403 7860 1406
rect 7916 1403 7968 1406
rect 8024 1403 8076 1406
rect 8132 1403 8184 1406
rect 8240 1403 8292 1406
rect 8348 1403 8400 1406
rect 8456 1403 8508 1406
rect 8564 1403 8616 1406
rect 8672 1403 8724 1406
rect 8780 1403 8832 1406
rect 9206 1403 9258 1406
rect 9314 1403 9366 1406
rect 9422 1403 9474 1406
rect 9530 1403 9582 1406
rect 9638 1403 9690 1406
rect 9746 1403 9798 1406
rect 9854 1403 9906 1406
rect 9962 1403 10014 1406
rect 10070 1403 10122 1406
rect 10178 1403 10230 1406
rect 10286 1403 10338 1406
rect 10394 1403 10446 1406
rect 10502 1403 10554 1406
rect 10610 1403 10662 1406
rect 10718 1403 10770 1406
rect 10826 1403 10878 1406
rect 10934 1403 10986 1406
rect 11042 1403 11094 1406
rect 11150 1403 11202 1406
rect 12051 6711 12103 6763
rect 12159 6711 12211 6763
rect 12267 6711 12319 6763
rect 12051 6603 12103 6655
rect 12159 6603 12211 6655
rect 12267 6603 12319 6655
rect 12051 6495 12103 6547
rect 12159 6495 12211 6547
rect 12267 6495 12319 6547
rect 12051 6387 12103 6439
rect 12159 6387 12211 6439
rect 12267 6387 12319 6439
rect 12051 6279 12103 6331
rect 12159 6279 12211 6331
rect 12267 6279 12319 6331
rect 12051 6171 12103 6223
rect 12159 6171 12211 6223
rect 12267 6171 12319 6223
rect 12051 6063 12103 6115
rect 12159 6063 12211 6115
rect 12267 6063 12319 6115
rect 12051 5955 12103 6007
rect 12159 5955 12211 6007
rect 12267 5955 12319 6007
rect 12051 5847 12103 5899
rect 12159 5847 12211 5899
rect 12267 5847 12319 5899
rect 12051 5739 12103 5791
rect 12159 5739 12211 5791
rect 12267 5739 12319 5791
rect 12051 5631 12103 5683
rect 12159 5631 12211 5683
rect 12267 5631 12319 5683
rect 12051 5523 12103 5575
rect 12159 5523 12211 5575
rect 12267 5523 12319 5575
rect 12051 5415 12103 5467
rect 12159 5415 12211 5467
rect 12267 5415 12319 5467
rect 12051 5307 12103 5359
rect 12159 5307 12211 5359
rect 12267 5307 12319 5359
rect 12051 5199 12103 5251
rect 12159 5199 12211 5251
rect 12267 5199 12319 5251
rect 12051 5091 12103 5143
rect 12159 5091 12211 5143
rect 12267 5091 12319 5143
rect 12051 4983 12103 5035
rect 12159 4983 12211 5035
rect 12267 4983 12319 5035
rect 12051 4875 12103 4927
rect 12159 4875 12211 4927
rect 12267 4875 12319 4927
rect 12051 4767 12103 4819
rect 12159 4767 12211 4819
rect 12267 4767 12319 4819
rect 12051 4659 12103 4711
rect 12159 4659 12211 4711
rect 12267 4659 12319 4711
rect 12051 4551 12103 4603
rect 12159 4551 12211 4603
rect 12267 4551 12319 4603
rect 12051 4443 12103 4495
rect 12159 4443 12211 4495
rect 12267 4443 12319 4495
rect 12051 4335 12103 4387
rect 12159 4335 12211 4387
rect 12267 4335 12319 4387
rect 12051 4227 12103 4279
rect 12159 4227 12211 4279
rect 12267 4227 12319 4279
rect 12051 4119 12103 4171
rect 12159 4119 12211 4171
rect 12267 4119 12319 4171
rect 12051 4011 12103 4063
rect 12159 4011 12211 4063
rect 12267 4011 12319 4063
rect 12051 3903 12103 3955
rect 12159 3903 12211 3955
rect 12267 3903 12319 3955
rect 12051 3795 12103 3847
rect 12159 3795 12211 3847
rect 12267 3795 12319 3847
rect 12051 3687 12103 3739
rect 12159 3687 12211 3739
rect 12267 3687 12319 3739
rect 12051 3579 12103 3631
rect 12159 3579 12211 3631
rect 12267 3579 12319 3631
rect 12051 3471 12103 3523
rect 12159 3471 12211 3523
rect 12267 3471 12319 3523
rect 12051 3363 12103 3415
rect 12159 3363 12211 3415
rect 12267 3363 12319 3415
rect 12051 3255 12103 3307
rect 12159 3255 12211 3307
rect 12267 3255 12319 3307
rect 12051 3147 12103 3199
rect 12159 3147 12211 3199
rect 12267 3147 12319 3199
rect 12051 3039 12103 3091
rect 12159 3039 12211 3091
rect 12267 3039 12319 3091
rect 12051 2931 12103 2983
rect 12159 2931 12211 2983
rect 12267 2931 12319 2983
rect 12051 2823 12103 2875
rect 12159 2823 12211 2875
rect 12267 2823 12319 2875
rect 12051 2715 12103 2767
rect 12159 2715 12211 2767
rect 12267 2715 12319 2767
rect 12051 2607 12103 2659
rect 12159 2607 12211 2659
rect 12267 2607 12319 2659
rect 12051 2499 12103 2551
rect 12159 2499 12211 2551
rect 12267 2499 12319 2551
rect 12051 2391 12103 2443
rect 12159 2391 12211 2443
rect 12267 2391 12319 2443
rect 12051 2283 12103 2335
rect 12159 2283 12211 2335
rect 12267 2283 12319 2335
rect 12051 2175 12103 2227
rect 12159 2175 12211 2227
rect 12267 2175 12319 2227
rect 12051 2067 12103 2119
rect 12159 2067 12211 2119
rect 12267 2067 12319 2119
rect 12051 1959 12103 2011
rect 12159 1959 12211 2011
rect 12267 1959 12319 2011
rect 12051 1851 12103 1903
rect 12159 1851 12211 1903
rect 12267 1851 12319 1903
rect 12051 1743 12103 1795
rect 12159 1743 12211 1795
rect 12267 1743 12319 1795
rect 12051 1635 12103 1687
rect 12159 1635 12211 1687
rect 12267 1635 12319 1687
rect 12051 1527 12103 1579
rect 12159 1527 12211 1579
rect 12267 1527 12319 1579
rect 12051 1419 12103 1471
rect 12159 1419 12211 1471
rect 12267 1419 12319 1471
rect 12051 1311 12103 1363
rect 12159 1311 12211 1363
rect 12267 1311 12319 1363
rect 12051 1203 12103 1255
rect 12159 1203 12211 1255
rect 12267 1203 12319 1255
rect 12051 1095 12103 1147
rect 12159 1095 12211 1147
rect 12267 1095 12319 1147
rect 643 879 695 931
rect 751 879 803 931
rect 859 879 911 931
rect 643 771 695 823
rect 751 771 803 823
rect 859 771 911 823
rect 643 663 695 715
rect 751 663 803 715
rect 859 663 911 715
rect 1760 909 1812 961
rect 1868 909 1920 961
rect 1976 909 2028 961
rect 2084 909 2136 961
rect 2192 909 2244 961
rect 2300 909 2352 961
rect 2408 909 2460 961
rect 2516 909 2568 961
rect 2624 909 2676 961
rect 2732 909 2784 961
rect 2840 909 2892 961
rect 2948 909 3000 961
rect 3056 909 3108 961
rect 3164 909 3216 961
rect 3272 909 3324 961
rect 3380 909 3432 961
rect 3488 909 3540 961
rect 3596 909 3648 961
rect 3704 909 3756 961
rect 4130 909 4182 961
rect 4238 909 4290 961
rect 4346 909 4398 961
rect 4454 909 4506 961
rect 4562 909 4614 961
rect 4670 909 4722 961
rect 4778 909 4830 961
rect 4886 909 4938 961
rect 4994 909 5046 961
rect 5102 909 5154 961
rect 5210 909 5262 961
rect 5318 909 5370 961
rect 5426 909 5478 961
rect 5534 909 5586 961
rect 5642 909 5694 961
rect 5750 909 5802 961
rect 5858 909 5910 961
rect 5966 909 6018 961
rect 6074 909 6126 961
rect 6836 909 6888 961
rect 6944 909 6996 961
rect 7052 909 7104 961
rect 7160 909 7212 961
rect 7268 909 7320 961
rect 7376 909 7428 961
rect 7484 909 7536 961
rect 7592 909 7644 961
rect 7700 909 7752 961
rect 7808 909 7860 961
rect 7916 909 7968 961
rect 8024 909 8076 961
rect 8132 909 8184 961
rect 8240 909 8292 961
rect 8348 909 8400 961
rect 8456 909 8508 961
rect 8564 909 8616 961
rect 8672 909 8724 961
rect 8780 909 8832 961
rect 9206 909 9258 961
rect 9314 909 9366 961
rect 9422 909 9474 961
rect 9530 909 9582 961
rect 9638 909 9690 961
rect 9746 909 9798 961
rect 9854 909 9906 961
rect 9962 909 10014 961
rect 10070 909 10122 961
rect 10178 909 10230 961
rect 10286 909 10338 961
rect 10394 909 10446 961
rect 10502 909 10554 961
rect 10610 909 10662 961
rect 10718 909 10770 961
rect 10826 909 10878 961
rect 10934 909 10986 961
rect 11042 909 11094 961
rect 11150 909 11202 961
rect 1760 801 1812 853
rect 1868 801 1920 853
rect 1976 801 2028 853
rect 2084 801 2136 853
rect 2192 801 2244 853
rect 2300 801 2352 853
rect 2408 801 2460 853
rect 2516 801 2568 853
rect 2624 801 2676 853
rect 2732 801 2784 853
rect 2840 801 2892 853
rect 2948 801 3000 853
rect 3056 801 3108 853
rect 3164 801 3216 853
rect 3272 801 3324 853
rect 3380 801 3432 853
rect 3488 801 3540 853
rect 3596 801 3648 853
rect 3704 801 3756 853
rect 4130 801 4182 853
rect 4238 801 4290 853
rect 4346 801 4398 853
rect 4454 801 4506 853
rect 4562 801 4614 853
rect 4670 801 4722 853
rect 4778 801 4830 853
rect 4886 801 4938 853
rect 4994 801 5046 853
rect 5102 801 5154 853
rect 5210 801 5262 853
rect 5318 801 5370 853
rect 5426 801 5478 853
rect 5534 801 5586 853
rect 5642 801 5694 853
rect 5750 801 5802 853
rect 5858 801 5910 853
rect 5966 801 6018 853
rect 6074 801 6126 853
rect 6836 801 6888 853
rect 6944 801 6996 853
rect 7052 801 7104 853
rect 7160 801 7212 853
rect 7268 801 7320 853
rect 7376 801 7428 853
rect 7484 801 7536 853
rect 7592 801 7644 853
rect 7700 801 7752 853
rect 7808 801 7860 853
rect 7916 801 7968 853
rect 8024 801 8076 853
rect 8132 801 8184 853
rect 8240 801 8292 853
rect 8348 801 8400 853
rect 8456 801 8508 853
rect 8564 801 8616 853
rect 8672 801 8724 853
rect 8780 801 8832 853
rect 9206 801 9258 853
rect 9314 801 9366 853
rect 9422 801 9474 853
rect 9530 801 9582 853
rect 9638 801 9690 853
rect 9746 801 9798 853
rect 9854 801 9906 853
rect 9962 801 10014 853
rect 10070 801 10122 853
rect 10178 801 10230 853
rect 10286 801 10338 853
rect 10394 801 10446 853
rect 10502 801 10554 853
rect 10610 801 10662 853
rect 10718 801 10770 853
rect 10826 801 10878 853
rect 10934 801 10986 853
rect 11042 801 11094 853
rect 11150 801 11202 853
rect 1760 693 1812 745
rect 1868 693 1920 745
rect 1976 693 2028 745
rect 2084 693 2136 745
rect 2192 693 2244 745
rect 2300 693 2352 745
rect 2408 693 2460 745
rect 2516 693 2568 745
rect 2624 693 2676 745
rect 2732 693 2784 745
rect 2840 693 2892 745
rect 2948 693 3000 745
rect 3056 693 3108 745
rect 3164 693 3216 745
rect 3272 693 3324 745
rect 3380 693 3432 745
rect 3488 693 3540 745
rect 3596 693 3648 745
rect 3704 693 3756 745
rect 4130 693 4182 745
rect 4238 693 4290 745
rect 4346 693 4398 745
rect 4454 693 4506 745
rect 4562 693 4614 745
rect 4670 693 4722 745
rect 4778 693 4830 745
rect 4886 693 4938 745
rect 4994 693 5046 745
rect 5102 693 5154 745
rect 5210 693 5262 745
rect 5318 693 5370 745
rect 5426 693 5478 745
rect 5534 693 5586 745
rect 5642 693 5694 745
rect 5750 693 5802 745
rect 5858 693 5910 745
rect 5966 693 6018 745
rect 6074 693 6126 745
rect 6836 693 6888 745
rect 6944 693 6996 745
rect 7052 693 7104 745
rect 7160 693 7212 745
rect 7268 693 7320 745
rect 7376 693 7428 745
rect 7484 693 7536 745
rect 7592 693 7644 745
rect 7700 693 7752 745
rect 7808 693 7860 745
rect 7916 693 7968 745
rect 8024 693 8076 745
rect 8132 693 8184 745
rect 8240 693 8292 745
rect 8348 693 8400 745
rect 8456 693 8508 745
rect 8564 693 8616 745
rect 8672 693 8724 745
rect 8780 693 8832 745
rect 9206 693 9258 745
rect 9314 693 9366 745
rect 9422 693 9474 745
rect 9530 693 9582 745
rect 9638 693 9690 745
rect 9746 693 9798 745
rect 9854 693 9906 745
rect 9962 693 10014 745
rect 10070 693 10122 745
rect 10178 693 10230 745
rect 10286 693 10338 745
rect 10394 693 10446 745
rect 10502 693 10554 745
rect 10610 693 10662 745
rect 10718 693 10770 745
rect 10826 693 10878 745
rect 10934 693 10986 745
rect 11042 693 11094 745
rect 11150 693 11202 745
rect 12051 987 12103 1039
rect 12159 987 12211 1039
rect 12267 987 12319 1039
rect 12051 879 12103 931
rect 12159 879 12211 931
rect 12267 879 12319 931
rect 12051 771 12103 823
rect 12159 771 12211 823
rect 12267 771 12319 823
rect 12051 663 12103 715
rect 12159 663 12211 715
rect 12267 663 12319 715
rect 1493 309 1545 361
rect 1601 309 1653 361
rect 3863 309 3915 361
rect 3971 309 4023 361
rect 6239 309 6291 361
rect 6347 309 6399 361
rect 6455 309 6507 361
rect 6563 309 6615 361
rect 6671 309 6723 361
rect 8939 309 8991 361
rect 9047 309 9099 361
rect 11309 309 11361 361
rect 11417 309 11469 361
rect 1493 201 1545 253
rect 1601 201 1653 253
rect 3863 201 3915 253
rect 3971 201 4023 253
rect 6239 201 6291 253
rect 6347 201 6399 253
rect 6455 201 6507 253
rect 6563 201 6615 253
rect 6671 201 6723 253
rect 8939 201 8991 253
rect 9047 201 9099 253
rect 11309 201 11361 253
rect 11417 201 11469 253
rect 1493 93 1545 145
rect 1601 93 1653 145
rect 3863 93 3915 145
rect 3971 93 4023 145
rect 6239 93 6291 145
rect 6347 93 6399 145
rect 6455 93 6507 145
rect 6563 93 6615 145
rect 6671 93 6723 145
rect 8939 93 8991 145
rect 9047 93 9099 145
rect 11309 93 11361 145
rect 11417 93 11469 145
<< metal2 >>
rect -747 24691 1153 25617
rect -747 24639 643 24691
rect 695 24639 751 24691
rect 803 24639 859 24691
rect 911 24639 1153 24691
rect -747 24583 1153 24639
rect -747 24531 643 24583
rect 695 24531 751 24583
rect 803 24531 859 24583
rect 911 24531 1153 24583
rect -747 24475 1153 24531
rect -747 24423 643 24475
rect 695 24423 751 24475
rect 803 24423 859 24475
rect 911 24423 1153 24475
rect -747 24367 1153 24423
rect -747 24315 643 24367
rect 695 24315 751 24367
rect 803 24315 859 24367
rect 911 24315 1153 24367
rect -747 24259 1153 24315
rect -747 24207 643 24259
rect 695 24207 751 24259
rect 803 24207 859 24259
rect 911 24207 1153 24259
rect -747 24151 1153 24207
rect -747 24099 643 24151
rect 695 24099 751 24151
rect 803 24099 859 24151
rect 911 24099 1153 24151
rect -747 24043 1153 24099
rect -747 23991 643 24043
rect 695 23991 751 24043
rect 803 23991 859 24043
rect 911 23991 1153 24043
rect -747 23935 1153 23991
rect -747 23883 643 23935
rect 695 23883 751 23935
rect 803 23883 859 23935
rect 911 23883 1153 23935
rect -747 23827 1153 23883
rect -747 23775 643 23827
rect 695 23775 751 23827
rect 803 23775 859 23827
rect 911 23775 1153 23827
rect -747 23719 1153 23775
rect -747 23667 643 23719
rect 695 23667 751 23719
rect 803 23667 859 23719
rect 911 23667 1153 23719
rect -747 23611 1153 23667
rect -747 23559 643 23611
rect 695 23559 751 23611
rect 803 23559 859 23611
rect 911 23559 1153 23611
rect -747 23503 1153 23559
rect -747 23451 643 23503
rect 695 23451 751 23503
rect 803 23451 859 23503
rect 911 23451 1153 23503
rect -747 23395 1153 23451
rect -747 23343 643 23395
rect 695 23343 751 23395
rect 803 23343 859 23395
rect 911 23343 1153 23395
rect -747 23287 1153 23343
rect -747 23235 643 23287
rect 695 23235 751 23287
rect 803 23235 859 23287
rect 911 23235 1153 23287
rect -747 23179 1153 23235
rect -747 23127 643 23179
rect 695 23127 751 23179
rect 803 23127 859 23179
rect 911 23127 1153 23179
rect -747 23071 1153 23127
rect -747 23019 643 23071
rect 695 23019 751 23071
rect 803 23019 859 23071
rect 911 23019 1153 23071
rect -747 22963 1153 23019
rect -747 22911 643 22963
rect 695 22911 751 22963
rect 803 22911 859 22963
rect 911 22911 1153 22963
rect -747 22855 1153 22911
rect -747 22803 643 22855
rect 695 22803 751 22855
rect 803 22803 859 22855
rect 911 22803 1153 22855
rect -747 22747 1153 22803
rect -747 22695 643 22747
rect 695 22695 751 22747
rect 803 22695 859 22747
rect 911 22695 1153 22747
rect -747 22639 1153 22695
rect -747 22587 643 22639
rect 695 22587 751 22639
rect 803 22587 859 22639
rect 911 22587 1153 22639
rect -747 22531 1153 22587
rect -747 22479 643 22531
rect 695 22479 751 22531
rect 803 22479 859 22531
rect 911 22479 1153 22531
rect -747 22423 1153 22479
rect -747 22371 643 22423
rect 695 22371 751 22423
rect 803 22371 859 22423
rect 911 22371 1153 22423
rect -747 22315 1153 22371
rect -747 22263 643 22315
rect 695 22263 751 22315
rect 803 22263 859 22315
rect 911 22263 1153 22315
rect -747 22207 1153 22263
rect -747 22155 643 22207
rect 695 22155 751 22207
rect 803 22155 859 22207
rect 911 22155 1153 22207
rect -747 22099 1153 22155
rect -747 22047 643 22099
rect 695 22047 751 22099
rect 803 22047 859 22099
rect 911 22047 1153 22099
rect -747 21991 1153 22047
rect -747 21939 643 21991
rect 695 21939 751 21991
rect 803 21939 859 21991
rect 911 21939 1153 21991
rect -747 21883 1153 21939
rect -747 21831 643 21883
rect 695 21831 751 21883
rect 803 21831 859 21883
rect 911 21831 1153 21883
rect -747 21775 1153 21831
rect -747 21723 643 21775
rect 695 21723 751 21775
rect 803 21723 859 21775
rect 911 21723 1153 21775
rect -747 21667 1153 21723
rect -747 21615 643 21667
rect 695 21615 751 21667
rect 803 21615 859 21667
rect 911 21615 1153 21667
rect -747 21559 1153 21615
rect -747 21507 643 21559
rect 695 21507 751 21559
rect 803 21507 859 21559
rect 911 21507 1153 21559
rect -747 21451 1153 21507
rect -747 21399 643 21451
rect 695 21399 751 21451
rect 803 21399 859 21451
rect 911 21399 1153 21451
rect -747 21343 1153 21399
rect -747 21291 643 21343
rect 695 21291 751 21343
rect 803 21291 859 21343
rect 911 21291 1153 21343
rect -747 21235 1153 21291
rect -747 21183 643 21235
rect 695 21183 751 21235
rect 803 21183 859 21235
rect 911 21183 1153 21235
rect -747 21127 1153 21183
rect -747 21075 643 21127
rect 695 21075 751 21127
rect 803 21075 859 21127
rect 911 21075 1153 21127
rect -747 21019 1153 21075
rect -747 20967 643 21019
rect 695 20967 751 21019
rect 803 20967 859 21019
rect 911 20967 1153 21019
rect -747 20911 1153 20967
rect -747 20859 643 20911
rect 695 20859 751 20911
rect 803 20859 859 20911
rect 911 20859 1153 20911
rect -747 20803 1153 20859
rect -747 20751 643 20803
rect 695 20751 751 20803
rect 803 20751 859 20803
rect 911 20751 1153 20803
rect -747 20695 1153 20751
rect -747 20643 643 20695
rect 695 20643 751 20695
rect 803 20643 859 20695
rect 911 20643 1153 20695
rect -747 20587 1153 20643
rect -747 20535 643 20587
rect 695 20535 751 20587
rect 803 20535 859 20587
rect 911 20535 1153 20587
rect -747 20479 1153 20535
rect -747 20427 643 20479
rect 695 20427 751 20479
rect 803 20427 859 20479
rect 911 20427 1153 20479
rect -747 20371 1153 20427
rect -747 20319 643 20371
rect 695 20319 751 20371
rect 803 20319 859 20371
rect 911 20319 1153 20371
rect -747 20263 1153 20319
rect -747 20211 643 20263
rect 695 20211 751 20263
rect 803 20211 859 20263
rect 911 20211 1153 20263
rect -747 20155 1153 20211
rect -747 20103 643 20155
rect 695 20103 751 20155
rect 803 20103 859 20155
rect 911 20103 1153 20155
rect -747 20047 1153 20103
rect -747 19995 643 20047
rect 695 19995 751 20047
rect 803 19995 859 20047
rect 911 19995 1153 20047
rect -747 19939 1153 19995
rect -747 19887 643 19939
rect 695 19887 751 19939
rect 803 19887 859 19939
rect 911 19887 1153 19939
rect -747 19831 1153 19887
rect -747 19779 643 19831
rect 695 19779 751 19831
rect 803 19779 859 19831
rect 911 19779 1153 19831
rect -747 19723 1153 19779
rect -747 19671 643 19723
rect 695 19671 751 19723
rect 803 19671 859 19723
rect 911 19671 1153 19723
rect -747 19615 1153 19671
rect -747 19563 643 19615
rect 695 19563 751 19615
rect 803 19563 859 19615
rect 911 19563 1153 19615
rect -747 19507 1153 19563
rect -747 19455 643 19507
rect 695 19455 751 19507
rect 803 19455 859 19507
rect 911 19455 1153 19507
rect -747 19399 1153 19455
rect -747 19347 643 19399
rect 695 19347 751 19399
rect 803 19347 859 19399
rect 911 19347 1153 19399
rect -747 19291 1153 19347
rect -747 19239 643 19291
rect 695 19239 751 19291
rect 803 19239 859 19291
rect 911 19239 1153 19291
rect -747 19183 1153 19239
rect -747 19131 643 19183
rect 695 19131 751 19183
rect 803 19131 859 19183
rect 911 19131 1153 19183
rect -747 19075 1153 19131
rect -747 19023 643 19075
rect 695 19023 751 19075
rect 803 19023 859 19075
rect 911 19023 1153 19075
rect -747 18967 1153 19023
rect -747 18915 643 18967
rect 695 18915 751 18967
rect 803 18915 859 18967
rect 911 18915 1153 18967
rect -747 18859 1153 18915
rect -747 18807 643 18859
rect 695 18807 751 18859
rect 803 18807 859 18859
rect 911 18807 1153 18859
rect -747 18751 1153 18807
rect -747 18699 643 18751
rect 695 18699 751 18751
rect 803 18699 859 18751
rect 911 18699 1153 18751
rect -747 18643 1153 18699
rect -747 18591 643 18643
rect 695 18591 751 18643
rect 803 18591 859 18643
rect 911 18591 1153 18643
rect -747 18535 1153 18591
rect -747 18483 643 18535
rect 695 18483 751 18535
rect 803 18483 859 18535
rect 911 18483 1153 18535
rect -747 18427 1153 18483
rect -747 18375 643 18427
rect 695 18375 751 18427
rect 803 18375 859 18427
rect 911 18375 1153 18427
rect -747 18319 1153 18375
rect -747 18267 643 18319
rect 695 18267 751 18319
rect 803 18267 859 18319
rect 911 18267 1153 18319
rect -747 18211 1153 18267
rect -747 18159 643 18211
rect 695 18159 751 18211
rect 803 18159 859 18211
rect 911 18159 1153 18211
rect -747 18103 1153 18159
rect -747 18051 643 18103
rect 695 18051 751 18103
rect 803 18051 859 18103
rect 911 18051 1153 18103
rect -747 17995 1153 18051
rect -747 17943 643 17995
rect 695 17943 751 17995
rect 803 17943 859 17995
rect 911 17943 1153 17995
rect -747 17887 1153 17943
rect -747 17835 643 17887
rect 695 17835 751 17887
rect 803 17835 859 17887
rect 911 17835 1153 17887
rect -747 17779 1153 17835
rect -747 17727 643 17779
rect 695 17727 751 17779
rect 803 17727 859 17779
rect 911 17727 1153 17779
rect -747 17671 1153 17727
rect -747 17619 643 17671
rect 695 17619 751 17671
rect 803 17619 859 17671
rect 911 17619 1153 17671
rect -747 17563 1153 17619
rect -747 17511 643 17563
rect 695 17511 751 17563
rect 803 17511 859 17563
rect 911 17511 1153 17563
rect -747 17455 1153 17511
rect -747 17403 643 17455
rect 695 17403 751 17455
rect 803 17403 859 17455
rect 911 17403 1153 17455
rect -747 17347 1153 17403
rect -747 17295 643 17347
rect 695 17295 751 17347
rect 803 17295 859 17347
rect 911 17295 1153 17347
rect -747 17239 1153 17295
rect -747 17187 643 17239
rect 695 17187 751 17239
rect 803 17187 859 17239
rect 911 17187 1153 17239
rect -747 17131 1153 17187
rect -747 17079 643 17131
rect 695 17079 751 17131
rect 803 17079 859 17131
rect 911 17079 1153 17131
rect -747 17023 1153 17079
rect -747 16971 643 17023
rect 695 16971 751 17023
rect 803 16971 859 17023
rect 911 16971 1153 17023
rect -747 16915 1153 16971
rect -747 16863 643 16915
rect 695 16863 751 16915
rect 803 16863 859 16915
rect 911 16863 1153 16915
rect -747 16807 1153 16863
rect -747 16755 643 16807
rect 695 16755 751 16807
rect 803 16755 859 16807
rect 911 16755 1153 16807
rect -747 16699 1153 16755
rect -747 16647 643 16699
rect 695 16647 751 16699
rect 803 16647 859 16699
rect 911 16647 1153 16699
rect -747 16591 1153 16647
rect -747 16539 643 16591
rect 695 16539 751 16591
rect 803 16539 859 16591
rect 911 16539 1153 16591
rect -747 16483 1153 16539
rect -747 16431 643 16483
rect 695 16431 751 16483
rect 803 16431 859 16483
rect 911 16431 1153 16483
rect -747 16375 1153 16431
rect -747 16323 643 16375
rect 695 16323 751 16375
rect 803 16323 859 16375
rect 911 16323 1153 16375
rect -747 16267 1153 16323
rect -747 16215 643 16267
rect 695 16215 751 16267
rect 803 16215 859 16267
rect 911 16215 1153 16267
rect -747 16159 1153 16215
rect -747 16107 643 16159
rect 695 16107 751 16159
rect 803 16107 859 16159
rect 911 16107 1153 16159
rect -747 16051 1153 16107
rect -747 15999 643 16051
rect 695 15999 751 16051
rect 803 15999 859 16051
rect 911 15999 1153 16051
rect -747 15943 1153 15999
rect -747 15891 643 15943
rect 695 15891 751 15943
rect 803 15891 859 15943
rect 911 15891 1153 15943
rect -747 15835 1153 15891
rect -747 15783 643 15835
rect 695 15783 751 15835
rect 803 15783 859 15835
rect 911 15783 1153 15835
rect -747 15727 1153 15783
rect -747 15675 643 15727
rect 695 15675 751 15727
rect 803 15675 859 15727
rect 911 15675 1153 15727
rect -747 15619 1153 15675
rect -747 15567 643 15619
rect 695 15567 751 15619
rect 803 15567 859 15619
rect 911 15567 1153 15619
rect -747 15511 1153 15567
rect -747 15459 643 15511
rect 695 15459 751 15511
rect 803 15459 859 15511
rect 911 15459 1153 15511
rect -747 15403 1153 15459
rect -747 15351 643 15403
rect 695 15351 751 15403
rect 803 15351 859 15403
rect 911 15351 1153 15403
rect -747 15295 1153 15351
rect -747 15243 643 15295
rect 695 15243 751 15295
rect 803 15243 859 15295
rect 911 15243 1153 15295
rect -747 15187 1153 15243
rect -747 15135 643 15187
rect 695 15135 751 15187
rect 803 15135 859 15187
rect 911 15135 1153 15187
rect -747 15079 1153 15135
rect -747 15027 643 15079
rect 695 15027 751 15079
rect 803 15027 859 15079
rect 911 15027 1153 15079
rect -747 14971 1153 15027
rect -747 14919 643 14971
rect 695 14919 751 14971
rect 803 14919 859 14971
rect 911 14919 1153 14971
rect -747 14863 1153 14919
rect -747 14811 643 14863
rect 695 14811 751 14863
rect 803 14811 859 14863
rect 911 14811 1153 14863
rect -747 14755 1153 14811
rect -747 14703 643 14755
rect 695 14703 751 14755
rect 803 14703 859 14755
rect 911 14703 1153 14755
rect -747 14647 1153 14703
rect -747 14595 643 14647
rect 695 14595 751 14647
rect 803 14595 859 14647
rect 911 14595 1153 14647
rect -747 14539 1153 14595
rect -747 14487 643 14539
rect 695 14487 751 14539
rect 803 14487 859 14539
rect 911 14487 1153 14539
rect -747 14431 1153 14487
rect -747 14379 643 14431
rect 695 14379 751 14431
rect 803 14379 859 14431
rect 911 14379 1153 14431
rect -747 14323 1153 14379
rect -747 14271 643 14323
rect 695 14271 751 14323
rect 803 14271 859 14323
rect 911 14271 1153 14323
rect -747 14215 1153 14271
rect -747 14163 643 14215
rect 695 14163 751 14215
rect 803 14163 859 14215
rect 911 14163 1153 14215
rect -747 14107 1153 14163
rect -747 14055 643 14107
rect 695 14055 751 14107
rect 803 14055 859 14107
rect 911 14055 1153 14107
rect -747 13999 1153 14055
rect -747 13947 643 13999
rect 695 13947 751 13999
rect 803 13947 859 13999
rect 911 13947 1153 13999
rect -747 13891 1153 13947
rect -747 13839 643 13891
rect 695 13839 751 13891
rect 803 13839 859 13891
rect 911 13839 1153 13891
rect -747 13783 1153 13839
rect -747 13731 643 13783
rect 695 13731 751 13783
rect 803 13731 859 13783
rect 911 13731 1153 13783
rect -747 13675 1153 13731
rect -747 13623 643 13675
rect 695 13623 751 13675
rect 803 13623 859 13675
rect 911 13623 1153 13675
rect -747 13567 1153 13623
rect -747 13515 643 13567
rect 695 13515 751 13567
rect 803 13515 859 13567
rect 911 13515 1153 13567
rect -747 13459 1153 13515
rect -747 13407 643 13459
rect 695 13407 751 13459
rect 803 13407 859 13459
rect 911 13407 1153 13459
rect -747 13351 1153 13407
rect -747 13299 643 13351
rect 695 13299 751 13351
rect 803 13299 859 13351
rect 911 13299 1153 13351
rect -747 13243 1153 13299
rect -747 13191 643 13243
rect 695 13191 751 13243
rect 803 13191 859 13243
rect 911 13191 1153 13243
rect -747 13135 1153 13191
rect -747 13083 643 13135
rect 695 13083 751 13135
rect 803 13083 859 13135
rect 911 13083 1153 13135
rect -747 13027 1153 13083
rect -747 12975 643 13027
rect 695 12975 751 13027
rect 803 12975 859 13027
rect 911 12975 1153 13027
rect -747 12919 1153 12975
rect -747 12867 643 12919
rect 695 12867 751 12919
rect 803 12867 859 12919
rect 911 12867 1153 12919
rect -747 12811 1153 12867
rect -747 12759 643 12811
rect 695 12759 751 12811
rect 803 12759 859 12811
rect 911 12759 1153 12811
rect -747 12703 1153 12759
rect -747 12651 643 12703
rect 695 12651 751 12703
rect 803 12651 859 12703
rect 911 12651 1153 12703
rect -747 12595 1153 12651
rect -747 12543 643 12595
rect 695 12543 751 12595
rect 803 12543 859 12595
rect 911 12543 1153 12595
rect -747 12487 1153 12543
rect -747 12435 643 12487
rect 695 12435 751 12487
rect 803 12435 859 12487
rect 911 12435 1153 12487
rect -747 12379 1153 12435
rect -747 12327 643 12379
rect 695 12327 751 12379
rect 803 12327 859 12379
rect 911 12327 1153 12379
rect -747 12271 1153 12327
rect -747 12219 643 12271
rect 695 12219 751 12271
rect 803 12219 859 12271
rect 911 12219 1153 12271
rect -747 12163 1153 12219
rect -747 12111 643 12163
rect 695 12111 751 12163
rect 803 12111 859 12163
rect 911 12111 1153 12163
rect -747 12055 1153 12111
rect -747 12003 643 12055
rect 695 12003 751 12055
rect 803 12003 859 12055
rect 911 12003 1153 12055
rect -747 11947 1153 12003
rect -747 11895 643 11947
rect 695 11895 751 11947
rect 803 11895 859 11947
rect 911 11895 1153 11947
rect -747 11839 1153 11895
rect -747 11787 643 11839
rect 695 11787 751 11839
rect 803 11787 859 11839
rect 911 11787 1153 11839
rect -747 11731 1153 11787
rect -747 11679 643 11731
rect 695 11679 751 11731
rect 803 11679 859 11731
rect 911 11679 1153 11731
rect -747 11623 1153 11679
rect -747 11571 643 11623
rect 695 11571 751 11623
rect 803 11571 859 11623
rect 911 11571 1153 11623
rect -747 11515 1153 11571
rect -747 11463 643 11515
rect 695 11463 751 11515
rect 803 11463 859 11515
rect 911 11463 1153 11515
rect -747 11407 1153 11463
rect -747 11355 643 11407
rect 695 11355 751 11407
rect 803 11355 859 11407
rect 911 11355 1153 11407
rect -747 11299 1153 11355
rect -747 11247 643 11299
rect 695 11247 751 11299
rect 803 11247 859 11299
rect 911 11247 1153 11299
rect -747 11191 1153 11247
rect -747 11139 643 11191
rect 695 11139 751 11191
rect 803 11139 859 11191
rect 911 11139 1153 11191
rect -747 11083 1153 11139
rect -747 11031 643 11083
rect 695 11031 751 11083
rect 803 11031 859 11083
rect 911 11031 1153 11083
rect -747 10975 1153 11031
rect -747 10923 643 10975
rect 695 10923 751 10975
rect 803 10923 859 10975
rect 911 10923 1153 10975
rect -747 10867 1153 10923
rect -747 10815 643 10867
rect 695 10815 751 10867
rect 803 10815 859 10867
rect 911 10815 1153 10867
rect -747 10759 1153 10815
rect -747 10707 643 10759
rect 695 10707 751 10759
rect 803 10707 859 10759
rect 911 10707 1153 10759
rect -747 10651 1153 10707
rect -747 10599 643 10651
rect 695 10599 751 10651
rect 803 10599 859 10651
rect 911 10599 1153 10651
rect -747 10543 1153 10599
rect -747 10491 643 10543
rect 695 10491 751 10543
rect 803 10491 859 10543
rect 911 10491 1153 10543
rect -747 10435 1153 10491
rect -747 10383 643 10435
rect 695 10383 751 10435
rect 803 10383 859 10435
rect 911 10383 1153 10435
rect -747 10327 1153 10383
rect -747 10275 643 10327
rect 695 10275 751 10327
rect 803 10275 859 10327
rect 911 10275 1153 10327
rect -747 10219 1153 10275
rect -747 10167 643 10219
rect 695 10167 751 10219
rect 803 10167 859 10219
rect 911 10167 1153 10219
rect -747 10111 1153 10167
rect -747 10059 643 10111
rect 695 10059 751 10111
rect 803 10059 859 10111
rect 911 10059 1153 10111
rect -747 10003 1153 10059
rect -747 9951 643 10003
rect 695 9951 751 10003
rect 803 9951 859 10003
rect 911 9951 1153 10003
rect -747 9895 1153 9951
rect -747 9843 643 9895
rect 695 9843 751 9895
rect 803 9843 859 9895
rect 911 9843 1153 9895
rect -747 9787 1153 9843
rect -747 9735 643 9787
rect 695 9735 751 9787
rect 803 9735 859 9787
rect 911 9735 1153 9787
rect -747 9679 1153 9735
rect -747 9627 643 9679
rect 695 9627 751 9679
rect 803 9627 859 9679
rect 911 9627 1153 9679
rect -747 9571 1153 9627
rect -747 9519 643 9571
rect 695 9519 751 9571
rect 803 9519 859 9571
rect 911 9519 1153 9571
rect -747 9463 1153 9519
rect -747 9411 643 9463
rect 695 9411 751 9463
rect 803 9411 859 9463
rect 911 9411 1153 9463
rect -747 9355 1153 9411
rect -747 9303 643 9355
rect 695 9303 751 9355
rect 803 9303 859 9355
rect 911 9303 1153 9355
rect -747 9247 1153 9303
rect -747 9195 643 9247
rect 695 9195 751 9247
rect 803 9195 859 9247
rect 911 9195 1153 9247
rect -747 9139 1153 9195
rect -747 9087 643 9139
rect 695 9087 751 9139
rect 803 9087 859 9139
rect 911 9087 1153 9139
rect -747 9031 1153 9087
rect -747 8979 643 9031
rect 695 8979 751 9031
rect 803 8979 859 9031
rect 911 8979 1153 9031
rect -747 8923 1153 8979
rect -747 8871 643 8923
rect 695 8871 751 8923
rect 803 8871 859 8923
rect 911 8871 1153 8923
rect -747 8815 1153 8871
rect -747 8763 643 8815
rect 695 8763 751 8815
rect 803 8763 859 8815
rect 911 8763 1153 8815
rect -747 8707 1153 8763
rect -747 8655 643 8707
rect 695 8655 751 8707
rect 803 8655 859 8707
rect 911 8655 1153 8707
rect -747 8599 1153 8655
rect -747 8547 643 8599
rect 695 8547 751 8599
rect 803 8547 859 8599
rect 911 8547 1153 8599
rect -747 8491 1153 8547
rect -747 8439 643 8491
rect 695 8439 751 8491
rect 803 8439 859 8491
rect 911 8439 1153 8491
rect -747 8383 1153 8439
rect -747 8331 643 8383
rect 695 8331 751 8383
rect 803 8331 859 8383
rect 911 8331 1153 8383
rect -747 8275 1153 8331
rect -747 8223 643 8275
rect 695 8223 751 8275
rect 803 8223 859 8275
rect 911 8223 1153 8275
rect -747 8167 1153 8223
rect -747 8115 643 8167
rect 695 8115 751 8167
rect 803 8115 859 8167
rect 911 8115 1153 8167
rect -747 8059 1153 8115
rect -747 8007 643 8059
rect 695 8007 751 8059
rect 803 8007 859 8059
rect 911 8007 1153 8059
rect -747 7951 1153 8007
rect -747 7899 643 7951
rect 695 7899 751 7951
rect 803 7899 859 7951
rect 911 7899 1153 7951
rect -747 7843 1153 7899
rect -747 7791 643 7843
rect 695 7791 751 7843
rect 803 7791 859 7843
rect 911 7791 1153 7843
rect -747 7735 1153 7791
rect -747 7683 643 7735
rect 695 7683 751 7735
rect 803 7683 859 7735
rect 911 7683 1153 7735
rect -747 7627 1153 7683
rect -747 7575 643 7627
rect 695 7575 751 7627
rect 803 7575 859 7627
rect 911 7575 1153 7627
rect -747 7519 1153 7575
rect -747 7467 643 7519
rect 695 7467 751 7519
rect 803 7467 859 7519
rect 911 7467 1153 7519
rect -747 7411 1153 7467
rect -747 7359 643 7411
rect 695 7359 751 7411
rect 803 7359 859 7411
rect 911 7359 1153 7411
rect -747 7303 1153 7359
rect -747 7251 643 7303
rect 695 7251 751 7303
rect 803 7251 859 7303
rect 911 7251 1153 7303
rect -747 7195 1153 7251
rect -747 7143 643 7195
rect 695 7143 751 7195
rect 803 7143 859 7195
rect 911 7143 1153 7195
rect -747 7087 1153 7143
rect -747 7035 643 7087
rect 695 7035 751 7087
rect 803 7035 859 7087
rect 911 7035 1153 7087
rect -747 6979 1153 7035
rect -747 6927 643 6979
rect 695 6927 751 6979
rect 803 6927 859 6979
rect 911 6927 1153 6979
rect -747 6871 1153 6927
rect -747 6819 643 6871
rect 695 6819 751 6871
rect 803 6819 859 6871
rect 911 6819 1153 6871
rect -747 6763 1153 6819
rect -747 6711 643 6763
rect 695 6711 751 6763
rect 803 6711 859 6763
rect 911 6711 1153 6763
rect -747 6655 1153 6711
rect -747 6603 643 6655
rect 695 6603 751 6655
rect 803 6603 859 6655
rect 911 6603 1153 6655
rect -747 6547 1153 6603
rect -747 6495 643 6547
rect 695 6495 751 6547
rect 803 6495 859 6547
rect 911 6495 1153 6547
rect -747 6439 1153 6495
rect -747 6387 643 6439
rect 695 6387 751 6439
rect 803 6387 859 6439
rect 911 6387 1153 6439
rect -747 6331 1153 6387
rect -747 6279 643 6331
rect 695 6279 751 6331
rect 803 6279 859 6331
rect 911 6279 1153 6331
rect -747 6223 1153 6279
rect -747 6171 643 6223
rect 695 6171 751 6223
rect 803 6171 859 6223
rect 911 6171 1153 6223
rect -747 6115 1153 6171
rect -747 6063 643 6115
rect 695 6063 751 6115
rect 803 6063 859 6115
rect 911 6063 1153 6115
rect -747 6007 1153 6063
rect -747 5955 643 6007
rect 695 5955 751 6007
rect 803 5955 859 6007
rect 911 5955 1153 6007
rect -747 5899 1153 5955
rect -747 5847 643 5899
rect 695 5847 751 5899
rect 803 5847 859 5899
rect 911 5847 1153 5899
rect -747 5791 1153 5847
rect -747 5739 643 5791
rect 695 5739 751 5791
rect 803 5739 859 5791
rect 911 5739 1153 5791
rect -747 5683 1153 5739
rect -747 5631 643 5683
rect 695 5631 751 5683
rect 803 5631 859 5683
rect 911 5631 1153 5683
rect -747 5575 1153 5631
rect -747 5523 643 5575
rect 695 5523 751 5575
rect 803 5523 859 5575
rect 911 5523 1153 5575
rect -747 5467 1153 5523
rect -747 5415 643 5467
rect 695 5415 751 5467
rect 803 5415 859 5467
rect 911 5415 1153 5467
rect -747 5359 1153 5415
rect -747 5307 643 5359
rect 695 5307 751 5359
rect 803 5307 859 5359
rect 911 5307 1153 5359
rect -747 5251 1153 5307
rect -747 5199 643 5251
rect 695 5199 751 5251
rect 803 5199 859 5251
rect 911 5199 1153 5251
rect -747 5143 1153 5199
rect -747 5091 643 5143
rect 695 5091 751 5143
rect 803 5091 859 5143
rect 911 5091 1153 5143
rect -747 5035 1153 5091
rect -747 4983 643 5035
rect 695 4983 751 5035
rect 803 4983 859 5035
rect 911 4983 1153 5035
rect -747 4927 1153 4983
rect -747 4875 643 4927
rect 695 4875 751 4927
rect 803 4875 859 4927
rect 911 4875 1153 4927
rect -747 4819 1153 4875
rect -747 4767 643 4819
rect 695 4767 751 4819
rect 803 4767 859 4819
rect 911 4767 1153 4819
rect -747 4711 1153 4767
rect -747 4659 643 4711
rect 695 4659 751 4711
rect 803 4659 859 4711
rect 911 4659 1153 4711
rect -747 4603 1153 4659
rect -747 4551 643 4603
rect 695 4551 751 4603
rect 803 4551 859 4603
rect 911 4551 1153 4603
rect -747 4495 1153 4551
rect -747 4443 643 4495
rect 695 4443 751 4495
rect 803 4443 859 4495
rect 911 4443 1153 4495
rect -747 4387 1153 4443
rect -747 4335 643 4387
rect 695 4335 751 4387
rect 803 4335 859 4387
rect 911 4335 1153 4387
rect -747 4279 1153 4335
rect -747 4227 643 4279
rect 695 4227 751 4279
rect 803 4227 859 4279
rect 911 4227 1153 4279
rect -747 4171 1153 4227
rect -747 4119 643 4171
rect 695 4119 751 4171
rect 803 4119 859 4171
rect 911 4119 1153 4171
rect -747 4063 1153 4119
rect -747 4011 643 4063
rect 695 4011 751 4063
rect 803 4011 859 4063
rect 911 4011 1153 4063
rect -747 3955 1153 4011
rect -747 3903 643 3955
rect 695 3903 751 3955
rect 803 3903 859 3955
rect 911 3903 1153 3955
rect -747 3847 1153 3903
rect -747 3795 643 3847
rect 695 3795 751 3847
rect 803 3795 859 3847
rect 911 3795 1153 3847
rect -747 3739 1153 3795
rect -747 3687 643 3739
rect 695 3687 751 3739
rect 803 3687 859 3739
rect 911 3687 1153 3739
rect -747 3631 1153 3687
rect -747 3579 643 3631
rect 695 3579 751 3631
rect 803 3579 859 3631
rect 911 3579 1153 3631
rect -747 3523 1153 3579
rect -747 3471 643 3523
rect 695 3471 751 3523
rect 803 3471 859 3523
rect 911 3471 1153 3523
rect -747 3415 1153 3471
rect -747 3363 643 3415
rect 695 3363 751 3415
rect 803 3363 859 3415
rect 911 3363 1153 3415
rect -747 3307 1153 3363
rect -747 3255 643 3307
rect 695 3255 751 3307
rect 803 3255 859 3307
rect 911 3255 1153 3307
rect -747 3199 1153 3255
rect -747 3147 643 3199
rect 695 3147 751 3199
rect 803 3147 859 3199
rect 911 3147 1153 3199
rect -747 3091 1153 3147
rect -747 3039 643 3091
rect 695 3039 751 3091
rect 803 3039 859 3091
rect 911 3039 1153 3091
rect -747 2983 1153 3039
rect -747 2931 643 2983
rect 695 2931 751 2983
rect 803 2931 859 2983
rect 911 2931 1153 2983
rect -747 2875 1153 2931
rect -747 2823 643 2875
rect 695 2823 751 2875
rect 803 2823 859 2875
rect 911 2823 1153 2875
rect -747 2767 1153 2823
rect -747 2715 643 2767
rect 695 2715 751 2767
rect 803 2715 859 2767
rect 911 2715 1153 2767
rect -747 2659 1153 2715
rect -747 2607 643 2659
rect 695 2607 751 2659
rect 803 2607 859 2659
rect 911 2607 1153 2659
rect -747 2551 1153 2607
rect -747 2499 643 2551
rect 695 2499 751 2551
rect 803 2499 859 2551
rect 911 2499 1153 2551
rect -747 2443 1153 2499
rect -747 2391 643 2443
rect 695 2391 751 2443
rect 803 2391 859 2443
rect 911 2391 1153 2443
rect -747 2335 1153 2391
rect -747 2283 643 2335
rect 695 2283 751 2335
rect 803 2283 859 2335
rect 911 2283 1153 2335
rect -747 2227 1153 2283
rect -747 2175 643 2227
rect 695 2175 751 2227
rect 803 2175 859 2227
rect 911 2175 1153 2227
rect -747 2119 1153 2175
rect -747 2067 643 2119
rect 695 2067 751 2119
rect 803 2067 859 2119
rect 911 2067 1153 2119
rect -747 2011 1153 2067
rect -747 1959 643 2011
rect 695 1959 751 2011
rect 803 1959 859 2011
rect 911 1959 1153 2011
rect -747 1903 1153 1959
rect -747 1851 643 1903
rect 695 1851 751 1903
rect 803 1851 859 1903
rect 911 1851 1153 1903
rect -747 1795 1153 1851
rect -747 1743 643 1795
rect 695 1743 751 1795
rect 803 1743 859 1795
rect 911 1743 1153 1795
rect -747 1687 1153 1743
rect -747 1635 643 1687
rect 695 1635 751 1687
rect 803 1635 859 1687
rect 911 1635 1153 1687
rect -747 1579 1153 1635
rect -747 1527 643 1579
rect 695 1527 751 1579
rect 803 1527 859 1579
rect 911 1527 1153 1579
rect -747 1471 1153 1527
rect -747 1419 643 1471
rect 695 1419 751 1471
rect 803 1419 859 1471
rect 911 1419 1153 1471
rect 1213 23887 1413 25617
rect 1213 23835 1233 23887
rect 1285 23835 1341 23887
rect 1393 23835 1413 23887
rect 1213 23779 1413 23835
rect 1213 23727 1233 23779
rect 1285 23727 1341 23779
rect 1393 23727 1413 23779
rect 1213 23671 1413 23727
rect 1213 23619 1233 23671
rect 1285 23619 1341 23671
rect 1393 23619 1413 23671
rect 1213 23563 1413 23619
rect 1213 23511 1233 23563
rect 1285 23511 1341 23563
rect 1393 23511 1413 23563
rect 1213 23455 1413 23511
rect 1213 23403 1233 23455
rect 1285 23403 1341 23455
rect 1393 23403 1413 23455
rect 1213 23347 1413 23403
rect 1213 23295 1233 23347
rect 1285 23295 1341 23347
rect 1393 23295 1413 23347
rect 1213 23239 1413 23295
rect 1213 23187 1233 23239
rect 1285 23187 1341 23239
rect 1393 23187 1413 23239
rect 1213 23131 1413 23187
rect 1213 23079 1233 23131
rect 1285 23079 1341 23131
rect 1393 23079 1413 23131
rect 1213 23023 1413 23079
rect 1213 22971 1233 23023
rect 1285 22971 1341 23023
rect 1393 22971 1413 23023
rect 1213 22915 1413 22971
rect 1213 22863 1233 22915
rect 1285 22863 1341 22915
rect 1393 22863 1413 22915
rect 1213 22807 1413 22863
rect 1213 22755 1233 22807
rect 1285 22755 1341 22807
rect 1393 22755 1413 22807
rect 1213 22699 1413 22755
rect 1213 22647 1233 22699
rect 1285 22647 1341 22699
rect 1393 22647 1413 22699
rect 1213 22591 1413 22647
rect 1213 22539 1233 22591
rect 1285 22539 1341 22591
rect 1393 22539 1413 22591
rect 1213 22483 1413 22539
rect 1213 22431 1233 22483
rect 1285 22431 1341 22483
rect 1393 22431 1413 22483
rect 1213 22375 1413 22431
rect 1213 22323 1233 22375
rect 1285 22323 1341 22375
rect 1393 22323 1413 22375
rect 1213 22267 1413 22323
rect 1213 22215 1233 22267
rect 1285 22215 1341 22267
rect 1393 22215 1413 22267
rect 1213 22159 1413 22215
rect 1213 22107 1233 22159
rect 1285 22107 1341 22159
rect 1393 22107 1413 22159
rect 1213 22051 1413 22107
rect 1213 21999 1233 22051
rect 1285 21999 1341 22051
rect 1393 21999 1413 22051
rect 1213 21943 1413 21999
rect 1213 21891 1233 21943
rect 1285 21891 1341 21943
rect 1393 21891 1413 21943
rect 1213 21835 1413 21891
rect 1213 21783 1233 21835
rect 1285 21783 1341 21835
rect 1393 21783 1413 21835
rect 1213 21727 1413 21783
rect 1213 21675 1233 21727
rect 1285 21675 1341 21727
rect 1393 21675 1413 21727
rect 1213 21619 1413 21675
rect 1213 21567 1233 21619
rect 1285 21567 1341 21619
rect 1393 21567 1413 21619
rect 1213 21511 1413 21567
rect 1213 21459 1233 21511
rect 1285 21459 1341 21511
rect 1393 21459 1413 21511
rect 1213 21403 1413 21459
rect 1213 21351 1233 21403
rect 1285 21351 1341 21403
rect 1393 21351 1413 21403
rect 1213 21295 1413 21351
rect 1213 21243 1233 21295
rect 1285 21243 1341 21295
rect 1393 21243 1413 21295
rect 1213 21187 1413 21243
rect 1213 21135 1233 21187
rect 1285 21135 1341 21187
rect 1393 21135 1413 21187
rect 1213 21079 1413 21135
rect 1213 21027 1233 21079
rect 1285 21027 1341 21079
rect 1393 21027 1413 21079
rect 1213 20971 1413 21027
rect 1213 20919 1233 20971
rect 1285 20919 1341 20971
rect 1393 20919 1413 20971
rect 1213 20863 1413 20919
rect 1213 20811 1233 20863
rect 1285 20811 1341 20863
rect 1393 20811 1413 20863
rect 1213 20755 1413 20811
rect 1213 20703 1233 20755
rect 1285 20703 1341 20755
rect 1393 20703 1413 20755
rect 1213 20647 1413 20703
rect 1213 20595 1233 20647
rect 1285 20595 1341 20647
rect 1393 20595 1413 20647
rect 1213 20539 1413 20595
rect 1213 20487 1233 20539
rect 1285 20487 1341 20539
rect 1393 20487 1413 20539
rect 1213 20431 1413 20487
rect 1213 20379 1233 20431
rect 1285 20379 1341 20431
rect 1393 20379 1413 20431
rect 1213 20323 1413 20379
rect 1213 20271 1233 20323
rect 1285 20271 1341 20323
rect 1393 20271 1413 20323
rect 1213 20215 1413 20271
rect 1213 20163 1233 20215
rect 1285 20163 1341 20215
rect 1393 20163 1413 20215
rect 1213 20107 1413 20163
rect 1213 20055 1233 20107
rect 1285 20055 1341 20107
rect 1393 20055 1413 20107
rect 1213 19999 1413 20055
rect 1213 19947 1233 19999
rect 1285 19947 1341 19999
rect 1393 19947 1413 19999
rect 1213 19891 1413 19947
rect 1213 19839 1233 19891
rect 1285 19839 1341 19891
rect 1393 19839 1413 19891
rect 1213 19783 1413 19839
rect 1213 19731 1233 19783
rect 1285 19731 1341 19783
rect 1393 19731 1413 19783
rect 1213 19675 1413 19731
rect 1213 19623 1233 19675
rect 1285 19623 1341 19675
rect 1393 19623 1413 19675
rect 1213 19567 1413 19623
rect 1213 19515 1233 19567
rect 1285 19515 1341 19567
rect 1393 19515 1413 19567
rect 1213 19459 1413 19515
rect 1213 19407 1233 19459
rect 1285 19407 1341 19459
rect 1393 19407 1413 19459
rect 1213 19351 1413 19407
rect 1213 19299 1233 19351
rect 1285 19299 1341 19351
rect 1393 19299 1413 19351
rect 1213 19243 1413 19299
rect 1213 19191 1233 19243
rect 1285 19191 1341 19243
rect 1393 19191 1413 19243
rect 1213 19135 1413 19191
rect 1213 19083 1233 19135
rect 1285 19083 1341 19135
rect 1393 19083 1413 19135
rect 1213 18015 1413 19083
rect 1213 17963 1233 18015
rect 1285 17963 1341 18015
rect 1393 17963 1413 18015
rect 1213 17907 1413 17963
rect 1213 17855 1233 17907
rect 1285 17855 1341 17907
rect 1393 17855 1413 17907
rect 1213 17799 1413 17855
rect 1213 17747 1233 17799
rect 1285 17747 1341 17799
rect 1393 17747 1413 17799
rect 1213 17691 1413 17747
rect 1213 17639 1233 17691
rect 1285 17639 1341 17691
rect 1393 17639 1413 17691
rect 1213 17583 1413 17639
rect 1213 17531 1233 17583
rect 1285 17531 1341 17583
rect 1393 17531 1413 17583
rect 1213 17475 1413 17531
rect 1213 17423 1233 17475
rect 1285 17423 1341 17475
rect 1393 17423 1413 17475
rect 1213 17367 1413 17423
rect 1213 17315 1233 17367
rect 1285 17315 1341 17367
rect 1393 17315 1413 17367
rect 1213 17259 1413 17315
rect 1213 17207 1233 17259
rect 1285 17207 1341 17259
rect 1393 17207 1413 17259
rect 1213 17151 1413 17207
rect 1213 17099 1233 17151
rect 1285 17099 1341 17151
rect 1393 17099 1413 17151
rect 1213 17043 1413 17099
rect 1213 16991 1233 17043
rect 1285 16991 1341 17043
rect 1393 16991 1413 17043
rect 1213 16935 1413 16991
rect 1213 16883 1233 16935
rect 1285 16883 1341 16935
rect 1393 16883 1413 16935
rect 1213 16827 1413 16883
rect 1213 16775 1233 16827
rect 1285 16775 1341 16827
rect 1393 16775 1413 16827
rect 1213 16719 1413 16775
rect 1213 16667 1233 16719
rect 1285 16667 1341 16719
rect 1393 16667 1413 16719
rect 1213 16611 1413 16667
rect 1213 16559 1233 16611
rect 1285 16559 1341 16611
rect 1393 16559 1413 16611
rect 1213 16503 1413 16559
rect 1213 16451 1233 16503
rect 1285 16451 1341 16503
rect 1393 16451 1413 16503
rect 1213 16395 1413 16451
rect 1213 16343 1233 16395
rect 1285 16343 1341 16395
rect 1393 16343 1413 16395
rect 1213 16287 1413 16343
rect 1213 16235 1233 16287
rect 1285 16235 1341 16287
rect 1393 16235 1413 16287
rect 1213 16179 1413 16235
rect 1213 16127 1233 16179
rect 1285 16127 1341 16179
rect 1393 16127 1413 16179
rect 1213 16071 1413 16127
rect 1213 16019 1233 16071
rect 1285 16019 1341 16071
rect 1393 16019 1413 16071
rect 1213 15963 1413 16019
rect 1213 15911 1233 15963
rect 1285 15911 1341 15963
rect 1393 15911 1413 15963
rect 1213 15855 1413 15911
rect 1213 15803 1233 15855
rect 1285 15803 1341 15855
rect 1393 15803 1413 15855
rect 1213 15747 1413 15803
rect 1213 15695 1233 15747
rect 1285 15695 1341 15747
rect 1393 15695 1413 15747
rect 1213 15639 1413 15695
rect 1213 15587 1233 15639
rect 1285 15587 1341 15639
rect 1393 15587 1413 15639
rect 1213 15531 1413 15587
rect 1213 15479 1233 15531
rect 1285 15479 1341 15531
rect 1393 15479 1413 15531
rect 1213 15423 1413 15479
rect 1213 15371 1233 15423
rect 1285 15371 1341 15423
rect 1393 15371 1413 15423
rect 1213 15315 1413 15371
rect 1213 15263 1233 15315
rect 1285 15263 1341 15315
rect 1393 15263 1413 15315
rect 1213 15207 1413 15263
rect 1213 15155 1233 15207
rect 1285 15155 1341 15207
rect 1393 15155 1413 15207
rect 1213 15099 1413 15155
rect 1213 15047 1233 15099
rect 1285 15047 1341 15099
rect 1393 15047 1413 15099
rect 1213 14991 1413 15047
rect 1213 14939 1233 14991
rect 1285 14939 1341 14991
rect 1393 14939 1413 14991
rect 1213 14883 1413 14939
rect 1213 14831 1233 14883
rect 1285 14831 1341 14883
rect 1393 14831 1413 14883
rect 1213 14775 1413 14831
rect 1213 14723 1233 14775
rect 1285 14723 1341 14775
rect 1393 14723 1413 14775
rect 1213 14667 1413 14723
rect 1213 14615 1233 14667
rect 1285 14615 1341 14667
rect 1393 14615 1413 14667
rect 1213 14559 1413 14615
rect 1213 14507 1233 14559
rect 1285 14507 1341 14559
rect 1393 14507 1413 14559
rect 1213 14451 1413 14507
rect 1213 14399 1233 14451
rect 1285 14399 1341 14451
rect 1393 14399 1413 14451
rect 1213 14343 1413 14399
rect 1213 14291 1233 14343
rect 1285 14291 1341 14343
rect 1393 14291 1413 14343
rect 1213 14235 1413 14291
rect 1213 14183 1233 14235
rect 1285 14183 1341 14235
rect 1393 14183 1413 14235
rect 1213 14127 1413 14183
rect 1213 14075 1233 14127
rect 1285 14075 1341 14127
rect 1393 14075 1413 14127
rect 1213 14019 1413 14075
rect 1213 13967 1233 14019
rect 1285 13967 1341 14019
rect 1393 13967 1413 14019
rect 1213 13911 1413 13967
rect 1213 13859 1233 13911
rect 1285 13859 1341 13911
rect 1393 13859 1413 13911
rect 1213 13803 1413 13859
rect 1213 13751 1233 13803
rect 1285 13751 1341 13803
rect 1393 13751 1413 13803
rect 1213 13695 1413 13751
rect 1213 13643 1233 13695
rect 1285 13643 1341 13695
rect 1393 13643 1413 13695
rect 1213 13587 1413 13643
rect 1213 13535 1233 13587
rect 1285 13535 1341 13587
rect 1393 13535 1413 13587
rect 1213 13479 1413 13535
rect 1213 13427 1233 13479
rect 1285 13427 1341 13479
rect 1393 13427 1413 13479
rect 1213 13371 1413 13427
rect 1213 13319 1233 13371
rect 1285 13319 1341 13371
rect 1393 13319 1413 13371
rect 1213 13263 1413 13319
rect 1213 13211 1233 13263
rect 1285 13211 1341 13263
rect 1393 13211 1413 13263
rect 1213 12143 1413 13211
rect 1213 12091 1233 12143
rect 1285 12091 1341 12143
rect 1393 12091 1413 12143
rect 1213 12035 1413 12091
rect 1213 11983 1233 12035
rect 1285 11983 1341 12035
rect 1393 11983 1413 12035
rect 1213 11927 1413 11983
rect 1213 11875 1233 11927
rect 1285 11875 1341 11927
rect 1393 11875 1413 11927
rect 1213 11819 1413 11875
rect 1213 11767 1233 11819
rect 1285 11767 1341 11819
rect 1393 11767 1413 11819
rect 1213 11711 1413 11767
rect 1213 11659 1233 11711
rect 1285 11659 1341 11711
rect 1393 11659 1413 11711
rect 1213 11603 1413 11659
rect 1213 11551 1233 11603
rect 1285 11551 1341 11603
rect 1393 11551 1413 11603
rect 1213 11495 1413 11551
rect 1213 11443 1233 11495
rect 1285 11443 1341 11495
rect 1393 11443 1413 11495
rect 1213 11387 1413 11443
rect 1213 11335 1233 11387
rect 1285 11335 1341 11387
rect 1393 11335 1413 11387
rect 1213 11279 1413 11335
rect 1213 11227 1233 11279
rect 1285 11227 1341 11279
rect 1393 11227 1413 11279
rect 1213 11171 1413 11227
rect 1213 11119 1233 11171
rect 1285 11119 1341 11171
rect 1393 11119 1413 11171
rect 1213 11063 1413 11119
rect 1213 11011 1233 11063
rect 1285 11011 1341 11063
rect 1393 11011 1413 11063
rect 1213 10955 1413 11011
rect 1213 10903 1233 10955
rect 1285 10903 1341 10955
rect 1393 10903 1413 10955
rect 1213 10847 1413 10903
rect 1213 10795 1233 10847
rect 1285 10795 1341 10847
rect 1393 10795 1413 10847
rect 1213 10739 1413 10795
rect 1213 10687 1233 10739
rect 1285 10687 1341 10739
rect 1393 10687 1413 10739
rect 1213 10631 1413 10687
rect 1213 10579 1233 10631
rect 1285 10579 1341 10631
rect 1393 10579 1413 10631
rect 1213 10523 1413 10579
rect 1213 10471 1233 10523
rect 1285 10471 1341 10523
rect 1393 10471 1413 10523
rect 1213 10415 1413 10471
rect 1213 10363 1233 10415
rect 1285 10363 1341 10415
rect 1393 10363 1413 10415
rect 1213 10307 1413 10363
rect 1213 10255 1233 10307
rect 1285 10255 1341 10307
rect 1393 10255 1413 10307
rect 1213 10199 1413 10255
rect 1213 10147 1233 10199
rect 1285 10147 1341 10199
rect 1393 10147 1413 10199
rect 1213 10091 1413 10147
rect 1213 10039 1233 10091
rect 1285 10039 1341 10091
rect 1393 10039 1413 10091
rect 1213 9983 1413 10039
rect 1213 9931 1233 9983
rect 1285 9931 1341 9983
rect 1393 9931 1413 9983
rect 1213 9875 1413 9931
rect 1213 9823 1233 9875
rect 1285 9823 1341 9875
rect 1393 9823 1413 9875
rect 1213 9767 1413 9823
rect 1213 9715 1233 9767
rect 1285 9715 1341 9767
rect 1393 9715 1413 9767
rect 1213 9659 1413 9715
rect 1213 9607 1233 9659
rect 1285 9607 1341 9659
rect 1393 9607 1413 9659
rect 1213 9551 1413 9607
rect 1213 9499 1233 9551
rect 1285 9499 1341 9551
rect 1393 9499 1413 9551
rect 1213 9443 1413 9499
rect 1213 9391 1233 9443
rect 1285 9391 1341 9443
rect 1393 9391 1413 9443
rect 1213 9335 1413 9391
rect 1213 9283 1233 9335
rect 1285 9283 1341 9335
rect 1393 9283 1413 9335
rect 1213 9227 1413 9283
rect 1213 9175 1233 9227
rect 1285 9175 1341 9227
rect 1393 9175 1413 9227
rect 1213 9119 1413 9175
rect 1213 9067 1233 9119
rect 1285 9067 1341 9119
rect 1393 9067 1413 9119
rect 1213 9011 1413 9067
rect 1213 8959 1233 9011
rect 1285 8959 1341 9011
rect 1393 8959 1413 9011
rect 1213 8903 1413 8959
rect 1213 8851 1233 8903
rect 1285 8851 1341 8903
rect 1393 8851 1413 8903
rect 1213 8795 1413 8851
rect 1213 8743 1233 8795
rect 1285 8743 1341 8795
rect 1393 8743 1413 8795
rect 1213 8687 1413 8743
rect 1213 8635 1233 8687
rect 1285 8635 1341 8687
rect 1393 8635 1413 8687
rect 1213 8579 1413 8635
rect 1213 8527 1233 8579
rect 1285 8527 1341 8579
rect 1393 8527 1413 8579
rect 1213 8471 1413 8527
rect 1213 8419 1233 8471
rect 1285 8419 1341 8471
rect 1393 8419 1413 8471
rect 1213 8363 1413 8419
rect 1213 8311 1233 8363
rect 1285 8311 1341 8363
rect 1393 8311 1413 8363
rect 1213 8255 1413 8311
rect 1213 8203 1233 8255
rect 1285 8203 1341 8255
rect 1393 8203 1413 8255
rect 1213 8147 1413 8203
rect 1213 8095 1233 8147
rect 1285 8095 1341 8147
rect 1393 8095 1413 8147
rect 1213 8039 1413 8095
rect 1213 7987 1233 8039
rect 1285 7987 1341 8039
rect 1393 7987 1413 8039
rect 1213 7931 1413 7987
rect 1213 7879 1233 7931
rect 1285 7879 1341 7931
rect 1393 7879 1413 7931
rect 1213 7823 1413 7879
rect 1213 7771 1233 7823
rect 1285 7771 1341 7823
rect 1393 7771 1413 7823
rect 1213 7715 1413 7771
rect 1213 7663 1233 7715
rect 1285 7663 1341 7715
rect 1393 7663 1413 7715
rect 1213 7607 1413 7663
rect 1213 7555 1233 7607
rect 1285 7555 1341 7607
rect 1393 7555 1413 7607
rect 1213 7499 1413 7555
rect 1213 7447 1233 7499
rect 1285 7447 1341 7499
rect 1393 7447 1413 7499
rect 1213 7391 1413 7447
rect 1213 7339 1233 7391
rect 1285 7339 1341 7391
rect 1393 7339 1413 7391
rect 1213 6271 1413 7339
rect 1213 6219 1233 6271
rect 1285 6219 1341 6271
rect 1393 6219 1413 6271
rect 1213 6163 1413 6219
rect 1213 6111 1233 6163
rect 1285 6111 1341 6163
rect 1393 6111 1413 6163
rect 1213 6055 1413 6111
rect 1213 6003 1233 6055
rect 1285 6003 1341 6055
rect 1393 6003 1413 6055
rect 1213 5947 1413 6003
rect 1213 5895 1233 5947
rect 1285 5895 1341 5947
rect 1393 5895 1413 5947
rect 1213 5839 1413 5895
rect 1213 5787 1233 5839
rect 1285 5787 1341 5839
rect 1393 5787 1413 5839
rect 1213 5731 1413 5787
rect 1213 5679 1233 5731
rect 1285 5679 1341 5731
rect 1393 5679 1413 5731
rect 1213 5623 1413 5679
rect 1213 5571 1233 5623
rect 1285 5571 1341 5623
rect 1393 5571 1413 5623
rect 1213 5515 1413 5571
rect 1213 5463 1233 5515
rect 1285 5463 1341 5515
rect 1393 5463 1413 5515
rect 1213 5407 1413 5463
rect 1213 5355 1233 5407
rect 1285 5355 1341 5407
rect 1393 5355 1413 5407
rect 1213 5299 1413 5355
rect 1213 5247 1233 5299
rect 1285 5247 1341 5299
rect 1393 5247 1413 5299
rect 1213 5191 1413 5247
rect 1213 5139 1233 5191
rect 1285 5139 1341 5191
rect 1393 5139 1413 5191
rect 1213 5083 1413 5139
rect 1213 5031 1233 5083
rect 1285 5031 1341 5083
rect 1393 5031 1413 5083
rect 1213 4975 1413 5031
rect 1213 4923 1233 4975
rect 1285 4923 1341 4975
rect 1393 4923 1413 4975
rect 1213 4867 1413 4923
rect 1213 4815 1233 4867
rect 1285 4815 1341 4867
rect 1393 4815 1413 4867
rect 1213 4759 1413 4815
rect 1213 4707 1233 4759
rect 1285 4707 1341 4759
rect 1393 4707 1413 4759
rect 1213 4651 1413 4707
rect 1213 4599 1233 4651
rect 1285 4599 1341 4651
rect 1393 4599 1413 4651
rect 1213 4543 1413 4599
rect 1213 4491 1233 4543
rect 1285 4491 1341 4543
rect 1393 4491 1413 4543
rect 1213 4435 1413 4491
rect 1213 4383 1233 4435
rect 1285 4383 1341 4435
rect 1393 4383 1413 4435
rect 1213 4327 1413 4383
rect 1213 4275 1233 4327
rect 1285 4275 1341 4327
rect 1393 4275 1413 4327
rect 1213 4219 1413 4275
rect 1213 4167 1233 4219
rect 1285 4167 1341 4219
rect 1393 4167 1413 4219
rect 1213 4111 1413 4167
rect 1213 4059 1233 4111
rect 1285 4059 1341 4111
rect 1393 4059 1413 4111
rect 1213 4003 1413 4059
rect 1213 3951 1233 4003
rect 1285 3951 1341 4003
rect 1393 3951 1413 4003
rect 1213 3895 1413 3951
rect 1213 3843 1233 3895
rect 1285 3843 1341 3895
rect 1393 3843 1413 3895
rect 1213 3787 1413 3843
rect 1213 3735 1233 3787
rect 1285 3735 1341 3787
rect 1393 3735 1413 3787
rect 1213 3679 1413 3735
rect 1213 3627 1233 3679
rect 1285 3627 1341 3679
rect 1393 3627 1413 3679
rect 1213 3571 1413 3627
rect 1213 3519 1233 3571
rect 1285 3519 1341 3571
rect 1393 3519 1413 3571
rect 1213 3463 1413 3519
rect 1213 3411 1233 3463
rect 1285 3411 1341 3463
rect 1393 3411 1413 3463
rect 1213 3355 1413 3411
rect 1213 3303 1233 3355
rect 1285 3303 1341 3355
rect 1393 3303 1413 3355
rect 1213 3247 1413 3303
rect 1213 3195 1233 3247
rect 1285 3195 1341 3247
rect 1393 3195 1413 3247
rect 1213 3139 1413 3195
rect 1213 3087 1233 3139
rect 1285 3087 1341 3139
rect 1393 3087 1413 3139
rect 1213 3031 1413 3087
rect 1213 2979 1233 3031
rect 1285 2979 1341 3031
rect 1393 2979 1413 3031
rect 1213 2923 1413 2979
rect 1213 2871 1233 2923
rect 1285 2871 1341 2923
rect 1393 2871 1413 2923
rect 1213 2815 1413 2871
rect 1213 2763 1233 2815
rect 1285 2763 1341 2815
rect 1393 2763 1413 2815
rect 1213 2707 1413 2763
rect 1213 2655 1233 2707
rect 1285 2655 1341 2707
rect 1393 2655 1413 2707
rect 1213 2599 1413 2655
rect 1213 2547 1233 2599
rect 1285 2547 1341 2599
rect 1393 2547 1413 2599
rect 1213 2491 1413 2547
rect 1213 2439 1233 2491
rect 1285 2439 1341 2491
rect 1393 2439 1413 2491
rect 1213 2383 1413 2439
rect 1213 2331 1233 2383
rect 1285 2331 1341 2383
rect 1393 2331 1413 2383
rect 1213 2275 1413 2331
rect 1213 2223 1233 2275
rect 1285 2223 1341 2275
rect 1393 2223 1413 2275
rect 1213 2167 1413 2223
rect 1213 2115 1233 2167
rect 1285 2115 1341 2167
rect 1393 2115 1413 2167
rect 1213 2059 1413 2115
rect 1213 2007 1233 2059
rect 1285 2007 1341 2059
rect 1393 2007 1413 2059
rect 1213 1951 1413 2007
rect 1213 1899 1233 1951
rect 1285 1899 1341 1951
rect 1393 1899 1413 1951
rect 1213 1843 1413 1899
rect 1213 1791 1233 1843
rect 1285 1791 1341 1843
rect 1393 1791 1413 1843
rect 1213 1735 1413 1791
rect 1213 1683 1233 1735
rect 1285 1683 1341 1735
rect 1393 1683 1413 1735
rect 1213 1627 1413 1683
rect 1213 1575 1233 1627
rect 1285 1575 1341 1627
rect 1393 1575 1413 1627
rect 1213 1519 1413 1575
rect 1213 1467 1233 1519
rect 1285 1467 1341 1519
rect 1393 1467 1413 1519
rect 1213 1455 1413 1467
rect 1473 25261 1673 25617
rect 1473 25209 1493 25261
rect 1545 25209 1601 25261
rect 1653 25209 1673 25261
rect 1473 25153 1673 25209
rect 1473 25101 1493 25153
rect 1545 25101 1601 25153
rect 1653 25101 1673 25153
rect 1473 25045 1673 25101
rect 1473 24993 1493 25045
rect 1545 24993 1601 25045
rect 1653 24993 1673 25045
rect 1473 23707 1673 24993
rect 1473 23655 1493 23707
rect 1545 23655 1601 23707
rect 1653 23655 1673 23707
rect 1473 23219 1673 23655
rect 1473 23167 1493 23219
rect 1545 23167 1601 23219
rect 1653 23167 1673 23219
rect 1473 22731 1673 23167
rect 1473 22679 1493 22731
rect 1545 22679 1601 22731
rect 1653 22679 1673 22731
rect 1473 22243 1673 22679
rect 1473 22191 1493 22243
rect 1545 22191 1601 22243
rect 1653 22191 1673 22243
rect 1473 21755 1673 22191
rect 1473 21703 1493 21755
rect 1545 21703 1601 21755
rect 1653 21703 1673 21755
rect 1473 21267 1673 21703
rect 1473 21215 1493 21267
rect 1545 21215 1601 21267
rect 1653 21215 1673 21267
rect 1473 20779 1673 21215
rect 1473 20727 1493 20779
rect 1545 20727 1601 20779
rect 1653 20727 1673 20779
rect 1473 20291 1673 20727
rect 1473 20239 1493 20291
rect 1545 20239 1601 20291
rect 1653 20239 1673 20291
rect 1473 19803 1673 20239
rect 1473 19751 1493 19803
rect 1545 19751 1601 19803
rect 1653 19751 1673 19803
rect 1473 19315 1673 19751
rect 1473 19263 1493 19315
rect 1545 19263 1601 19315
rect 1653 19263 1673 19315
rect 1473 17835 1673 19263
rect 1473 17783 1493 17835
rect 1545 17783 1601 17835
rect 1653 17783 1673 17835
rect 1473 17347 1673 17783
rect 1473 17295 1493 17347
rect 1545 17295 1601 17347
rect 1653 17295 1673 17347
rect 1473 16859 1673 17295
rect 1473 16807 1493 16859
rect 1545 16807 1601 16859
rect 1653 16807 1673 16859
rect 1473 16371 1673 16807
rect 1473 16319 1493 16371
rect 1545 16319 1601 16371
rect 1653 16319 1673 16371
rect 1473 15883 1673 16319
rect 1473 15831 1493 15883
rect 1545 15831 1601 15883
rect 1653 15831 1673 15883
rect 1473 15395 1673 15831
rect 1473 15343 1493 15395
rect 1545 15343 1601 15395
rect 1653 15343 1673 15395
rect 1473 14907 1673 15343
rect 1473 14855 1493 14907
rect 1545 14855 1601 14907
rect 1653 14855 1673 14907
rect 1473 14419 1673 14855
rect 1473 14367 1493 14419
rect 1545 14367 1601 14419
rect 1653 14367 1673 14419
rect 1473 13931 1673 14367
rect 1473 13879 1493 13931
rect 1545 13879 1601 13931
rect 1653 13879 1673 13931
rect 1473 13443 1673 13879
rect 1473 13391 1493 13443
rect 1545 13391 1601 13443
rect 1653 13391 1673 13443
rect 1473 11963 1673 13391
rect 1473 11911 1493 11963
rect 1545 11911 1601 11963
rect 1653 11911 1673 11963
rect 1473 11475 1673 11911
rect 1473 11423 1493 11475
rect 1545 11423 1601 11475
rect 1653 11423 1673 11475
rect 1473 10987 1673 11423
rect 1473 10935 1493 10987
rect 1545 10935 1601 10987
rect 1653 10935 1673 10987
rect 1473 10499 1673 10935
rect 1473 10447 1493 10499
rect 1545 10447 1601 10499
rect 1653 10447 1673 10499
rect 1473 10011 1673 10447
rect 1473 9959 1493 10011
rect 1545 9959 1601 10011
rect 1653 9959 1673 10011
rect 1473 9523 1673 9959
rect 1473 9471 1493 9523
rect 1545 9471 1601 9523
rect 1653 9471 1673 9523
rect 1473 9035 1673 9471
rect 1473 8983 1493 9035
rect 1545 8983 1601 9035
rect 1653 8983 1673 9035
rect 1473 8547 1673 8983
rect 1473 8495 1493 8547
rect 1545 8495 1601 8547
rect 1653 8495 1673 8547
rect 1473 8059 1673 8495
rect 1473 8007 1493 8059
rect 1545 8007 1601 8059
rect 1653 8007 1673 8059
rect 1473 7571 1673 8007
rect 1473 7519 1493 7571
rect 1545 7519 1601 7571
rect 1653 7519 1673 7571
rect 1473 6091 1673 7519
rect 1473 6039 1493 6091
rect 1545 6039 1601 6091
rect 1653 6039 1673 6091
rect 1473 5603 1673 6039
rect 1473 5551 1493 5603
rect 1545 5551 1601 5603
rect 1653 5551 1673 5603
rect 1473 5115 1673 5551
rect 1473 5063 1493 5115
rect 1545 5063 1601 5115
rect 1653 5063 1673 5115
rect 1473 4627 1673 5063
rect 1473 4575 1493 4627
rect 1545 4575 1601 4627
rect 1653 4575 1673 4627
rect 1473 4139 1673 4575
rect 1473 4087 1493 4139
rect 1545 4087 1601 4139
rect 1653 4087 1673 4139
rect 1473 3651 1673 4087
rect 1473 3599 1493 3651
rect 1545 3599 1601 3651
rect 1653 3599 1673 3651
rect 1473 3163 1673 3599
rect 1473 3111 1493 3163
rect 1545 3111 1601 3163
rect 1653 3111 1673 3163
rect 1473 2675 1673 3111
rect 1473 2623 1493 2675
rect 1545 2623 1601 2675
rect 1653 2623 1673 2675
rect 1473 2187 1673 2623
rect 1473 2135 1493 2187
rect 1545 2135 1601 2187
rect 1653 2135 1673 2187
rect 1473 1699 1673 2135
rect 1473 1647 1493 1699
rect 1545 1647 1601 1699
rect 1653 1647 1673 1699
rect -747 1363 1153 1419
rect -747 1311 643 1363
rect 695 1311 751 1363
rect 803 1311 859 1363
rect 911 1311 1153 1363
rect -747 1255 1153 1311
rect -747 1203 643 1255
rect 695 1203 751 1255
rect 803 1203 859 1255
rect 911 1203 1153 1255
rect -747 1147 1153 1203
rect -747 1095 643 1147
rect 695 1095 751 1147
rect 803 1095 859 1147
rect 911 1095 1153 1147
rect -747 1039 1153 1095
rect -747 987 643 1039
rect 695 987 751 1039
rect 803 987 859 1039
rect 911 987 1153 1039
rect -747 931 1153 987
rect -747 879 643 931
rect 695 879 751 931
rect 803 879 859 931
rect 911 879 1153 931
rect -747 823 1153 879
rect -747 771 643 823
rect 695 771 751 823
rect 803 771 859 823
rect 911 771 1153 823
rect -747 715 1153 771
rect -747 663 643 715
rect 695 663 751 715
rect 803 663 859 715
rect 911 663 1153 715
rect -747 43 1153 663
rect 1473 361 1673 1647
rect 1473 309 1493 361
rect 1545 309 1601 361
rect 1653 309 1673 361
rect 1473 253 1673 309
rect 1473 201 1493 253
rect 1545 201 1601 253
rect 1653 201 1673 253
rect 1473 145 1673 201
rect 1473 93 1493 145
rect 1545 93 1601 145
rect 1653 93 1673 145
rect 1473 43 1673 93
rect 1733 24661 3783 25617
rect 1733 24609 1760 24661
rect 1812 24609 1868 24661
rect 1920 24609 1976 24661
rect 2028 24609 2084 24661
rect 2136 24609 2192 24661
rect 2244 24609 2300 24661
rect 2352 24609 2408 24661
rect 2460 24609 2516 24661
rect 2568 24609 2624 24661
rect 2676 24609 2732 24661
rect 2784 24609 2840 24661
rect 2892 24609 2948 24661
rect 3000 24609 3056 24661
rect 3108 24609 3164 24661
rect 3216 24609 3272 24661
rect 3324 24609 3380 24661
rect 3432 24609 3488 24661
rect 3540 24609 3596 24661
rect 3648 24609 3704 24661
rect 3756 24609 3783 24661
rect 1733 24553 3783 24609
rect 1733 24501 1760 24553
rect 1812 24501 1868 24553
rect 1920 24501 1976 24553
rect 2028 24501 2084 24553
rect 2136 24501 2192 24553
rect 2244 24501 2300 24553
rect 2352 24501 2408 24553
rect 2460 24501 2516 24553
rect 2568 24501 2624 24553
rect 2676 24501 2732 24553
rect 2784 24501 2840 24553
rect 2892 24501 2948 24553
rect 3000 24501 3056 24553
rect 3108 24501 3164 24553
rect 3216 24501 3272 24553
rect 3324 24501 3380 24553
rect 3432 24501 3488 24553
rect 3540 24501 3596 24553
rect 3648 24501 3704 24553
rect 3756 24501 3783 24553
rect 1733 24445 3783 24501
rect 1733 24393 1760 24445
rect 1812 24393 1868 24445
rect 1920 24393 1976 24445
rect 2028 24393 2084 24445
rect 2136 24393 2192 24445
rect 2244 24393 2300 24445
rect 2352 24393 2408 24445
rect 2460 24393 2516 24445
rect 2568 24393 2624 24445
rect 2676 24393 2732 24445
rect 2784 24393 2840 24445
rect 2892 24393 2948 24445
rect 3000 24393 3056 24445
rect 3108 24393 3164 24445
rect 3216 24393 3272 24445
rect 3324 24393 3380 24445
rect 3432 24393 3488 24445
rect 3540 24393 3596 24445
rect 3648 24393 3704 24445
rect 3756 24393 3783 24445
rect 1733 23951 3783 24393
rect 1733 23899 1760 23951
rect 1812 23899 1868 23951
rect 1920 23899 1976 23951
rect 2028 23899 2084 23951
rect 2136 23899 2192 23951
rect 2244 23899 2300 23951
rect 2352 23899 2408 23951
rect 2460 23899 2516 23951
rect 2568 23899 2624 23951
rect 2676 23899 2732 23951
rect 2784 23899 2840 23951
rect 2892 23899 2948 23951
rect 3000 23899 3056 23951
rect 3108 23899 3164 23951
rect 3216 23899 3272 23951
rect 3324 23899 3380 23951
rect 3432 23899 3488 23951
rect 3540 23899 3596 23951
rect 3648 23899 3704 23951
rect 3756 23899 3783 23951
rect 1733 23463 3783 23899
rect 1733 23411 1760 23463
rect 1812 23411 1868 23463
rect 1920 23411 1976 23463
rect 2028 23411 2084 23463
rect 2136 23411 2192 23463
rect 2244 23411 2300 23463
rect 2352 23411 2408 23463
rect 2460 23411 2516 23463
rect 2568 23411 2624 23463
rect 2676 23411 2732 23463
rect 2784 23411 2840 23463
rect 2892 23411 2948 23463
rect 3000 23411 3056 23463
rect 3108 23411 3164 23463
rect 3216 23411 3272 23463
rect 3324 23411 3380 23463
rect 3432 23411 3488 23463
rect 3540 23411 3596 23463
rect 3648 23411 3704 23463
rect 3756 23411 3783 23463
rect 1733 22975 3783 23411
rect 1733 22923 1760 22975
rect 1812 22923 1868 22975
rect 1920 22923 1976 22975
rect 2028 22923 2084 22975
rect 2136 22923 2192 22975
rect 2244 22923 2300 22975
rect 2352 22923 2408 22975
rect 2460 22923 2516 22975
rect 2568 22923 2624 22975
rect 2676 22923 2732 22975
rect 2784 22923 2840 22975
rect 2892 22923 2948 22975
rect 3000 22923 3056 22975
rect 3108 22923 3164 22975
rect 3216 22923 3272 22975
rect 3324 22923 3380 22975
rect 3432 22923 3488 22975
rect 3540 22923 3596 22975
rect 3648 22923 3704 22975
rect 3756 22923 3783 22975
rect 1733 22487 3783 22923
rect 1733 22435 1760 22487
rect 1812 22435 1868 22487
rect 1920 22435 1976 22487
rect 2028 22435 2084 22487
rect 2136 22435 2192 22487
rect 2244 22435 2300 22487
rect 2352 22435 2408 22487
rect 2460 22435 2516 22487
rect 2568 22435 2624 22487
rect 2676 22435 2732 22487
rect 2784 22435 2840 22487
rect 2892 22435 2948 22487
rect 3000 22435 3056 22487
rect 3108 22435 3164 22487
rect 3216 22435 3272 22487
rect 3324 22435 3380 22487
rect 3432 22435 3488 22487
rect 3540 22435 3596 22487
rect 3648 22435 3704 22487
rect 3756 22435 3783 22487
rect 1733 21999 3783 22435
rect 1733 21947 1760 21999
rect 1812 21947 1868 21999
rect 1920 21947 1976 21999
rect 2028 21947 2084 21999
rect 2136 21947 2192 21999
rect 2244 21947 2300 21999
rect 2352 21947 2408 21999
rect 2460 21947 2516 21999
rect 2568 21947 2624 21999
rect 2676 21947 2732 21999
rect 2784 21947 2840 21999
rect 2892 21947 2948 21999
rect 3000 21947 3056 21999
rect 3108 21947 3164 21999
rect 3216 21947 3272 21999
rect 3324 21947 3380 21999
rect 3432 21947 3488 21999
rect 3540 21947 3596 21999
rect 3648 21947 3704 21999
rect 3756 21947 3783 21999
rect 1733 21511 3783 21947
rect 1733 21459 1760 21511
rect 1812 21459 1868 21511
rect 1920 21459 1976 21511
rect 2028 21459 2084 21511
rect 2136 21459 2192 21511
rect 2244 21459 2300 21511
rect 2352 21459 2408 21511
rect 2460 21459 2516 21511
rect 2568 21459 2624 21511
rect 2676 21459 2732 21511
rect 2784 21459 2840 21511
rect 2892 21459 2948 21511
rect 3000 21459 3056 21511
rect 3108 21459 3164 21511
rect 3216 21459 3272 21511
rect 3324 21459 3380 21511
rect 3432 21459 3488 21511
rect 3540 21459 3596 21511
rect 3648 21459 3704 21511
rect 3756 21459 3783 21511
rect 1733 21023 3783 21459
rect 1733 20971 1760 21023
rect 1812 20971 1868 21023
rect 1920 20971 1976 21023
rect 2028 20971 2084 21023
rect 2136 20971 2192 21023
rect 2244 20971 2300 21023
rect 2352 20971 2408 21023
rect 2460 20971 2516 21023
rect 2568 20971 2624 21023
rect 2676 20971 2732 21023
rect 2784 20971 2840 21023
rect 2892 20971 2948 21023
rect 3000 20971 3056 21023
rect 3108 20971 3164 21023
rect 3216 20971 3272 21023
rect 3324 20971 3380 21023
rect 3432 20971 3488 21023
rect 3540 20971 3596 21023
rect 3648 20971 3704 21023
rect 3756 20971 3783 21023
rect 1733 20535 3783 20971
rect 1733 20483 1760 20535
rect 1812 20483 1868 20535
rect 1920 20483 1976 20535
rect 2028 20483 2084 20535
rect 2136 20483 2192 20535
rect 2244 20483 2300 20535
rect 2352 20483 2408 20535
rect 2460 20483 2516 20535
rect 2568 20483 2624 20535
rect 2676 20483 2732 20535
rect 2784 20483 2840 20535
rect 2892 20483 2948 20535
rect 3000 20483 3056 20535
rect 3108 20483 3164 20535
rect 3216 20483 3272 20535
rect 3324 20483 3380 20535
rect 3432 20483 3488 20535
rect 3540 20483 3596 20535
rect 3648 20483 3704 20535
rect 3756 20483 3783 20535
rect 1733 20047 3783 20483
rect 1733 19995 1760 20047
rect 1812 19995 1868 20047
rect 1920 19995 1976 20047
rect 2028 19995 2084 20047
rect 2136 19995 2192 20047
rect 2244 19995 2300 20047
rect 2352 19995 2408 20047
rect 2460 19995 2516 20047
rect 2568 19995 2624 20047
rect 2676 19995 2732 20047
rect 2784 19995 2840 20047
rect 2892 19995 2948 20047
rect 3000 19995 3056 20047
rect 3108 19995 3164 20047
rect 3216 19995 3272 20047
rect 3324 19995 3380 20047
rect 3432 19995 3488 20047
rect 3540 19995 3596 20047
rect 3648 19995 3704 20047
rect 3756 19995 3783 20047
rect 1733 19559 3783 19995
rect 1733 19507 1760 19559
rect 1812 19507 1868 19559
rect 1920 19507 1976 19559
rect 2028 19507 2084 19559
rect 2136 19507 2192 19559
rect 2244 19507 2300 19559
rect 2352 19507 2408 19559
rect 2460 19507 2516 19559
rect 2568 19507 2624 19559
rect 2676 19507 2732 19559
rect 2784 19507 2840 19559
rect 2892 19507 2948 19559
rect 3000 19507 3056 19559
rect 3108 19507 3164 19559
rect 3216 19507 3272 19559
rect 3324 19507 3380 19559
rect 3432 19507 3488 19559
rect 3540 19507 3596 19559
rect 3648 19507 3704 19559
rect 3756 19507 3783 19559
rect 1733 19071 3783 19507
rect 1733 19019 1760 19071
rect 1812 19019 1868 19071
rect 1920 19019 1976 19071
rect 2028 19019 2084 19071
rect 2136 19019 2192 19071
rect 2244 19019 2300 19071
rect 2352 19019 2408 19071
rect 2460 19019 2516 19071
rect 2568 19019 2624 19071
rect 2676 19019 2732 19071
rect 2784 19019 2840 19071
rect 2892 19019 2948 19071
rect 3000 19019 3056 19071
rect 3108 19019 3164 19071
rect 3216 19019 3272 19071
rect 3324 19019 3380 19071
rect 3432 19019 3488 19071
rect 3540 19019 3596 19071
rect 3648 19019 3704 19071
rect 3756 19019 3783 19071
rect 1733 18629 3783 19019
rect 1733 18577 1760 18629
rect 1812 18577 1868 18629
rect 1920 18577 1976 18629
rect 2028 18577 2084 18629
rect 2136 18577 2192 18629
rect 2244 18577 2300 18629
rect 2352 18577 2408 18629
rect 2460 18577 2516 18629
rect 2568 18577 2624 18629
rect 2676 18577 2732 18629
rect 2784 18577 2840 18629
rect 2892 18577 2948 18629
rect 3000 18577 3056 18629
rect 3108 18577 3164 18629
rect 3216 18577 3272 18629
rect 3324 18577 3380 18629
rect 3432 18577 3488 18629
rect 3540 18577 3596 18629
rect 3648 18577 3704 18629
rect 3756 18577 3783 18629
rect 1733 18521 3783 18577
rect 1733 18469 1760 18521
rect 1812 18469 1868 18521
rect 1920 18469 1976 18521
rect 2028 18469 2084 18521
rect 2136 18469 2192 18521
rect 2244 18469 2300 18521
rect 2352 18469 2408 18521
rect 2460 18469 2516 18521
rect 2568 18469 2624 18521
rect 2676 18469 2732 18521
rect 2784 18469 2840 18521
rect 2892 18469 2948 18521
rect 3000 18469 3056 18521
rect 3108 18469 3164 18521
rect 3216 18469 3272 18521
rect 3324 18469 3380 18521
rect 3432 18469 3488 18521
rect 3540 18469 3596 18521
rect 3648 18469 3704 18521
rect 3756 18469 3783 18521
rect 1733 18079 3783 18469
rect 1733 18027 1760 18079
rect 1812 18027 1868 18079
rect 1920 18027 1976 18079
rect 2028 18027 2084 18079
rect 2136 18027 2192 18079
rect 2244 18027 2300 18079
rect 2352 18027 2408 18079
rect 2460 18027 2516 18079
rect 2568 18027 2624 18079
rect 2676 18027 2732 18079
rect 2784 18027 2840 18079
rect 2892 18027 2948 18079
rect 3000 18027 3056 18079
rect 3108 18027 3164 18079
rect 3216 18027 3272 18079
rect 3324 18027 3380 18079
rect 3432 18027 3488 18079
rect 3540 18027 3596 18079
rect 3648 18027 3704 18079
rect 3756 18027 3783 18079
rect 1733 17591 3783 18027
rect 1733 17539 1760 17591
rect 1812 17539 1868 17591
rect 1920 17539 1976 17591
rect 2028 17539 2084 17591
rect 2136 17539 2192 17591
rect 2244 17539 2300 17591
rect 2352 17539 2408 17591
rect 2460 17539 2516 17591
rect 2568 17539 2624 17591
rect 2676 17539 2732 17591
rect 2784 17539 2840 17591
rect 2892 17539 2948 17591
rect 3000 17539 3056 17591
rect 3108 17539 3164 17591
rect 3216 17539 3272 17591
rect 3324 17539 3380 17591
rect 3432 17539 3488 17591
rect 3540 17539 3596 17591
rect 3648 17539 3704 17591
rect 3756 17539 3783 17591
rect 1733 17103 3783 17539
rect 1733 17051 1760 17103
rect 1812 17051 1868 17103
rect 1920 17051 1976 17103
rect 2028 17051 2084 17103
rect 2136 17051 2192 17103
rect 2244 17051 2300 17103
rect 2352 17051 2408 17103
rect 2460 17051 2516 17103
rect 2568 17051 2624 17103
rect 2676 17051 2732 17103
rect 2784 17051 2840 17103
rect 2892 17051 2948 17103
rect 3000 17051 3056 17103
rect 3108 17051 3164 17103
rect 3216 17051 3272 17103
rect 3324 17051 3380 17103
rect 3432 17051 3488 17103
rect 3540 17051 3596 17103
rect 3648 17051 3704 17103
rect 3756 17051 3783 17103
rect 1733 16615 3783 17051
rect 1733 16563 1760 16615
rect 1812 16563 1868 16615
rect 1920 16563 1976 16615
rect 2028 16563 2084 16615
rect 2136 16563 2192 16615
rect 2244 16563 2300 16615
rect 2352 16563 2408 16615
rect 2460 16563 2516 16615
rect 2568 16563 2624 16615
rect 2676 16563 2732 16615
rect 2784 16563 2840 16615
rect 2892 16563 2948 16615
rect 3000 16563 3056 16615
rect 3108 16563 3164 16615
rect 3216 16563 3272 16615
rect 3324 16563 3380 16615
rect 3432 16563 3488 16615
rect 3540 16563 3596 16615
rect 3648 16563 3704 16615
rect 3756 16563 3783 16615
rect 1733 16127 3783 16563
rect 1733 16075 1760 16127
rect 1812 16075 1868 16127
rect 1920 16075 1976 16127
rect 2028 16075 2084 16127
rect 2136 16075 2192 16127
rect 2244 16075 2300 16127
rect 2352 16075 2408 16127
rect 2460 16075 2516 16127
rect 2568 16075 2624 16127
rect 2676 16075 2732 16127
rect 2784 16075 2840 16127
rect 2892 16075 2948 16127
rect 3000 16075 3056 16127
rect 3108 16075 3164 16127
rect 3216 16075 3272 16127
rect 3324 16075 3380 16127
rect 3432 16075 3488 16127
rect 3540 16075 3596 16127
rect 3648 16075 3704 16127
rect 3756 16075 3783 16127
rect 1733 15639 3783 16075
rect 1733 15587 1760 15639
rect 1812 15587 1868 15639
rect 1920 15587 1976 15639
rect 2028 15587 2084 15639
rect 2136 15587 2192 15639
rect 2244 15587 2300 15639
rect 2352 15587 2408 15639
rect 2460 15587 2516 15639
rect 2568 15587 2624 15639
rect 2676 15587 2732 15639
rect 2784 15587 2840 15639
rect 2892 15587 2948 15639
rect 3000 15587 3056 15639
rect 3108 15587 3164 15639
rect 3216 15587 3272 15639
rect 3324 15587 3380 15639
rect 3432 15587 3488 15639
rect 3540 15587 3596 15639
rect 3648 15587 3704 15639
rect 3756 15587 3783 15639
rect 1733 15151 3783 15587
rect 1733 15099 1760 15151
rect 1812 15099 1868 15151
rect 1920 15099 1976 15151
rect 2028 15099 2084 15151
rect 2136 15099 2192 15151
rect 2244 15099 2300 15151
rect 2352 15099 2408 15151
rect 2460 15099 2516 15151
rect 2568 15099 2624 15151
rect 2676 15099 2732 15151
rect 2784 15099 2840 15151
rect 2892 15099 2948 15151
rect 3000 15099 3056 15151
rect 3108 15099 3164 15151
rect 3216 15099 3272 15151
rect 3324 15099 3380 15151
rect 3432 15099 3488 15151
rect 3540 15099 3596 15151
rect 3648 15099 3704 15151
rect 3756 15099 3783 15151
rect 1733 14663 3783 15099
rect 1733 14611 1760 14663
rect 1812 14611 1868 14663
rect 1920 14611 1976 14663
rect 2028 14611 2084 14663
rect 2136 14611 2192 14663
rect 2244 14611 2300 14663
rect 2352 14611 2408 14663
rect 2460 14611 2516 14663
rect 2568 14611 2624 14663
rect 2676 14611 2732 14663
rect 2784 14611 2840 14663
rect 2892 14611 2948 14663
rect 3000 14611 3056 14663
rect 3108 14611 3164 14663
rect 3216 14611 3272 14663
rect 3324 14611 3380 14663
rect 3432 14611 3488 14663
rect 3540 14611 3596 14663
rect 3648 14611 3704 14663
rect 3756 14611 3783 14663
rect 1733 14175 3783 14611
rect 1733 14123 1760 14175
rect 1812 14123 1868 14175
rect 1920 14123 1976 14175
rect 2028 14123 2084 14175
rect 2136 14123 2192 14175
rect 2244 14123 2300 14175
rect 2352 14123 2408 14175
rect 2460 14123 2516 14175
rect 2568 14123 2624 14175
rect 2676 14123 2732 14175
rect 2784 14123 2840 14175
rect 2892 14123 2948 14175
rect 3000 14123 3056 14175
rect 3108 14123 3164 14175
rect 3216 14123 3272 14175
rect 3324 14123 3380 14175
rect 3432 14123 3488 14175
rect 3540 14123 3596 14175
rect 3648 14123 3704 14175
rect 3756 14123 3783 14175
rect 1733 13687 3783 14123
rect 1733 13635 1760 13687
rect 1812 13635 1868 13687
rect 1920 13635 1976 13687
rect 2028 13635 2084 13687
rect 2136 13635 2192 13687
rect 2244 13635 2300 13687
rect 2352 13635 2408 13687
rect 2460 13635 2516 13687
rect 2568 13635 2624 13687
rect 2676 13635 2732 13687
rect 2784 13635 2840 13687
rect 2892 13635 2948 13687
rect 3000 13635 3056 13687
rect 3108 13635 3164 13687
rect 3216 13635 3272 13687
rect 3324 13635 3380 13687
rect 3432 13635 3488 13687
rect 3540 13635 3596 13687
rect 3648 13635 3704 13687
rect 3756 13635 3783 13687
rect 1733 13199 3783 13635
rect 1733 13147 1760 13199
rect 1812 13147 1868 13199
rect 1920 13147 1976 13199
rect 2028 13147 2084 13199
rect 2136 13147 2192 13199
rect 2244 13147 2300 13199
rect 2352 13147 2408 13199
rect 2460 13147 2516 13199
rect 2568 13147 2624 13199
rect 2676 13147 2732 13199
rect 2784 13147 2840 13199
rect 2892 13147 2948 13199
rect 3000 13147 3056 13199
rect 3108 13147 3164 13199
rect 3216 13147 3272 13199
rect 3324 13147 3380 13199
rect 3432 13147 3488 13199
rect 3540 13147 3596 13199
rect 3648 13147 3704 13199
rect 3756 13147 3783 13199
rect 1733 12757 3783 13147
rect 1733 12705 1760 12757
rect 1812 12705 1868 12757
rect 1920 12705 1976 12757
rect 2028 12705 2084 12757
rect 2136 12705 2192 12757
rect 2244 12705 2300 12757
rect 2352 12705 2408 12757
rect 2460 12705 2516 12757
rect 2568 12705 2624 12757
rect 2676 12705 2732 12757
rect 2784 12705 2840 12757
rect 2892 12705 2948 12757
rect 3000 12705 3056 12757
rect 3108 12705 3164 12757
rect 3216 12705 3272 12757
rect 3324 12705 3380 12757
rect 3432 12705 3488 12757
rect 3540 12705 3596 12757
rect 3648 12705 3704 12757
rect 3756 12705 3783 12757
rect 1733 12649 3783 12705
rect 1733 12597 1760 12649
rect 1812 12597 1868 12649
rect 1920 12597 1976 12649
rect 2028 12597 2084 12649
rect 2136 12597 2192 12649
rect 2244 12597 2300 12649
rect 2352 12597 2408 12649
rect 2460 12597 2516 12649
rect 2568 12597 2624 12649
rect 2676 12597 2732 12649
rect 2784 12597 2840 12649
rect 2892 12597 2948 12649
rect 3000 12597 3056 12649
rect 3108 12597 3164 12649
rect 3216 12597 3272 12649
rect 3324 12597 3380 12649
rect 3432 12597 3488 12649
rect 3540 12597 3596 12649
rect 3648 12597 3704 12649
rect 3756 12597 3783 12649
rect 1733 12207 3783 12597
rect 1733 12155 1760 12207
rect 1812 12155 1868 12207
rect 1920 12155 1976 12207
rect 2028 12155 2084 12207
rect 2136 12155 2192 12207
rect 2244 12155 2300 12207
rect 2352 12155 2408 12207
rect 2460 12155 2516 12207
rect 2568 12155 2624 12207
rect 2676 12155 2732 12207
rect 2784 12155 2840 12207
rect 2892 12155 2948 12207
rect 3000 12155 3056 12207
rect 3108 12155 3164 12207
rect 3216 12155 3272 12207
rect 3324 12155 3380 12207
rect 3432 12155 3488 12207
rect 3540 12155 3596 12207
rect 3648 12155 3704 12207
rect 3756 12155 3783 12207
rect 1733 11719 3783 12155
rect 1733 11667 1760 11719
rect 1812 11667 1868 11719
rect 1920 11667 1976 11719
rect 2028 11667 2084 11719
rect 2136 11667 2192 11719
rect 2244 11667 2300 11719
rect 2352 11667 2408 11719
rect 2460 11667 2516 11719
rect 2568 11667 2624 11719
rect 2676 11667 2732 11719
rect 2784 11667 2840 11719
rect 2892 11667 2948 11719
rect 3000 11667 3056 11719
rect 3108 11667 3164 11719
rect 3216 11667 3272 11719
rect 3324 11667 3380 11719
rect 3432 11667 3488 11719
rect 3540 11667 3596 11719
rect 3648 11667 3704 11719
rect 3756 11667 3783 11719
rect 1733 11231 3783 11667
rect 1733 11179 1760 11231
rect 1812 11179 1868 11231
rect 1920 11179 1976 11231
rect 2028 11179 2084 11231
rect 2136 11179 2192 11231
rect 2244 11179 2300 11231
rect 2352 11179 2408 11231
rect 2460 11179 2516 11231
rect 2568 11179 2624 11231
rect 2676 11179 2732 11231
rect 2784 11179 2840 11231
rect 2892 11179 2948 11231
rect 3000 11179 3056 11231
rect 3108 11179 3164 11231
rect 3216 11179 3272 11231
rect 3324 11179 3380 11231
rect 3432 11179 3488 11231
rect 3540 11179 3596 11231
rect 3648 11179 3704 11231
rect 3756 11179 3783 11231
rect 1733 10743 3783 11179
rect 1733 10691 1760 10743
rect 1812 10691 1868 10743
rect 1920 10691 1976 10743
rect 2028 10691 2084 10743
rect 2136 10691 2192 10743
rect 2244 10691 2300 10743
rect 2352 10691 2408 10743
rect 2460 10691 2516 10743
rect 2568 10691 2624 10743
rect 2676 10691 2732 10743
rect 2784 10691 2840 10743
rect 2892 10691 2948 10743
rect 3000 10691 3056 10743
rect 3108 10691 3164 10743
rect 3216 10691 3272 10743
rect 3324 10691 3380 10743
rect 3432 10691 3488 10743
rect 3540 10691 3596 10743
rect 3648 10691 3704 10743
rect 3756 10691 3783 10743
rect 1733 10255 3783 10691
rect 1733 10203 1760 10255
rect 1812 10203 1868 10255
rect 1920 10203 1976 10255
rect 2028 10203 2084 10255
rect 2136 10203 2192 10255
rect 2244 10203 2300 10255
rect 2352 10203 2408 10255
rect 2460 10203 2516 10255
rect 2568 10203 2624 10255
rect 2676 10203 2732 10255
rect 2784 10203 2840 10255
rect 2892 10203 2948 10255
rect 3000 10203 3056 10255
rect 3108 10203 3164 10255
rect 3216 10203 3272 10255
rect 3324 10203 3380 10255
rect 3432 10203 3488 10255
rect 3540 10203 3596 10255
rect 3648 10203 3704 10255
rect 3756 10203 3783 10255
rect 1733 9767 3783 10203
rect 1733 9715 1760 9767
rect 1812 9715 1868 9767
rect 1920 9715 1976 9767
rect 2028 9715 2084 9767
rect 2136 9715 2192 9767
rect 2244 9715 2300 9767
rect 2352 9715 2408 9767
rect 2460 9715 2516 9767
rect 2568 9715 2624 9767
rect 2676 9715 2732 9767
rect 2784 9715 2840 9767
rect 2892 9715 2948 9767
rect 3000 9715 3056 9767
rect 3108 9715 3164 9767
rect 3216 9715 3272 9767
rect 3324 9715 3380 9767
rect 3432 9715 3488 9767
rect 3540 9715 3596 9767
rect 3648 9715 3704 9767
rect 3756 9715 3783 9767
rect 1733 9279 3783 9715
rect 1733 9227 1760 9279
rect 1812 9227 1868 9279
rect 1920 9227 1976 9279
rect 2028 9227 2084 9279
rect 2136 9227 2192 9279
rect 2244 9227 2300 9279
rect 2352 9227 2408 9279
rect 2460 9227 2516 9279
rect 2568 9227 2624 9279
rect 2676 9227 2732 9279
rect 2784 9227 2840 9279
rect 2892 9227 2948 9279
rect 3000 9227 3056 9279
rect 3108 9227 3164 9279
rect 3216 9227 3272 9279
rect 3324 9227 3380 9279
rect 3432 9227 3488 9279
rect 3540 9227 3596 9279
rect 3648 9227 3704 9279
rect 3756 9227 3783 9279
rect 1733 8791 3783 9227
rect 1733 8739 1760 8791
rect 1812 8739 1868 8791
rect 1920 8739 1976 8791
rect 2028 8739 2084 8791
rect 2136 8739 2192 8791
rect 2244 8739 2300 8791
rect 2352 8739 2408 8791
rect 2460 8739 2516 8791
rect 2568 8739 2624 8791
rect 2676 8739 2732 8791
rect 2784 8739 2840 8791
rect 2892 8739 2948 8791
rect 3000 8739 3056 8791
rect 3108 8739 3164 8791
rect 3216 8739 3272 8791
rect 3324 8739 3380 8791
rect 3432 8739 3488 8791
rect 3540 8739 3596 8791
rect 3648 8739 3704 8791
rect 3756 8739 3783 8791
rect 1733 8303 3783 8739
rect 1733 8251 1760 8303
rect 1812 8251 1868 8303
rect 1920 8251 1976 8303
rect 2028 8251 2084 8303
rect 2136 8251 2192 8303
rect 2244 8251 2300 8303
rect 2352 8251 2408 8303
rect 2460 8251 2516 8303
rect 2568 8251 2624 8303
rect 2676 8251 2732 8303
rect 2784 8251 2840 8303
rect 2892 8251 2948 8303
rect 3000 8251 3056 8303
rect 3108 8251 3164 8303
rect 3216 8251 3272 8303
rect 3324 8251 3380 8303
rect 3432 8251 3488 8303
rect 3540 8251 3596 8303
rect 3648 8251 3704 8303
rect 3756 8251 3783 8303
rect 1733 7815 3783 8251
rect 1733 7763 1760 7815
rect 1812 7763 1868 7815
rect 1920 7763 1976 7815
rect 2028 7763 2084 7815
rect 2136 7763 2192 7815
rect 2244 7763 2300 7815
rect 2352 7763 2408 7815
rect 2460 7763 2516 7815
rect 2568 7763 2624 7815
rect 2676 7763 2732 7815
rect 2784 7763 2840 7815
rect 2892 7763 2948 7815
rect 3000 7763 3056 7815
rect 3108 7763 3164 7815
rect 3216 7763 3272 7815
rect 3324 7763 3380 7815
rect 3432 7763 3488 7815
rect 3540 7763 3596 7815
rect 3648 7763 3704 7815
rect 3756 7763 3783 7815
rect 1733 7327 3783 7763
rect 1733 7275 1760 7327
rect 1812 7275 1868 7327
rect 1920 7275 1976 7327
rect 2028 7275 2084 7327
rect 2136 7275 2192 7327
rect 2244 7275 2300 7327
rect 2352 7275 2408 7327
rect 2460 7275 2516 7327
rect 2568 7275 2624 7327
rect 2676 7275 2732 7327
rect 2784 7275 2840 7327
rect 2892 7275 2948 7327
rect 3000 7275 3056 7327
rect 3108 7275 3164 7327
rect 3216 7275 3272 7327
rect 3324 7275 3380 7327
rect 3432 7275 3488 7327
rect 3540 7275 3596 7327
rect 3648 7275 3704 7327
rect 3756 7275 3783 7327
rect 1733 6885 3783 7275
rect 1733 6833 1760 6885
rect 1812 6833 1868 6885
rect 1920 6833 1976 6885
rect 2028 6833 2084 6885
rect 2136 6833 2192 6885
rect 2244 6833 2300 6885
rect 2352 6833 2408 6885
rect 2460 6833 2516 6885
rect 2568 6833 2624 6885
rect 2676 6833 2732 6885
rect 2784 6833 2840 6885
rect 2892 6833 2948 6885
rect 3000 6833 3056 6885
rect 3108 6833 3164 6885
rect 3216 6833 3272 6885
rect 3324 6833 3380 6885
rect 3432 6833 3488 6885
rect 3540 6833 3596 6885
rect 3648 6833 3704 6885
rect 3756 6833 3783 6885
rect 1733 6777 3783 6833
rect 1733 6725 1760 6777
rect 1812 6725 1868 6777
rect 1920 6725 1976 6777
rect 2028 6725 2084 6777
rect 2136 6725 2192 6777
rect 2244 6725 2300 6777
rect 2352 6725 2408 6777
rect 2460 6725 2516 6777
rect 2568 6725 2624 6777
rect 2676 6725 2732 6777
rect 2784 6725 2840 6777
rect 2892 6725 2948 6777
rect 3000 6725 3056 6777
rect 3108 6725 3164 6777
rect 3216 6725 3272 6777
rect 3324 6725 3380 6777
rect 3432 6725 3488 6777
rect 3540 6725 3596 6777
rect 3648 6725 3704 6777
rect 3756 6725 3783 6777
rect 1733 6335 3783 6725
rect 1733 6283 1760 6335
rect 1812 6283 1868 6335
rect 1920 6283 1976 6335
rect 2028 6283 2084 6335
rect 2136 6283 2192 6335
rect 2244 6283 2300 6335
rect 2352 6283 2408 6335
rect 2460 6283 2516 6335
rect 2568 6283 2624 6335
rect 2676 6283 2732 6335
rect 2784 6283 2840 6335
rect 2892 6283 2948 6335
rect 3000 6283 3056 6335
rect 3108 6283 3164 6335
rect 3216 6283 3272 6335
rect 3324 6283 3380 6335
rect 3432 6283 3488 6335
rect 3540 6283 3596 6335
rect 3648 6283 3704 6335
rect 3756 6283 3783 6335
rect 1733 5847 3783 6283
rect 1733 5795 1760 5847
rect 1812 5795 1868 5847
rect 1920 5795 1976 5847
rect 2028 5795 2084 5847
rect 2136 5795 2192 5847
rect 2244 5795 2300 5847
rect 2352 5795 2408 5847
rect 2460 5795 2516 5847
rect 2568 5795 2624 5847
rect 2676 5795 2732 5847
rect 2784 5795 2840 5847
rect 2892 5795 2948 5847
rect 3000 5795 3056 5847
rect 3108 5795 3164 5847
rect 3216 5795 3272 5847
rect 3324 5795 3380 5847
rect 3432 5795 3488 5847
rect 3540 5795 3596 5847
rect 3648 5795 3704 5847
rect 3756 5795 3783 5847
rect 1733 5359 3783 5795
rect 1733 5307 1760 5359
rect 1812 5307 1868 5359
rect 1920 5307 1976 5359
rect 2028 5307 2084 5359
rect 2136 5307 2192 5359
rect 2244 5307 2300 5359
rect 2352 5307 2408 5359
rect 2460 5307 2516 5359
rect 2568 5307 2624 5359
rect 2676 5307 2732 5359
rect 2784 5307 2840 5359
rect 2892 5307 2948 5359
rect 3000 5307 3056 5359
rect 3108 5307 3164 5359
rect 3216 5307 3272 5359
rect 3324 5307 3380 5359
rect 3432 5307 3488 5359
rect 3540 5307 3596 5359
rect 3648 5307 3704 5359
rect 3756 5307 3783 5359
rect 1733 4871 3783 5307
rect 1733 4819 1760 4871
rect 1812 4819 1868 4871
rect 1920 4819 1976 4871
rect 2028 4819 2084 4871
rect 2136 4819 2192 4871
rect 2244 4819 2300 4871
rect 2352 4819 2408 4871
rect 2460 4819 2516 4871
rect 2568 4819 2624 4871
rect 2676 4819 2732 4871
rect 2784 4819 2840 4871
rect 2892 4819 2948 4871
rect 3000 4819 3056 4871
rect 3108 4819 3164 4871
rect 3216 4819 3272 4871
rect 3324 4819 3380 4871
rect 3432 4819 3488 4871
rect 3540 4819 3596 4871
rect 3648 4819 3704 4871
rect 3756 4819 3783 4871
rect 1733 4383 3783 4819
rect 1733 4331 1760 4383
rect 1812 4331 1868 4383
rect 1920 4331 1976 4383
rect 2028 4331 2084 4383
rect 2136 4331 2192 4383
rect 2244 4331 2300 4383
rect 2352 4331 2408 4383
rect 2460 4331 2516 4383
rect 2568 4331 2624 4383
rect 2676 4331 2732 4383
rect 2784 4331 2840 4383
rect 2892 4331 2948 4383
rect 3000 4331 3056 4383
rect 3108 4331 3164 4383
rect 3216 4331 3272 4383
rect 3324 4331 3380 4383
rect 3432 4331 3488 4383
rect 3540 4331 3596 4383
rect 3648 4331 3704 4383
rect 3756 4331 3783 4383
rect 1733 3895 3783 4331
rect 1733 3843 1760 3895
rect 1812 3843 1868 3895
rect 1920 3843 1976 3895
rect 2028 3843 2084 3895
rect 2136 3843 2192 3895
rect 2244 3843 2300 3895
rect 2352 3843 2408 3895
rect 2460 3843 2516 3895
rect 2568 3843 2624 3895
rect 2676 3843 2732 3895
rect 2784 3843 2840 3895
rect 2892 3843 2948 3895
rect 3000 3843 3056 3895
rect 3108 3843 3164 3895
rect 3216 3843 3272 3895
rect 3324 3843 3380 3895
rect 3432 3843 3488 3895
rect 3540 3843 3596 3895
rect 3648 3843 3704 3895
rect 3756 3843 3783 3895
rect 1733 3407 3783 3843
rect 1733 3355 1760 3407
rect 1812 3355 1868 3407
rect 1920 3355 1976 3407
rect 2028 3355 2084 3407
rect 2136 3355 2192 3407
rect 2244 3355 2300 3407
rect 2352 3355 2408 3407
rect 2460 3355 2516 3407
rect 2568 3355 2624 3407
rect 2676 3355 2732 3407
rect 2784 3355 2840 3407
rect 2892 3355 2948 3407
rect 3000 3355 3056 3407
rect 3108 3355 3164 3407
rect 3216 3355 3272 3407
rect 3324 3355 3380 3407
rect 3432 3355 3488 3407
rect 3540 3355 3596 3407
rect 3648 3355 3704 3407
rect 3756 3355 3783 3407
rect 1733 2919 3783 3355
rect 1733 2867 1760 2919
rect 1812 2867 1868 2919
rect 1920 2867 1976 2919
rect 2028 2867 2084 2919
rect 2136 2867 2192 2919
rect 2244 2867 2300 2919
rect 2352 2867 2408 2919
rect 2460 2867 2516 2919
rect 2568 2867 2624 2919
rect 2676 2867 2732 2919
rect 2784 2867 2840 2919
rect 2892 2867 2948 2919
rect 3000 2867 3056 2919
rect 3108 2867 3164 2919
rect 3216 2867 3272 2919
rect 3324 2867 3380 2919
rect 3432 2867 3488 2919
rect 3540 2867 3596 2919
rect 3648 2867 3704 2919
rect 3756 2867 3783 2919
rect 1733 2431 3783 2867
rect 1733 2379 1760 2431
rect 1812 2379 1868 2431
rect 1920 2379 1976 2431
rect 2028 2379 2084 2431
rect 2136 2379 2192 2431
rect 2244 2379 2300 2431
rect 2352 2379 2408 2431
rect 2460 2379 2516 2431
rect 2568 2379 2624 2431
rect 2676 2379 2732 2431
rect 2784 2379 2840 2431
rect 2892 2379 2948 2431
rect 3000 2379 3056 2431
rect 3108 2379 3164 2431
rect 3216 2379 3272 2431
rect 3324 2379 3380 2431
rect 3432 2379 3488 2431
rect 3540 2379 3596 2431
rect 3648 2379 3704 2431
rect 3756 2379 3783 2431
rect 1733 1943 3783 2379
rect 1733 1891 1760 1943
rect 1812 1891 1868 1943
rect 1920 1891 1976 1943
rect 2028 1891 2084 1943
rect 2136 1891 2192 1943
rect 2244 1891 2300 1943
rect 2352 1891 2408 1943
rect 2460 1891 2516 1943
rect 2568 1891 2624 1943
rect 2676 1891 2732 1943
rect 2784 1891 2840 1943
rect 2892 1891 2948 1943
rect 3000 1891 3056 1943
rect 3108 1891 3164 1943
rect 3216 1891 3272 1943
rect 3324 1891 3380 1943
rect 3432 1891 3488 1943
rect 3540 1891 3596 1943
rect 3648 1891 3704 1943
rect 3756 1891 3783 1943
rect 1733 1455 3783 1891
rect 1733 1403 1760 1455
rect 1812 1403 1868 1455
rect 1920 1403 1976 1455
rect 2028 1403 2084 1455
rect 2136 1403 2192 1455
rect 2244 1403 2300 1455
rect 2352 1403 2408 1455
rect 2460 1403 2516 1455
rect 2568 1403 2624 1455
rect 2676 1403 2732 1455
rect 2784 1403 2840 1455
rect 2892 1403 2948 1455
rect 3000 1403 3056 1455
rect 3108 1403 3164 1455
rect 3216 1403 3272 1455
rect 3324 1403 3380 1455
rect 3432 1403 3488 1455
rect 3540 1403 3596 1455
rect 3648 1403 3704 1455
rect 3756 1403 3783 1455
rect 1733 961 3783 1403
rect 1733 909 1760 961
rect 1812 909 1868 961
rect 1920 909 1976 961
rect 2028 909 2084 961
rect 2136 909 2192 961
rect 2244 909 2300 961
rect 2352 909 2408 961
rect 2460 909 2516 961
rect 2568 909 2624 961
rect 2676 909 2732 961
rect 2784 909 2840 961
rect 2892 909 2948 961
rect 3000 909 3056 961
rect 3108 909 3164 961
rect 3216 909 3272 961
rect 3324 909 3380 961
rect 3432 909 3488 961
rect 3540 909 3596 961
rect 3648 909 3704 961
rect 3756 909 3783 961
rect 1733 853 3783 909
rect 1733 801 1760 853
rect 1812 801 1868 853
rect 1920 801 1976 853
rect 2028 801 2084 853
rect 2136 801 2192 853
rect 2244 801 2300 853
rect 2352 801 2408 853
rect 2460 801 2516 853
rect 2568 801 2624 853
rect 2676 801 2732 853
rect 2784 801 2840 853
rect 2892 801 2948 853
rect 3000 801 3056 853
rect 3108 801 3164 853
rect 3216 801 3272 853
rect 3324 801 3380 853
rect 3432 801 3488 853
rect 3540 801 3596 853
rect 3648 801 3704 853
rect 3756 801 3783 853
rect 1733 745 3783 801
rect 1733 693 1760 745
rect 1812 693 1868 745
rect 1920 693 1976 745
rect 2028 693 2084 745
rect 2136 693 2192 745
rect 2244 693 2300 745
rect 2352 693 2408 745
rect 2460 693 2516 745
rect 2568 693 2624 745
rect 2676 693 2732 745
rect 2784 693 2840 745
rect 2892 693 2948 745
rect 3000 693 3056 745
rect 3108 693 3164 745
rect 3216 693 3272 745
rect 3324 693 3380 745
rect 3432 693 3488 745
rect 3540 693 3596 745
rect 3648 693 3704 745
rect 3756 693 3783 745
rect 1733 43 3783 693
rect 3843 25261 4043 25617
rect 3843 25209 3863 25261
rect 3915 25209 3971 25261
rect 4023 25209 4043 25261
rect 3843 25153 4043 25209
rect 3843 25101 3863 25153
rect 3915 25101 3971 25153
rect 4023 25101 4043 25153
rect 3843 25045 4043 25101
rect 3843 24993 3863 25045
rect 3915 24993 3971 25045
rect 4023 24993 4043 25045
rect 3843 23707 4043 24993
rect 3843 23655 3863 23707
rect 3915 23655 3971 23707
rect 4023 23655 4043 23707
rect 3843 23219 4043 23655
rect 3843 23167 3863 23219
rect 3915 23167 3971 23219
rect 4023 23167 4043 23219
rect 3843 22731 4043 23167
rect 3843 22679 3863 22731
rect 3915 22679 3971 22731
rect 4023 22679 4043 22731
rect 3843 22243 4043 22679
rect 3843 22191 3863 22243
rect 3915 22191 3971 22243
rect 4023 22191 4043 22243
rect 3843 21755 4043 22191
rect 3843 21703 3863 21755
rect 3915 21703 3971 21755
rect 4023 21703 4043 21755
rect 3843 21267 4043 21703
rect 3843 21215 3863 21267
rect 3915 21215 3971 21267
rect 4023 21215 4043 21267
rect 3843 20779 4043 21215
rect 3843 20727 3863 20779
rect 3915 20727 3971 20779
rect 4023 20727 4043 20779
rect 3843 20291 4043 20727
rect 3843 20239 3863 20291
rect 3915 20239 3971 20291
rect 4023 20239 4043 20291
rect 3843 19803 4043 20239
rect 3843 19751 3863 19803
rect 3915 19751 3971 19803
rect 4023 19751 4043 19803
rect 3843 19315 4043 19751
rect 3843 19263 3863 19315
rect 3915 19263 3971 19315
rect 4023 19263 4043 19315
rect 3843 17835 4043 19263
rect 3843 17783 3863 17835
rect 3915 17783 3971 17835
rect 4023 17783 4043 17835
rect 3843 17347 4043 17783
rect 3843 17295 3863 17347
rect 3915 17295 3971 17347
rect 4023 17295 4043 17347
rect 3843 16859 4043 17295
rect 3843 16807 3863 16859
rect 3915 16807 3971 16859
rect 4023 16807 4043 16859
rect 3843 16371 4043 16807
rect 3843 16319 3863 16371
rect 3915 16319 3971 16371
rect 4023 16319 4043 16371
rect 3843 15883 4043 16319
rect 3843 15831 3863 15883
rect 3915 15831 3971 15883
rect 4023 15831 4043 15883
rect 3843 15395 4043 15831
rect 3843 15343 3863 15395
rect 3915 15343 3971 15395
rect 4023 15343 4043 15395
rect 3843 14907 4043 15343
rect 3843 14855 3863 14907
rect 3915 14855 3971 14907
rect 4023 14855 4043 14907
rect 3843 14419 4043 14855
rect 3843 14367 3863 14419
rect 3915 14367 3971 14419
rect 4023 14367 4043 14419
rect 3843 13931 4043 14367
rect 3843 13879 3863 13931
rect 3915 13879 3971 13931
rect 4023 13879 4043 13931
rect 3843 13443 4043 13879
rect 3843 13391 3863 13443
rect 3915 13391 3971 13443
rect 4023 13391 4043 13443
rect 3843 11963 4043 13391
rect 3843 11911 3863 11963
rect 3915 11911 3971 11963
rect 4023 11911 4043 11963
rect 3843 11475 4043 11911
rect 3843 11423 3863 11475
rect 3915 11423 3971 11475
rect 4023 11423 4043 11475
rect 3843 10987 4043 11423
rect 3843 10935 3863 10987
rect 3915 10935 3971 10987
rect 4023 10935 4043 10987
rect 3843 10499 4043 10935
rect 3843 10447 3863 10499
rect 3915 10447 3971 10499
rect 4023 10447 4043 10499
rect 3843 10011 4043 10447
rect 3843 9959 3863 10011
rect 3915 9959 3971 10011
rect 4023 9959 4043 10011
rect 3843 9523 4043 9959
rect 3843 9471 3863 9523
rect 3915 9471 3971 9523
rect 4023 9471 4043 9523
rect 3843 9035 4043 9471
rect 3843 8983 3863 9035
rect 3915 8983 3971 9035
rect 4023 8983 4043 9035
rect 3843 8547 4043 8983
rect 3843 8495 3863 8547
rect 3915 8495 3971 8547
rect 4023 8495 4043 8547
rect 3843 8059 4043 8495
rect 3843 8007 3863 8059
rect 3915 8007 3971 8059
rect 4023 8007 4043 8059
rect 3843 7571 4043 8007
rect 3843 7519 3863 7571
rect 3915 7519 3971 7571
rect 4023 7519 4043 7571
rect 3843 6091 4043 7519
rect 3843 6039 3863 6091
rect 3915 6039 3971 6091
rect 4023 6039 4043 6091
rect 3843 5603 4043 6039
rect 3843 5551 3863 5603
rect 3915 5551 3971 5603
rect 4023 5551 4043 5603
rect 3843 5115 4043 5551
rect 3843 5063 3863 5115
rect 3915 5063 3971 5115
rect 4023 5063 4043 5115
rect 3843 4627 4043 5063
rect 3843 4575 3863 4627
rect 3915 4575 3971 4627
rect 4023 4575 4043 4627
rect 3843 4139 4043 4575
rect 3843 4087 3863 4139
rect 3915 4087 3971 4139
rect 4023 4087 4043 4139
rect 3843 3651 4043 4087
rect 3843 3599 3863 3651
rect 3915 3599 3971 3651
rect 4023 3599 4043 3651
rect 3843 3163 4043 3599
rect 3843 3111 3863 3163
rect 3915 3111 3971 3163
rect 4023 3111 4043 3163
rect 3843 2675 4043 3111
rect 3843 2623 3863 2675
rect 3915 2623 3971 2675
rect 4023 2623 4043 2675
rect 3843 2187 4043 2623
rect 3843 2135 3863 2187
rect 3915 2135 3971 2187
rect 4023 2135 4043 2187
rect 3843 1699 4043 2135
rect 3843 1647 3863 1699
rect 3915 1647 3971 1699
rect 4023 1647 4043 1699
rect 3843 361 4043 1647
rect 3843 309 3863 361
rect 3915 309 3971 361
rect 4023 309 4043 361
rect 3843 253 4043 309
rect 3843 201 3863 253
rect 3915 201 3971 253
rect 4023 201 4043 253
rect 3843 145 4043 201
rect 3843 93 3863 145
rect 3915 93 3971 145
rect 4023 93 4043 145
rect 3843 43 4043 93
rect 4103 24661 6153 25617
rect 4103 24609 4130 24661
rect 4182 24609 4238 24661
rect 4290 24609 4346 24661
rect 4398 24609 4454 24661
rect 4506 24609 4562 24661
rect 4614 24609 4670 24661
rect 4722 24609 4778 24661
rect 4830 24609 4886 24661
rect 4938 24609 4994 24661
rect 5046 24609 5102 24661
rect 5154 24609 5210 24661
rect 5262 24609 5318 24661
rect 5370 24609 5426 24661
rect 5478 24609 5534 24661
rect 5586 24609 5642 24661
rect 5694 24609 5750 24661
rect 5802 24609 5858 24661
rect 5910 24609 5966 24661
rect 6018 24609 6074 24661
rect 6126 24609 6153 24661
rect 4103 24553 6153 24609
rect 4103 24501 4130 24553
rect 4182 24501 4238 24553
rect 4290 24501 4346 24553
rect 4398 24501 4454 24553
rect 4506 24501 4562 24553
rect 4614 24501 4670 24553
rect 4722 24501 4778 24553
rect 4830 24501 4886 24553
rect 4938 24501 4994 24553
rect 5046 24501 5102 24553
rect 5154 24501 5210 24553
rect 5262 24501 5318 24553
rect 5370 24501 5426 24553
rect 5478 24501 5534 24553
rect 5586 24501 5642 24553
rect 5694 24501 5750 24553
rect 5802 24501 5858 24553
rect 5910 24501 5966 24553
rect 6018 24501 6074 24553
rect 6126 24501 6153 24553
rect 4103 24445 6153 24501
rect 4103 24393 4130 24445
rect 4182 24393 4238 24445
rect 4290 24393 4346 24445
rect 4398 24393 4454 24445
rect 4506 24393 4562 24445
rect 4614 24393 4670 24445
rect 4722 24393 4778 24445
rect 4830 24393 4886 24445
rect 4938 24393 4994 24445
rect 5046 24393 5102 24445
rect 5154 24393 5210 24445
rect 5262 24393 5318 24445
rect 5370 24393 5426 24445
rect 5478 24393 5534 24445
rect 5586 24393 5642 24445
rect 5694 24393 5750 24445
rect 5802 24393 5858 24445
rect 5910 24393 5966 24445
rect 6018 24393 6074 24445
rect 6126 24393 6153 24445
rect 4103 23951 6153 24393
rect 4103 23899 4130 23951
rect 4182 23899 4238 23951
rect 4290 23899 4346 23951
rect 4398 23899 4454 23951
rect 4506 23899 4562 23951
rect 4614 23899 4670 23951
rect 4722 23899 4778 23951
rect 4830 23899 4886 23951
rect 4938 23899 4994 23951
rect 5046 23899 5102 23951
rect 5154 23899 5210 23951
rect 5262 23899 5318 23951
rect 5370 23899 5426 23951
rect 5478 23899 5534 23951
rect 5586 23899 5642 23951
rect 5694 23899 5750 23951
rect 5802 23899 5858 23951
rect 5910 23899 5966 23951
rect 6018 23899 6074 23951
rect 6126 23899 6153 23951
rect 4103 23463 6153 23899
rect 4103 23411 4130 23463
rect 4182 23411 4238 23463
rect 4290 23411 4346 23463
rect 4398 23411 4454 23463
rect 4506 23411 4562 23463
rect 4614 23411 4670 23463
rect 4722 23411 4778 23463
rect 4830 23411 4886 23463
rect 4938 23411 4994 23463
rect 5046 23411 5102 23463
rect 5154 23411 5210 23463
rect 5262 23411 5318 23463
rect 5370 23411 5426 23463
rect 5478 23411 5534 23463
rect 5586 23411 5642 23463
rect 5694 23411 5750 23463
rect 5802 23411 5858 23463
rect 5910 23411 5966 23463
rect 6018 23411 6074 23463
rect 6126 23411 6153 23463
rect 4103 22975 6153 23411
rect 4103 22923 4130 22975
rect 4182 22923 4238 22975
rect 4290 22923 4346 22975
rect 4398 22923 4454 22975
rect 4506 22923 4562 22975
rect 4614 22923 4670 22975
rect 4722 22923 4778 22975
rect 4830 22923 4886 22975
rect 4938 22923 4994 22975
rect 5046 22923 5102 22975
rect 5154 22923 5210 22975
rect 5262 22923 5318 22975
rect 5370 22923 5426 22975
rect 5478 22923 5534 22975
rect 5586 22923 5642 22975
rect 5694 22923 5750 22975
rect 5802 22923 5858 22975
rect 5910 22923 5966 22975
rect 6018 22923 6074 22975
rect 6126 22923 6153 22975
rect 4103 22487 6153 22923
rect 4103 22435 4130 22487
rect 4182 22435 4238 22487
rect 4290 22435 4346 22487
rect 4398 22435 4454 22487
rect 4506 22435 4562 22487
rect 4614 22435 4670 22487
rect 4722 22435 4778 22487
rect 4830 22435 4886 22487
rect 4938 22435 4994 22487
rect 5046 22435 5102 22487
rect 5154 22435 5210 22487
rect 5262 22435 5318 22487
rect 5370 22435 5426 22487
rect 5478 22435 5534 22487
rect 5586 22435 5642 22487
rect 5694 22435 5750 22487
rect 5802 22435 5858 22487
rect 5910 22435 5966 22487
rect 6018 22435 6074 22487
rect 6126 22435 6153 22487
rect 4103 21999 6153 22435
rect 4103 21947 4130 21999
rect 4182 21947 4238 21999
rect 4290 21947 4346 21999
rect 4398 21947 4454 21999
rect 4506 21947 4562 21999
rect 4614 21947 4670 21999
rect 4722 21947 4778 21999
rect 4830 21947 4886 21999
rect 4938 21947 4994 21999
rect 5046 21947 5102 21999
rect 5154 21947 5210 21999
rect 5262 21947 5318 21999
rect 5370 21947 5426 21999
rect 5478 21947 5534 21999
rect 5586 21947 5642 21999
rect 5694 21947 5750 21999
rect 5802 21947 5858 21999
rect 5910 21947 5966 21999
rect 6018 21947 6074 21999
rect 6126 21947 6153 21999
rect 4103 21511 6153 21947
rect 4103 21459 4130 21511
rect 4182 21459 4238 21511
rect 4290 21459 4346 21511
rect 4398 21459 4454 21511
rect 4506 21459 4562 21511
rect 4614 21459 4670 21511
rect 4722 21459 4778 21511
rect 4830 21459 4886 21511
rect 4938 21459 4994 21511
rect 5046 21459 5102 21511
rect 5154 21459 5210 21511
rect 5262 21459 5318 21511
rect 5370 21459 5426 21511
rect 5478 21459 5534 21511
rect 5586 21459 5642 21511
rect 5694 21459 5750 21511
rect 5802 21459 5858 21511
rect 5910 21459 5966 21511
rect 6018 21459 6074 21511
rect 6126 21459 6153 21511
rect 4103 21023 6153 21459
rect 4103 20971 4130 21023
rect 4182 20971 4238 21023
rect 4290 20971 4346 21023
rect 4398 20971 4454 21023
rect 4506 20971 4562 21023
rect 4614 20971 4670 21023
rect 4722 20971 4778 21023
rect 4830 20971 4886 21023
rect 4938 20971 4994 21023
rect 5046 20971 5102 21023
rect 5154 20971 5210 21023
rect 5262 20971 5318 21023
rect 5370 20971 5426 21023
rect 5478 20971 5534 21023
rect 5586 20971 5642 21023
rect 5694 20971 5750 21023
rect 5802 20971 5858 21023
rect 5910 20971 5966 21023
rect 6018 20971 6074 21023
rect 6126 20971 6153 21023
rect 4103 20535 6153 20971
rect 4103 20483 4130 20535
rect 4182 20483 4238 20535
rect 4290 20483 4346 20535
rect 4398 20483 4454 20535
rect 4506 20483 4562 20535
rect 4614 20483 4670 20535
rect 4722 20483 4778 20535
rect 4830 20483 4886 20535
rect 4938 20483 4994 20535
rect 5046 20483 5102 20535
rect 5154 20483 5210 20535
rect 5262 20483 5318 20535
rect 5370 20483 5426 20535
rect 5478 20483 5534 20535
rect 5586 20483 5642 20535
rect 5694 20483 5750 20535
rect 5802 20483 5858 20535
rect 5910 20483 5966 20535
rect 6018 20483 6074 20535
rect 6126 20483 6153 20535
rect 4103 20047 6153 20483
rect 4103 19995 4130 20047
rect 4182 19995 4238 20047
rect 4290 19995 4346 20047
rect 4398 19995 4454 20047
rect 4506 19995 4562 20047
rect 4614 19995 4670 20047
rect 4722 19995 4778 20047
rect 4830 19995 4886 20047
rect 4938 19995 4994 20047
rect 5046 19995 5102 20047
rect 5154 19995 5210 20047
rect 5262 19995 5318 20047
rect 5370 19995 5426 20047
rect 5478 19995 5534 20047
rect 5586 19995 5642 20047
rect 5694 19995 5750 20047
rect 5802 19995 5858 20047
rect 5910 19995 5966 20047
rect 6018 19995 6074 20047
rect 6126 19995 6153 20047
rect 4103 19559 6153 19995
rect 4103 19507 4130 19559
rect 4182 19507 4238 19559
rect 4290 19507 4346 19559
rect 4398 19507 4454 19559
rect 4506 19507 4562 19559
rect 4614 19507 4670 19559
rect 4722 19507 4778 19559
rect 4830 19507 4886 19559
rect 4938 19507 4994 19559
rect 5046 19507 5102 19559
rect 5154 19507 5210 19559
rect 5262 19507 5318 19559
rect 5370 19507 5426 19559
rect 5478 19507 5534 19559
rect 5586 19507 5642 19559
rect 5694 19507 5750 19559
rect 5802 19507 5858 19559
rect 5910 19507 5966 19559
rect 6018 19507 6074 19559
rect 6126 19507 6153 19559
rect 4103 19071 6153 19507
rect 4103 19019 4130 19071
rect 4182 19019 4238 19071
rect 4290 19019 4346 19071
rect 4398 19019 4454 19071
rect 4506 19019 4562 19071
rect 4614 19019 4670 19071
rect 4722 19019 4778 19071
rect 4830 19019 4886 19071
rect 4938 19019 4994 19071
rect 5046 19019 5102 19071
rect 5154 19019 5210 19071
rect 5262 19019 5318 19071
rect 5370 19019 5426 19071
rect 5478 19019 5534 19071
rect 5586 19019 5642 19071
rect 5694 19019 5750 19071
rect 5802 19019 5858 19071
rect 5910 19019 5966 19071
rect 6018 19019 6074 19071
rect 6126 19019 6153 19071
rect 4103 18629 6153 19019
rect 4103 18577 4130 18629
rect 4182 18577 4238 18629
rect 4290 18577 4346 18629
rect 4398 18577 4454 18629
rect 4506 18577 4562 18629
rect 4614 18577 4670 18629
rect 4722 18577 4778 18629
rect 4830 18577 4886 18629
rect 4938 18577 4994 18629
rect 5046 18577 5102 18629
rect 5154 18577 5210 18629
rect 5262 18577 5318 18629
rect 5370 18577 5426 18629
rect 5478 18577 5534 18629
rect 5586 18577 5642 18629
rect 5694 18577 5750 18629
rect 5802 18577 5858 18629
rect 5910 18577 5966 18629
rect 6018 18577 6074 18629
rect 6126 18577 6153 18629
rect 4103 18521 6153 18577
rect 4103 18469 4130 18521
rect 4182 18469 4238 18521
rect 4290 18469 4346 18521
rect 4398 18469 4454 18521
rect 4506 18469 4562 18521
rect 4614 18469 4670 18521
rect 4722 18469 4778 18521
rect 4830 18469 4886 18521
rect 4938 18469 4994 18521
rect 5046 18469 5102 18521
rect 5154 18469 5210 18521
rect 5262 18469 5318 18521
rect 5370 18469 5426 18521
rect 5478 18469 5534 18521
rect 5586 18469 5642 18521
rect 5694 18469 5750 18521
rect 5802 18469 5858 18521
rect 5910 18469 5966 18521
rect 6018 18469 6074 18521
rect 6126 18469 6153 18521
rect 4103 18079 6153 18469
rect 4103 18027 4130 18079
rect 4182 18027 4238 18079
rect 4290 18027 4346 18079
rect 4398 18027 4454 18079
rect 4506 18027 4562 18079
rect 4614 18027 4670 18079
rect 4722 18027 4778 18079
rect 4830 18027 4886 18079
rect 4938 18027 4994 18079
rect 5046 18027 5102 18079
rect 5154 18027 5210 18079
rect 5262 18027 5318 18079
rect 5370 18027 5426 18079
rect 5478 18027 5534 18079
rect 5586 18027 5642 18079
rect 5694 18027 5750 18079
rect 5802 18027 5858 18079
rect 5910 18027 5966 18079
rect 6018 18027 6074 18079
rect 6126 18027 6153 18079
rect 4103 17591 6153 18027
rect 4103 17539 4130 17591
rect 4182 17539 4238 17591
rect 4290 17539 4346 17591
rect 4398 17539 4454 17591
rect 4506 17539 4562 17591
rect 4614 17539 4670 17591
rect 4722 17539 4778 17591
rect 4830 17539 4886 17591
rect 4938 17539 4994 17591
rect 5046 17539 5102 17591
rect 5154 17539 5210 17591
rect 5262 17539 5318 17591
rect 5370 17539 5426 17591
rect 5478 17539 5534 17591
rect 5586 17539 5642 17591
rect 5694 17539 5750 17591
rect 5802 17539 5858 17591
rect 5910 17539 5966 17591
rect 6018 17539 6074 17591
rect 6126 17539 6153 17591
rect 4103 17103 6153 17539
rect 4103 17051 4130 17103
rect 4182 17051 4238 17103
rect 4290 17051 4346 17103
rect 4398 17051 4454 17103
rect 4506 17051 4562 17103
rect 4614 17051 4670 17103
rect 4722 17051 4778 17103
rect 4830 17051 4886 17103
rect 4938 17051 4994 17103
rect 5046 17051 5102 17103
rect 5154 17051 5210 17103
rect 5262 17051 5318 17103
rect 5370 17051 5426 17103
rect 5478 17051 5534 17103
rect 5586 17051 5642 17103
rect 5694 17051 5750 17103
rect 5802 17051 5858 17103
rect 5910 17051 5966 17103
rect 6018 17051 6074 17103
rect 6126 17051 6153 17103
rect 4103 16615 6153 17051
rect 4103 16563 4130 16615
rect 4182 16563 4238 16615
rect 4290 16563 4346 16615
rect 4398 16563 4454 16615
rect 4506 16563 4562 16615
rect 4614 16563 4670 16615
rect 4722 16563 4778 16615
rect 4830 16563 4886 16615
rect 4938 16563 4994 16615
rect 5046 16563 5102 16615
rect 5154 16563 5210 16615
rect 5262 16563 5318 16615
rect 5370 16563 5426 16615
rect 5478 16563 5534 16615
rect 5586 16563 5642 16615
rect 5694 16563 5750 16615
rect 5802 16563 5858 16615
rect 5910 16563 5966 16615
rect 6018 16563 6074 16615
rect 6126 16563 6153 16615
rect 4103 16127 6153 16563
rect 4103 16075 4130 16127
rect 4182 16075 4238 16127
rect 4290 16075 4346 16127
rect 4398 16075 4454 16127
rect 4506 16075 4562 16127
rect 4614 16075 4670 16127
rect 4722 16075 4778 16127
rect 4830 16075 4886 16127
rect 4938 16075 4994 16127
rect 5046 16075 5102 16127
rect 5154 16075 5210 16127
rect 5262 16075 5318 16127
rect 5370 16075 5426 16127
rect 5478 16075 5534 16127
rect 5586 16075 5642 16127
rect 5694 16075 5750 16127
rect 5802 16075 5858 16127
rect 5910 16075 5966 16127
rect 6018 16075 6074 16127
rect 6126 16075 6153 16127
rect 4103 15639 6153 16075
rect 4103 15587 4130 15639
rect 4182 15587 4238 15639
rect 4290 15587 4346 15639
rect 4398 15587 4454 15639
rect 4506 15587 4562 15639
rect 4614 15587 4670 15639
rect 4722 15587 4778 15639
rect 4830 15587 4886 15639
rect 4938 15587 4994 15639
rect 5046 15587 5102 15639
rect 5154 15587 5210 15639
rect 5262 15587 5318 15639
rect 5370 15587 5426 15639
rect 5478 15587 5534 15639
rect 5586 15587 5642 15639
rect 5694 15587 5750 15639
rect 5802 15587 5858 15639
rect 5910 15587 5966 15639
rect 6018 15587 6074 15639
rect 6126 15587 6153 15639
rect 4103 15151 6153 15587
rect 4103 15099 4130 15151
rect 4182 15099 4238 15151
rect 4290 15099 4346 15151
rect 4398 15099 4454 15151
rect 4506 15099 4562 15151
rect 4614 15099 4670 15151
rect 4722 15099 4778 15151
rect 4830 15099 4886 15151
rect 4938 15099 4994 15151
rect 5046 15099 5102 15151
rect 5154 15099 5210 15151
rect 5262 15099 5318 15151
rect 5370 15099 5426 15151
rect 5478 15099 5534 15151
rect 5586 15099 5642 15151
rect 5694 15099 5750 15151
rect 5802 15099 5858 15151
rect 5910 15099 5966 15151
rect 6018 15099 6074 15151
rect 6126 15099 6153 15151
rect 4103 14663 6153 15099
rect 4103 14611 4130 14663
rect 4182 14611 4238 14663
rect 4290 14611 4346 14663
rect 4398 14611 4454 14663
rect 4506 14611 4562 14663
rect 4614 14611 4670 14663
rect 4722 14611 4778 14663
rect 4830 14611 4886 14663
rect 4938 14611 4994 14663
rect 5046 14611 5102 14663
rect 5154 14611 5210 14663
rect 5262 14611 5318 14663
rect 5370 14611 5426 14663
rect 5478 14611 5534 14663
rect 5586 14611 5642 14663
rect 5694 14611 5750 14663
rect 5802 14611 5858 14663
rect 5910 14611 5966 14663
rect 6018 14611 6074 14663
rect 6126 14611 6153 14663
rect 4103 14175 6153 14611
rect 4103 14123 4130 14175
rect 4182 14123 4238 14175
rect 4290 14123 4346 14175
rect 4398 14123 4454 14175
rect 4506 14123 4562 14175
rect 4614 14123 4670 14175
rect 4722 14123 4778 14175
rect 4830 14123 4886 14175
rect 4938 14123 4994 14175
rect 5046 14123 5102 14175
rect 5154 14123 5210 14175
rect 5262 14123 5318 14175
rect 5370 14123 5426 14175
rect 5478 14123 5534 14175
rect 5586 14123 5642 14175
rect 5694 14123 5750 14175
rect 5802 14123 5858 14175
rect 5910 14123 5966 14175
rect 6018 14123 6074 14175
rect 6126 14123 6153 14175
rect 4103 13687 6153 14123
rect 4103 13635 4130 13687
rect 4182 13635 4238 13687
rect 4290 13635 4346 13687
rect 4398 13635 4454 13687
rect 4506 13635 4562 13687
rect 4614 13635 4670 13687
rect 4722 13635 4778 13687
rect 4830 13635 4886 13687
rect 4938 13635 4994 13687
rect 5046 13635 5102 13687
rect 5154 13635 5210 13687
rect 5262 13635 5318 13687
rect 5370 13635 5426 13687
rect 5478 13635 5534 13687
rect 5586 13635 5642 13687
rect 5694 13635 5750 13687
rect 5802 13635 5858 13687
rect 5910 13635 5966 13687
rect 6018 13635 6074 13687
rect 6126 13635 6153 13687
rect 4103 13199 6153 13635
rect 4103 13147 4130 13199
rect 4182 13147 4238 13199
rect 4290 13147 4346 13199
rect 4398 13147 4454 13199
rect 4506 13147 4562 13199
rect 4614 13147 4670 13199
rect 4722 13147 4778 13199
rect 4830 13147 4886 13199
rect 4938 13147 4994 13199
rect 5046 13147 5102 13199
rect 5154 13147 5210 13199
rect 5262 13147 5318 13199
rect 5370 13147 5426 13199
rect 5478 13147 5534 13199
rect 5586 13147 5642 13199
rect 5694 13147 5750 13199
rect 5802 13147 5858 13199
rect 5910 13147 5966 13199
rect 6018 13147 6074 13199
rect 6126 13147 6153 13199
rect 4103 12757 6153 13147
rect 4103 12705 4130 12757
rect 4182 12705 4238 12757
rect 4290 12705 4346 12757
rect 4398 12705 4454 12757
rect 4506 12705 4562 12757
rect 4614 12705 4670 12757
rect 4722 12705 4778 12757
rect 4830 12705 4886 12757
rect 4938 12705 4994 12757
rect 5046 12705 5102 12757
rect 5154 12705 5210 12757
rect 5262 12705 5318 12757
rect 5370 12705 5426 12757
rect 5478 12705 5534 12757
rect 5586 12705 5642 12757
rect 5694 12705 5750 12757
rect 5802 12705 5858 12757
rect 5910 12705 5966 12757
rect 6018 12705 6074 12757
rect 6126 12705 6153 12757
rect 4103 12649 6153 12705
rect 4103 12597 4130 12649
rect 4182 12597 4238 12649
rect 4290 12597 4346 12649
rect 4398 12597 4454 12649
rect 4506 12597 4562 12649
rect 4614 12597 4670 12649
rect 4722 12597 4778 12649
rect 4830 12597 4886 12649
rect 4938 12597 4994 12649
rect 5046 12597 5102 12649
rect 5154 12597 5210 12649
rect 5262 12597 5318 12649
rect 5370 12597 5426 12649
rect 5478 12597 5534 12649
rect 5586 12597 5642 12649
rect 5694 12597 5750 12649
rect 5802 12597 5858 12649
rect 5910 12597 5966 12649
rect 6018 12597 6074 12649
rect 6126 12597 6153 12649
rect 4103 12207 6153 12597
rect 4103 12155 4130 12207
rect 4182 12155 4238 12207
rect 4290 12155 4346 12207
rect 4398 12155 4454 12207
rect 4506 12155 4562 12207
rect 4614 12155 4670 12207
rect 4722 12155 4778 12207
rect 4830 12155 4886 12207
rect 4938 12155 4994 12207
rect 5046 12155 5102 12207
rect 5154 12155 5210 12207
rect 5262 12155 5318 12207
rect 5370 12155 5426 12207
rect 5478 12155 5534 12207
rect 5586 12155 5642 12207
rect 5694 12155 5750 12207
rect 5802 12155 5858 12207
rect 5910 12155 5966 12207
rect 6018 12155 6074 12207
rect 6126 12155 6153 12207
rect 4103 11719 6153 12155
rect 4103 11667 4130 11719
rect 4182 11667 4238 11719
rect 4290 11667 4346 11719
rect 4398 11667 4454 11719
rect 4506 11667 4562 11719
rect 4614 11667 4670 11719
rect 4722 11667 4778 11719
rect 4830 11667 4886 11719
rect 4938 11667 4994 11719
rect 5046 11667 5102 11719
rect 5154 11667 5210 11719
rect 5262 11667 5318 11719
rect 5370 11667 5426 11719
rect 5478 11667 5534 11719
rect 5586 11667 5642 11719
rect 5694 11667 5750 11719
rect 5802 11667 5858 11719
rect 5910 11667 5966 11719
rect 6018 11667 6074 11719
rect 6126 11667 6153 11719
rect 4103 11231 6153 11667
rect 4103 11179 4130 11231
rect 4182 11179 4238 11231
rect 4290 11179 4346 11231
rect 4398 11179 4454 11231
rect 4506 11179 4562 11231
rect 4614 11179 4670 11231
rect 4722 11179 4778 11231
rect 4830 11179 4886 11231
rect 4938 11179 4994 11231
rect 5046 11179 5102 11231
rect 5154 11179 5210 11231
rect 5262 11179 5318 11231
rect 5370 11179 5426 11231
rect 5478 11179 5534 11231
rect 5586 11179 5642 11231
rect 5694 11179 5750 11231
rect 5802 11179 5858 11231
rect 5910 11179 5966 11231
rect 6018 11179 6074 11231
rect 6126 11179 6153 11231
rect 4103 10743 6153 11179
rect 4103 10691 4130 10743
rect 4182 10691 4238 10743
rect 4290 10691 4346 10743
rect 4398 10691 4454 10743
rect 4506 10691 4562 10743
rect 4614 10691 4670 10743
rect 4722 10691 4778 10743
rect 4830 10691 4886 10743
rect 4938 10691 4994 10743
rect 5046 10691 5102 10743
rect 5154 10691 5210 10743
rect 5262 10691 5318 10743
rect 5370 10691 5426 10743
rect 5478 10691 5534 10743
rect 5586 10691 5642 10743
rect 5694 10691 5750 10743
rect 5802 10691 5858 10743
rect 5910 10691 5966 10743
rect 6018 10691 6074 10743
rect 6126 10691 6153 10743
rect 4103 10255 6153 10691
rect 4103 10203 4130 10255
rect 4182 10203 4238 10255
rect 4290 10203 4346 10255
rect 4398 10203 4454 10255
rect 4506 10203 4562 10255
rect 4614 10203 4670 10255
rect 4722 10203 4778 10255
rect 4830 10203 4886 10255
rect 4938 10203 4994 10255
rect 5046 10203 5102 10255
rect 5154 10203 5210 10255
rect 5262 10203 5318 10255
rect 5370 10203 5426 10255
rect 5478 10203 5534 10255
rect 5586 10203 5642 10255
rect 5694 10203 5750 10255
rect 5802 10203 5858 10255
rect 5910 10203 5966 10255
rect 6018 10203 6074 10255
rect 6126 10203 6153 10255
rect 4103 9767 6153 10203
rect 4103 9715 4130 9767
rect 4182 9715 4238 9767
rect 4290 9715 4346 9767
rect 4398 9715 4454 9767
rect 4506 9715 4562 9767
rect 4614 9715 4670 9767
rect 4722 9715 4778 9767
rect 4830 9715 4886 9767
rect 4938 9715 4994 9767
rect 5046 9715 5102 9767
rect 5154 9715 5210 9767
rect 5262 9715 5318 9767
rect 5370 9715 5426 9767
rect 5478 9715 5534 9767
rect 5586 9715 5642 9767
rect 5694 9715 5750 9767
rect 5802 9715 5858 9767
rect 5910 9715 5966 9767
rect 6018 9715 6074 9767
rect 6126 9715 6153 9767
rect 4103 9279 6153 9715
rect 4103 9227 4130 9279
rect 4182 9227 4238 9279
rect 4290 9227 4346 9279
rect 4398 9227 4454 9279
rect 4506 9227 4562 9279
rect 4614 9227 4670 9279
rect 4722 9227 4778 9279
rect 4830 9227 4886 9279
rect 4938 9227 4994 9279
rect 5046 9227 5102 9279
rect 5154 9227 5210 9279
rect 5262 9227 5318 9279
rect 5370 9227 5426 9279
rect 5478 9227 5534 9279
rect 5586 9227 5642 9279
rect 5694 9227 5750 9279
rect 5802 9227 5858 9279
rect 5910 9227 5966 9279
rect 6018 9227 6074 9279
rect 6126 9227 6153 9279
rect 4103 8791 6153 9227
rect 4103 8739 4130 8791
rect 4182 8739 4238 8791
rect 4290 8739 4346 8791
rect 4398 8739 4454 8791
rect 4506 8739 4562 8791
rect 4614 8739 4670 8791
rect 4722 8739 4778 8791
rect 4830 8739 4886 8791
rect 4938 8739 4994 8791
rect 5046 8739 5102 8791
rect 5154 8739 5210 8791
rect 5262 8739 5318 8791
rect 5370 8739 5426 8791
rect 5478 8739 5534 8791
rect 5586 8739 5642 8791
rect 5694 8739 5750 8791
rect 5802 8739 5858 8791
rect 5910 8739 5966 8791
rect 6018 8739 6074 8791
rect 6126 8739 6153 8791
rect 4103 8303 6153 8739
rect 4103 8251 4130 8303
rect 4182 8251 4238 8303
rect 4290 8251 4346 8303
rect 4398 8251 4454 8303
rect 4506 8251 4562 8303
rect 4614 8251 4670 8303
rect 4722 8251 4778 8303
rect 4830 8251 4886 8303
rect 4938 8251 4994 8303
rect 5046 8251 5102 8303
rect 5154 8251 5210 8303
rect 5262 8251 5318 8303
rect 5370 8251 5426 8303
rect 5478 8251 5534 8303
rect 5586 8251 5642 8303
rect 5694 8251 5750 8303
rect 5802 8251 5858 8303
rect 5910 8251 5966 8303
rect 6018 8251 6074 8303
rect 6126 8251 6153 8303
rect 4103 7815 6153 8251
rect 4103 7763 4130 7815
rect 4182 7763 4238 7815
rect 4290 7763 4346 7815
rect 4398 7763 4454 7815
rect 4506 7763 4562 7815
rect 4614 7763 4670 7815
rect 4722 7763 4778 7815
rect 4830 7763 4886 7815
rect 4938 7763 4994 7815
rect 5046 7763 5102 7815
rect 5154 7763 5210 7815
rect 5262 7763 5318 7815
rect 5370 7763 5426 7815
rect 5478 7763 5534 7815
rect 5586 7763 5642 7815
rect 5694 7763 5750 7815
rect 5802 7763 5858 7815
rect 5910 7763 5966 7815
rect 6018 7763 6074 7815
rect 6126 7763 6153 7815
rect 4103 7327 6153 7763
rect 4103 7275 4130 7327
rect 4182 7275 4238 7327
rect 4290 7275 4346 7327
rect 4398 7275 4454 7327
rect 4506 7275 4562 7327
rect 4614 7275 4670 7327
rect 4722 7275 4778 7327
rect 4830 7275 4886 7327
rect 4938 7275 4994 7327
rect 5046 7275 5102 7327
rect 5154 7275 5210 7327
rect 5262 7275 5318 7327
rect 5370 7275 5426 7327
rect 5478 7275 5534 7327
rect 5586 7275 5642 7327
rect 5694 7275 5750 7327
rect 5802 7275 5858 7327
rect 5910 7275 5966 7327
rect 6018 7275 6074 7327
rect 6126 7275 6153 7327
rect 4103 6885 6153 7275
rect 4103 6833 4130 6885
rect 4182 6833 4238 6885
rect 4290 6833 4346 6885
rect 4398 6833 4454 6885
rect 4506 6833 4562 6885
rect 4614 6833 4670 6885
rect 4722 6833 4778 6885
rect 4830 6833 4886 6885
rect 4938 6833 4994 6885
rect 5046 6833 5102 6885
rect 5154 6833 5210 6885
rect 5262 6833 5318 6885
rect 5370 6833 5426 6885
rect 5478 6833 5534 6885
rect 5586 6833 5642 6885
rect 5694 6833 5750 6885
rect 5802 6833 5858 6885
rect 5910 6833 5966 6885
rect 6018 6833 6074 6885
rect 6126 6833 6153 6885
rect 4103 6777 6153 6833
rect 4103 6725 4130 6777
rect 4182 6725 4238 6777
rect 4290 6725 4346 6777
rect 4398 6725 4454 6777
rect 4506 6725 4562 6777
rect 4614 6725 4670 6777
rect 4722 6725 4778 6777
rect 4830 6725 4886 6777
rect 4938 6725 4994 6777
rect 5046 6725 5102 6777
rect 5154 6725 5210 6777
rect 5262 6725 5318 6777
rect 5370 6725 5426 6777
rect 5478 6725 5534 6777
rect 5586 6725 5642 6777
rect 5694 6725 5750 6777
rect 5802 6725 5858 6777
rect 5910 6725 5966 6777
rect 6018 6725 6074 6777
rect 6126 6725 6153 6777
rect 4103 6335 6153 6725
rect 4103 6283 4130 6335
rect 4182 6283 4238 6335
rect 4290 6283 4346 6335
rect 4398 6283 4454 6335
rect 4506 6283 4562 6335
rect 4614 6283 4670 6335
rect 4722 6283 4778 6335
rect 4830 6283 4886 6335
rect 4938 6283 4994 6335
rect 5046 6283 5102 6335
rect 5154 6283 5210 6335
rect 5262 6283 5318 6335
rect 5370 6283 5426 6335
rect 5478 6283 5534 6335
rect 5586 6283 5642 6335
rect 5694 6283 5750 6335
rect 5802 6283 5858 6335
rect 5910 6283 5966 6335
rect 6018 6283 6074 6335
rect 6126 6283 6153 6335
rect 4103 5847 6153 6283
rect 4103 5795 4130 5847
rect 4182 5795 4238 5847
rect 4290 5795 4346 5847
rect 4398 5795 4454 5847
rect 4506 5795 4562 5847
rect 4614 5795 4670 5847
rect 4722 5795 4778 5847
rect 4830 5795 4886 5847
rect 4938 5795 4994 5847
rect 5046 5795 5102 5847
rect 5154 5795 5210 5847
rect 5262 5795 5318 5847
rect 5370 5795 5426 5847
rect 5478 5795 5534 5847
rect 5586 5795 5642 5847
rect 5694 5795 5750 5847
rect 5802 5795 5858 5847
rect 5910 5795 5966 5847
rect 6018 5795 6074 5847
rect 6126 5795 6153 5847
rect 4103 5359 6153 5795
rect 4103 5307 4130 5359
rect 4182 5307 4238 5359
rect 4290 5307 4346 5359
rect 4398 5307 4454 5359
rect 4506 5307 4562 5359
rect 4614 5307 4670 5359
rect 4722 5307 4778 5359
rect 4830 5307 4886 5359
rect 4938 5307 4994 5359
rect 5046 5307 5102 5359
rect 5154 5307 5210 5359
rect 5262 5307 5318 5359
rect 5370 5307 5426 5359
rect 5478 5307 5534 5359
rect 5586 5307 5642 5359
rect 5694 5307 5750 5359
rect 5802 5307 5858 5359
rect 5910 5307 5966 5359
rect 6018 5307 6074 5359
rect 6126 5307 6153 5359
rect 4103 4871 6153 5307
rect 4103 4819 4130 4871
rect 4182 4819 4238 4871
rect 4290 4819 4346 4871
rect 4398 4819 4454 4871
rect 4506 4819 4562 4871
rect 4614 4819 4670 4871
rect 4722 4819 4778 4871
rect 4830 4819 4886 4871
rect 4938 4819 4994 4871
rect 5046 4819 5102 4871
rect 5154 4819 5210 4871
rect 5262 4819 5318 4871
rect 5370 4819 5426 4871
rect 5478 4819 5534 4871
rect 5586 4819 5642 4871
rect 5694 4819 5750 4871
rect 5802 4819 5858 4871
rect 5910 4819 5966 4871
rect 6018 4819 6074 4871
rect 6126 4819 6153 4871
rect 4103 4383 6153 4819
rect 4103 4331 4130 4383
rect 4182 4331 4238 4383
rect 4290 4331 4346 4383
rect 4398 4331 4454 4383
rect 4506 4331 4562 4383
rect 4614 4331 4670 4383
rect 4722 4331 4778 4383
rect 4830 4331 4886 4383
rect 4938 4331 4994 4383
rect 5046 4331 5102 4383
rect 5154 4331 5210 4383
rect 5262 4331 5318 4383
rect 5370 4331 5426 4383
rect 5478 4331 5534 4383
rect 5586 4331 5642 4383
rect 5694 4331 5750 4383
rect 5802 4331 5858 4383
rect 5910 4331 5966 4383
rect 6018 4331 6074 4383
rect 6126 4331 6153 4383
rect 4103 3895 6153 4331
rect 4103 3843 4130 3895
rect 4182 3843 4238 3895
rect 4290 3843 4346 3895
rect 4398 3843 4454 3895
rect 4506 3843 4562 3895
rect 4614 3843 4670 3895
rect 4722 3843 4778 3895
rect 4830 3843 4886 3895
rect 4938 3843 4994 3895
rect 5046 3843 5102 3895
rect 5154 3843 5210 3895
rect 5262 3843 5318 3895
rect 5370 3843 5426 3895
rect 5478 3843 5534 3895
rect 5586 3843 5642 3895
rect 5694 3843 5750 3895
rect 5802 3843 5858 3895
rect 5910 3843 5966 3895
rect 6018 3843 6074 3895
rect 6126 3843 6153 3895
rect 4103 3407 6153 3843
rect 4103 3355 4130 3407
rect 4182 3355 4238 3407
rect 4290 3355 4346 3407
rect 4398 3355 4454 3407
rect 4506 3355 4562 3407
rect 4614 3355 4670 3407
rect 4722 3355 4778 3407
rect 4830 3355 4886 3407
rect 4938 3355 4994 3407
rect 5046 3355 5102 3407
rect 5154 3355 5210 3407
rect 5262 3355 5318 3407
rect 5370 3355 5426 3407
rect 5478 3355 5534 3407
rect 5586 3355 5642 3407
rect 5694 3355 5750 3407
rect 5802 3355 5858 3407
rect 5910 3355 5966 3407
rect 6018 3355 6074 3407
rect 6126 3355 6153 3407
rect 4103 2919 6153 3355
rect 4103 2867 4130 2919
rect 4182 2867 4238 2919
rect 4290 2867 4346 2919
rect 4398 2867 4454 2919
rect 4506 2867 4562 2919
rect 4614 2867 4670 2919
rect 4722 2867 4778 2919
rect 4830 2867 4886 2919
rect 4938 2867 4994 2919
rect 5046 2867 5102 2919
rect 5154 2867 5210 2919
rect 5262 2867 5318 2919
rect 5370 2867 5426 2919
rect 5478 2867 5534 2919
rect 5586 2867 5642 2919
rect 5694 2867 5750 2919
rect 5802 2867 5858 2919
rect 5910 2867 5966 2919
rect 6018 2867 6074 2919
rect 6126 2867 6153 2919
rect 4103 2431 6153 2867
rect 4103 2379 4130 2431
rect 4182 2379 4238 2431
rect 4290 2379 4346 2431
rect 4398 2379 4454 2431
rect 4506 2379 4562 2431
rect 4614 2379 4670 2431
rect 4722 2379 4778 2431
rect 4830 2379 4886 2431
rect 4938 2379 4994 2431
rect 5046 2379 5102 2431
rect 5154 2379 5210 2431
rect 5262 2379 5318 2431
rect 5370 2379 5426 2431
rect 5478 2379 5534 2431
rect 5586 2379 5642 2431
rect 5694 2379 5750 2431
rect 5802 2379 5858 2431
rect 5910 2379 5966 2431
rect 6018 2379 6074 2431
rect 6126 2379 6153 2431
rect 4103 1943 6153 2379
rect 4103 1891 4130 1943
rect 4182 1891 4238 1943
rect 4290 1891 4346 1943
rect 4398 1891 4454 1943
rect 4506 1891 4562 1943
rect 4614 1891 4670 1943
rect 4722 1891 4778 1943
rect 4830 1891 4886 1943
rect 4938 1891 4994 1943
rect 5046 1891 5102 1943
rect 5154 1891 5210 1943
rect 5262 1891 5318 1943
rect 5370 1891 5426 1943
rect 5478 1891 5534 1943
rect 5586 1891 5642 1943
rect 5694 1891 5750 1943
rect 5802 1891 5858 1943
rect 5910 1891 5966 1943
rect 6018 1891 6074 1943
rect 6126 1891 6153 1943
rect 4103 1455 6153 1891
rect 4103 1403 4130 1455
rect 4182 1403 4238 1455
rect 4290 1403 4346 1455
rect 4398 1403 4454 1455
rect 4506 1403 4562 1455
rect 4614 1403 4670 1455
rect 4722 1403 4778 1455
rect 4830 1403 4886 1455
rect 4938 1403 4994 1455
rect 5046 1403 5102 1455
rect 5154 1403 5210 1455
rect 5262 1403 5318 1455
rect 5370 1403 5426 1455
rect 5478 1403 5534 1455
rect 5586 1403 5642 1455
rect 5694 1403 5750 1455
rect 5802 1403 5858 1455
rect 5910 1403 5966 1455
rect 6018 1403 6074 1455
rect 6126 1403 6153 1455
rect 4103 961 6153 1403
rect 4103 909 4130 961
rect 4182 909 4238 961
rect 4290 909 4346 961
rect 4398 909 4454 961
rect 4506 909 4562 961
rect 4614 909 4670 961
rect 4722 909 4778 961
rect 4830 909 4886 961
rect 4938 909 4994 961
rect 5046 909 5102 961
rect 5154 909 5210 961
rect 5262 909 5318 961
rect 5370 909 5426 961
rect 5478 909 5534 961
rect 5586 909 5642 961
rect 5694 909 5750 961
rect 5802 909 5858 961
rect 5910 909 5966 961
rect 6018 909 6074 961
rect 6126 909 6153 961
rect 4103 853 6153 909
rect 4103 801 4130 853
rect 4182 801 4238 853
rect 4290 801 4346 853
rect 4398 801 4454 853
rect 4506 801 4562 853
rect 4614 801 4670 853
rect 4722 801 4778 853
rect 4830 801 4886 853
rect 4938 801 4994 853
rect 5046 801 5102 853
rect 5154 801 5210 853
rect 5262 801 5318 853
rect 5370 801 5426 853
rect 5478 801 5534 853
rect 5586 801 5642 853
rect 5694 801 5750 853
rect 5802 801 5858 853
rect 5910 801 5966 853
rect 6018 801 6074 853
rect 6126 801 6153 853
rect 4103 745 6153 801
rect 4103 693 4130 745
rect 4182 693 4238 745
rect 4290 693 4346 745
rect 4398 693 4454 745
rect 4506 693 4562 745
rect 4614 693 4670 745
rect 4722 693 4778 745
rect 4830 693 4886 745
rect 4938 693 4994 745
rect 5046 693 5102 745
rect 5154 693 5210 745
rect 5262 693 5318 745
rect 5370 693 5426 745
rect 5478 693 5534 745
rect 5586 693 5642 745
rect 5694 693 5750 745
rect 5802 693 5858 745
rect 5910 693 5966 745
rect 6018 693 6074 745
rect 6126 693 6153 745
rect 4103 43 6153 693
rect 6213 25261 6749 25617
rect 6213 25209 6239 25261
rect 6291 25209 6347 25261
rect 6399 25209 6455 25261
rect 6507 25209 6563 25261
rect 6615 25209 6671 25261
rect 6723 25209 6749 25261
rect 6213 25153 6749 25209
rect 6213 25101 6239 25153
rect 6291 25101 6347 25153
rect 6399 25101 6455 25153
rect 6507 25101 6563 25153
rect 6615 25101 6671 25153
rect 6723 25101 6749 25153
rect 6213 25045 6749 25101
rect 6213 24993 6239 25045
rect 6291 24993 6347 25045
rect 6399 24993 6455 25045
rect 6507 24993 6563 25045
rect 6615 24993 6671 25045
rect 6723 24993 6749 25045
rect 6213 23707 6749 24993
rect 6213 23655 6239 23707
rect 6291 23655 6347 23707
rect 6399 23655 6455 23707
rect 6507 23655 6563 23707
rect 6615 23655 6671 23707
rect 6723 23655 6749 23707
rect 6213 23219 6749 23655
rect 6213 23167 6239 23219
rect 6291 23167 6347 23219
rect 6399 23167 6455 23219
rect 6507 23167 6563 23219
rect 6615 23167 6671 23219
rect 6723 23167 6749 23219
rect 6213 22731 6749 23167
rect 6213 22679 6239 22731
rect 6291 22679 6347 22731
rect 6399 22679 6455 22731
rect 6507 22679 6563 22731
rect 6615 22679 6671 22731
rect 6723 22679 6749 22731
rect 6213 22243 6749 22679
rect 6213 22191 6239 22243
rect 6291 22191 6347 22243
rect 6399 22191 6455 22243
rect 6507 22191 6563 22243
rect 6615 22191 6671 22243
rect 6723 22191 6749 22243
rect 6213 21755 6749 22191
rect 6213 21703 6239 21755
rect 6291 21703 6347 21755
rect 6399 21703 6455 21755
rect 6507 21703 6563 21755
rect 6615 21703 6671 21755
rect 6723 21703 6749 21755
rect 6213 21267 6749 21703
rect 6213 21215 6239 21267
rect 6291 21215 6347 21267
rect 6399 21215 6455 21267
rect 6507 21215 6563 21267
rect 6615 21215 6671 21267
rect 6723 21215 6749 21267
rect 6213 20779 6749 21215
rect 6213 20727 6239 20779
rect 6291 20727 6347 20779
rect 6399 20727 6455 20779
rect 6507 20727 6563 20779
rect 6615 20727 6671 20779
rect 6723 20727 6749 20779
rect 6213 20291 6749 20727
rect 6213 20239 6239 20291
rect 6291 20239 6347 20291
rect 6399 20239 6455 20291
rect 6507 20239 6563 20291
rect 6615 20239 6671 20291
rect 6723 20239 6749 20291
rect 6213 19803 6749 20239
rect 6213 19751 6239 19803
rect 6291 19751 6347 19803
rect 6399 19751 6455 19803
rect 6507 19751 6563 19803
rect 6615 19751 6671 19803
rect 6723 19751 6749 19803
rect 6213 19315 6749 19751
rect 6213 19263 6239 19315
rect 6291 19263 6347 19315
rect 6399 19263 6455 19315
rect 6507 19263 6563 19315
rect 6615 19263 6671 19315
rect 6723 19263 6749 19315
rect 6213 17835 6749 19263
rect 6213 17783 6239 17835
rect 6291 17783 6347 17835
rect 6399 17783 6455 17835
rect 6507 17783 6563 17835
rect 6615 17783 6671 17835
rect 6723 17783 6749 17835
rect 6213 17347 6749 17783
rect 6213 17295 6239 17347
rect 6291 17295 6347 17347
rect 6399 17295 6455 17347
rect 6507 17295 6563 17347
rect 6615 17295 6671 17347
rect 6723 17295 6749 17347
rect 6213 16859 6749 17295
rect 6213 16807 6239 16859
rect 6291 16807 6347 16859
rect 6399 16807 6455 16859
rect 6507 16807 6563 16859
rect 6615 16807 6671 16859
rect 6723 16807 6749 16859
rect 6213 16371 6749 16807
rect 6213 16319 6239 16371
rect 6291 16319 6347 16371
rect 6399 16319 6455 16371
rect 6507 16319 6563 16371
rect 6615 16319 6671 16371
rect 6723 16319 6749 16371
rect 6213 15883 6749 16319
rect 6213 15831 6239 15883
rect 6291 15831 6347 15883
rect 6399 15831 6455 15883
rect 6507 15831 6563 15883
rect 6615 15831 6671 15883
rect 6723 15831 6749 15883
rect 6213 15395 6749 15831
rect 6213 15343 6239 15395
rect 6291 15343 6347 15395
rect 6399 15343 6455 15395
rect 6507 15343 6563 15395
rect 6615 15343 6671 15395
rect 6723 15343 6749 15395
rect 6213 14907 6749 15343
rect 6213 14855 6239 14907
rect 6291 14855 6347 14907
rect 6399 14855 6455 14907
rect 6507 14855 6563 14907
rect 6615 14855 6671 14907
rect 6723 14855 6749 14907
rect 6213 14419 6749 14855
rect 6213 14367 6239 14419
rect 6291 14367 6347 14419
rect 6399 14367 6455 14419
rect 6507 14367 6563 14419
rect 6615 14367 6671 14419
rect 6723 14367 6749 14419
rect 6213 13931 6749 14367
rect 6213 13879 6239 13931
rect 6291 13879 6347 13931
rect 6399 13879 6455 13931
rect 6507 13879 6563 13931
rect 6615 13879 6671 13931
rect 6723 13879 6749 13931
rect 6213 13443 6749 13879
rect 6213 13391 6239 13443
rect 6291 13391 6347 13443
rect 6399 13391 6455 13443
rect 6507 13391 6563 13443
rect 6615 13391 6671 13443
rect 6723 13391 6749 13443
rect 6213 11963 6749 13391
rect 6213 11911 6239 11963
rect 6291 11911 6347 11963
rect 6399 11911 6455 11963
rect 6507 11911 6563 11963
rect 6615 11911 6671 11963
rect 6723 11911 6749 11963
rect 6213 11475 6749 11911
rect 6213 11423 6239 11475
rect 6291 11423 6347 11475
rect 6399 11423 6455 11475
rect 6507 11423 6563 11475
rect 6615 11423 6671 11475
rect 6723 11423 6749 11475
rect 6213 10987 6749 11423
rect 6213 10935 6239 10987
rect 6291 10935 6347 10987
rect 6399 10935 6455 10987
rect 6507 10935 6563 10987
rect 6615 10935 6671 10987
rect 6723 10935 6749 10987
rect 6213 10499 6749 10935
rect 6213 10447 6239 10499
rect 6291 10447 6347 10499
rect 6399 10447 6455 10499
rect 6507 10447 6563 10499
rect 6615 10447 6671 10499
rect 6723 10447 6749 10499
rect 6213 10011 6749 10447
rect 6213 9959 6239 10011
rect 6291 9959 6347 10011
rect 6399 9959 6455 10011
rect 6507 9959 6563 10011
rect 6615 9959 6671 10011
rect 6723 9959 6749 10011
rect 6213 9523 6749 9959
rect 6213 9471 6239 9523
rect 6291 9471 6347 9523
rect 6399 9471 6455 9523
rect 6507 9471 6563 9523
rect 6615 9471 6671 9523
rect 6723 9471 6749 9523
rect 6213 9035 6749 9471
rect 6213 8983 6239 9035
rect 6291 8983 6347 9035
rect 6399 8983 6455 9035
rect 6507 8983 6563 9035
rect 6615 8983 6671 9035
rect 6723 8983 6749 9035
rect 6213 8547 6749 8983
rect 6213 8495 6239 8547
rect 6291 8495 6347 8547
rect 6399 8495 6455 8547
rect 6507 8495 6563 8547
rect 6615 8495 6671 8547
rect 6723 8495 6749 8547
rect 6213 8059 6749 8495
rect 6213 8007 6239 8059
rect 6291 8007 6347 8059
rect 6399 8007 6455 8059
rect 6507 8007 6563 8059
rect 6615 8007 6671 8059
rect 6723 8007 6749 8059
rect 6213 7571 6749 8007
rect 6213 7519 6239 7571
rect 6291 7519 6347 7571
rect 6399 7519 6455 7571
rect 6507 7519 6563 7571
rect 6615 7519 6671 7571
rect 6723 7519 6749 7571
rect 6213 6091 6749 7519
rect 6213 6039 6239 6091
rect 6291 6039 6347 6091
rect 6399 6039 6455 6091
rect 6507 6039 6563 6091
rect 6615 6039 6671 6091
rect 6723 6039 6749 6091
rect 6213 5603 6749 6039
rect 6213 5551 6239 5603
rect 6291 5551 6347 5603
rect 6399 5551 6455 5603
rect 6507 5551 6563 5603
rect 6615 5551 6671 5603
rect 6723 5551 6749 5603
rect 6213 5115 6749 5551
rect 6213 5063 6239 5115
rect 6291 5063 6347 5115
rect 6399 5063 6455 5115
rect 6507 5063 6563 5115
rect 6615 5063 6671 5115
rect 6723 5063 6749 5115
rect 6213 4627 6749 5063
rect 6213 4575 6239 4627
rect 6291 4575 6347 4627
rect 6399 4575 6455 4627
rect 6507 4575 6563 4627
rect 6615 4575 6671 4627
rect 6723 4575 6749 4627
rect 6213 4139 6749 4575
rect 6213 4087 6239 4139
rect 6291 4087 6347 4139
rect 6399 4087 6455 4139
rect 6507 4087 6563 4139
rect 6615 4087 6671 4139
rect 6723 4087 6749 4139
rect 6213 3651 6749 4087
rect 6213 3599 6239 3651
rect 6291 3599 6347 3651
rect 6399 3599 6455 3651
rect 6507 3599 6563 3651
rect 6615 3599 6671 3651
rect 6723 3599 6749 3651
rect 6213 3163 6749 3599
rect 6213 3111 6239 3163
rect 6291 3111 6347 3163
rect 6399 3111 6455 3163
rect 6507 3111 6563 3163
rect 6615 3111 6671 3163
rect 6723 3111 6749 3163
rect 6213 2675 6749 3111
rect 6213 2623 6239 2675
rect 6291 2623 6347 2675
rect 6399 2623 6455 2675
rect 6507 2623 6563 2675
rect 6615 2623 6671 2675
rect 6723 2623 6749 2675
rect 6213 2187 6749 2623
rect 6213 2135 6239 2187
rect 6291 2135 6347 2187
rect 6399 2135 6455 2187
rect 6507 2135 6563 2187
rect 6615 2135 6671 2187
rect 6723 2135 6749 2187
rect 6213 1699 6749 2135
rect 6213 1647 6239 1699
rect 6291 1647 6347 1699
rect 6399 1647 6455 1699
rect 6507 1647 6563 1699
rect 6615 1647 6671 1699
rect 6723 1647 6749 1699
rect 6213 361 6749 1647
rect 6213 309 6239 361
rect 6291 309 6347 361
rect 6399 309 6455 361
rect 6507 309 6563 361
rect 6615 309 6671 361
rect 6723 309 6749 361
rect 6213 253 6749 309
rect 6213 201 6239 253
rect 6291 201 6347 253
rect 6399 201 6455 253
rect 6507 201 6563 253
rect 6615 201 6671 253
rect 6723 201 6749 253
rect 6213 145 6749 201
rect 6213 93 6239 145
rect 6291 93 6347 145
rect 6399 93 6455 145
rect 6507 93 6563 145
rect 6615 93 6671 145
rect 6723 93 6749 145
rect 6213 43 6749 93
rect 6809 24661 8859 25617
rect 6809 24609 6836 24661
rect 6888 24609 6944 24661
rect 6996 24609 7052 24661
rect 7104 24609 7160 24661
rect 7212 24609 7268 24661
rect 7320 24609 7376 24661
rect 7428 24609 7484 24661
rect 7536 24609 7592 24661
rect 7644 24609 7700 24661
rect 7752 24609 7808 24661
rect 7860 24609 7916 24661
rect 7968 24609 8024 24661
rect 8076 24609 8132 24661
rect 8184 24609 8240 24661
rect 8292 24609 8348 24661
rect 8400 24609 8456 24661
rect 8508 24609 8564 24661
rect 8616 24609 8672 24661
rect 8724 24609 8780 24661
rect 8832 24609 8859 24661
rect 6809 24553 8859 24609
rect 6809 24501 6836 24553
rect 6888 24501 6944 24553
rect 6996 24501 7052 24553
rect 7104 24501 7160 24553
rect 7212 24501 7268 24553
rect 7320 24501 7376 24553
rect 7428 24501 7484 24553
rect 7536 24501 7592 24553
rect 7644 24501 7700 24553
rect 7752 24501 7808 24553
rect 7860 24501 7916 24553
rect 7968 24501 8024 24553
rect 8076 24501 8132 24553
rect 8184 24501 8240 24553
rect 8292 24501 8348 24553
rect 8400 24501 8456 24553
rect 8508 24501 8564 24553
rect 8616 24501 8672 24553
rect 8724 24501 8780 24553
rect 8832 24501 8859 24553
rect 6809 24445 8859 24501
rect 6809 24393 6836 24445
rect 6888 24393 6944 24445
rect 6996 24393 7052 24445
rect 7104 24393 7160 24445
rect 7212 24393 7268 24445
rect 7320 24393 7376 24445
rect 7428 24393 7484 24445
rect 7536 24393 7592 24445
rect 7644 24393 7700 24445
rect 7752 24393 7808 24445
rect 7860 24393 7916 24445
rect 7968 24393 8024 24445
rect 8076 24393 8132 24445
rect 8184 24393 8240 24445
rect 8292 24393 8348 24445
rect 8400 24393 8456 24445
rect 8508 24393 8564 24445
rect 8616 24393 8672 24445
rect 8724 24393 8780 24445
rect 8832 24393 8859 24445
rect 6809 23951 8859 24393
rect 6809 23899 6836 23951
rect 6888 23899 6944 23951
rect 6996 23899 7052 23951
rect 7104 23899 7160 23951
rect 7212 23899 7268 23951
rect 7320 23899 7376 23951
rect 7428 23899 7484 23951
rect 7536 23899 7592 23951
rect 7644 23899 7700 23951
rect 7752 23899 7808 23951
rect 7860 23899 7916 23951
rect 7968 23899 8024 23951
rect 8076 23899 8132 23951
rect 8184 23899 8240 23951
rect 8292 23899 8348 23951
rect 8400 23899 8456 23951
rect 8508 23899 8564 23951
rect 8616 23899 8672 23951
rect 8724 23899 8780 23951
rect 8832 23899 8859 23951
rect 6809 23463 8859 23899
rect 6809 23411 6836 23463
rect 6888 23411 6944 23463
rect 6996 23411 7052 23463
rect 7104 23411 7160 23463
rect 7212 23411 7268 23463
rect 7320 23411 7376 23463
rect 7428 23411 7484 23463
rect 7536 23411 7592 23463
rect 7644 23411 7700 23463
rect 7752 23411 7808 23463
rect 7860 23411 7916 23463
rect 7968 23411 8024 23463
rect 8076 23411 8132 23463
rect 8184 23411 8240 23463
rect 8292 23411 8348 23463
rect 8400 23411 8456 23463
rect 8508 23411 8564 23463
rect 8616 23411 8672 23463
rect 8724 23411 8780 23463
rect 8832 23411 8859 23463
rect 6809 22975 8859 23411
rect 6809 22923 6836 22975
rect 6888 22923 6944 22975
rect 6996 22923 7052 22975
rect 7104 22923 7160 22975
rect 7212 22923 7268 22975
rect 7320 22923 7376 22975
rect 7428 22923 7484 22975
rect 7536 22923 7592 22975
rect 7644 22923 7700 22975
rect 7752 22923 7808 22975
rect 7860 22923 7916 22975
rect 7968 22923 8024 22975
rect 8076 22923 8132 22975
rect 8184 22923 8240 22975
rect 8292 22923 8348 22975
rect 8400 22923 8456 22975
rect 8508 22923 8564 22975
rect 8616 22923 8672 22975
rect 8724 22923 8780 22975
rect 8832 22923 8859 22975
rect 6809 22487 8859 22923
rect 6809 22435 6836 22487
rect 6888 22435 6944 22487
rect 6996 22435 7052 22487
rect 7104 22435 7160 22487
rect 7212 22435 7268 22487
rect 7320 22435 7376 22487
rect 7428 22435 7484 22487
rect 7536 22435 7592 22487
rect 7644 22435 7700 22487
rect 7752 22435 7808 22487
rect 7860 22435 7916 22487
rect 7968 22435 8024 22487
rect 8076 22435 8132 22487
rect 8184 22435 8240 22487
rect 8292 22435 8348 22487
rect 8400 22435 8456 22487
rect 8508 22435 8564 22487
rect 8616 22435 8672 22487
rect 8724 22435 8780 22487
rect 8832 22435 8859 22487
rect 6809 21999 8859 22435
rect 6809 21947 6836 21999
rect 6888 21947 6944 21999
rect 6996 21947 7052 21999
rect 7104 21947 7160 21999
rect 7212 21947 7268 21999
rect 7320 21947 7376 21999
rect 7428 21947 7484 21999
rect 7536 21947 7592 21999
rect 7644 21947 7700 21999
rect 7752 21947 7808 21999
rect 7860 21947 7916 21999
rect 7968 21947 8024 21999
rect 8076 21947 8132 21999
rect 8184 21947 8240 21999
rect 8292 21947 8348 21999
rect 8400 21947 8456 21999
rect 8508 21947 8564 21999
rect 8616 21947 8672 21999
rect 8724 21947 8780 21999
rect 8832 21947 8859 21999
rect 6809 21511 8859 21947
rect 6809 21459 6836 21511
rect 6888 21459 6944 21511
rect 6996 21459 7052 21511
rect 7104 21459 7160 21511
rect 7212 21459 7268 21511
rect 7320 21459 7376 21511
rect 7428 21459 7484 21511
rect 7536 21459 7592 21511
rect 7644 21459 7700 21511
rect 7752 21459 7808 21511
rect 7860 21459 7916 21511
rect 7968 21459 8024 21511
rect 8076 21459 8132 21511
rect 8184 21459 8240 21511
rect 8292 21459 8348 21511
rect 8400 21459 8456 21511
rect 8508 21459 8564 21511
rect 8616 21459 8672 21511
rect 8724 21459 8780 21511
rect 8832 21459 8859 21511
rect 6809 21023 8859 21459
rect 6809 20971 6836 21023
rect 6888 20971 6944 21023
rect 6996 20971 7052 21023
rect 7104 20971 7160 21023
rect 7212 20971 7268 21023
rect 7320 20971 7376 21023
rect 7428 20971 7484 21023
rect 7536 20971 7592 21023
rect 7644 20971 7700 21023
rect 7752 20971 7808 21023
rect 7860 20971 7916 21023
rect 7968 20971 8024 21023
rect 8076 20971 8132 21023
rect 8184 20971 8240 21023
rect 8292 20971 8348 21023
rect 8400 20971 8456 21023
rect 8508 20971 8564 21023
rect 8616 20971 8672 21023
rect 8724 20971 8780 21023
rect 8832 20971 8859 21023
rect 6809 20535 8859 20971
rect 6809 20483 6836 20535
rect 6888 20483 6944 20535
rect 6996 20483 7052 20535
rect 7104 20483 7160 20535
rect 7212 20483 7268 20535
rect 7320 20483 7376 20535
rect 7428 20483 7484 20535
rect 7536 20483 7592 20535
rect 7644 20483 7700 20535
rect 7752 20483 7808 20535
rect 7860 20483 7916 20535
rect 7968 20483 8024 20535
rect 8076 20483 8132 20535
rect 8184 20483 8240 20535
rect 8292 20483 8348 20535
rect 8400 20483 8456 20535
rect 8508 20483 8564 20535
rect 8616 20483 8672 20535
rect 8724 20483 8780 20535
rect 8832 20483 8859 20535
rect 6809 20047 8859 20483
rect 6809 19995 6836 20047
rect 6888 19995 6944 20047
rect 6996 19995 7052 20047
rect 7104 19995 7160 20047
rect 7212 19995 7268 20047
rect 7320 19995 7376 20047
rect 7428 19995 7484 20047
rect 7536 19995 7592 20047
rect 7644 19995 7700 20047
rect 7752 19995 7808 20047
rect 7860 19995 7916 20047
rect 7968 19995 8024 20047
rect 8076 19995 8132 20047
rect 8184 19995 8240 20047
rect 8292 19995 8348 20047
rect 8400 19995 8456 20047
rect 8508 19995 8564 20047
rect 8616 19995 8672 20047
rect 8724 19995 8780 20047
rect 8832 19995 8859 20047
rect 6809 19559 8859 19995
rect 6809 19507 6836 19559
rect 6888 19507 6944 19559
rect 6996 19507 7052 19559
rect 7104 19507 7160 19559
rect 7212 19507 7268 19559
rect 7320 19507 7376 19559
rect 7428 19507 7484 19559
rect 7536 19507 7592 19559
rect 7644 19507 7700 19559
rect 7752 19507 7808 19559
rect 7860 19507 7916 19559
rect 7968 19507 8024 19559
rect 8076 19507 8132 19559
rect 8184 19507 8240 19559
rect 8292 19507 8348 19559
rect 8400 19507 8456 19559
rect 8508 19507 8564 19559
rect 8616 19507 8672 19559
rect 8724 19507 8780 19559
rect 8832 19507 8859 19559
rect 6809 19071 8859 19507
rect 6809 19019 6836 19071
rect 6888 19019 6944 19071
rect 6996 19019 7052 19071
rect 7104 19019 7160 19071
rect 7212 19019 7268 19071
rect 7320 19019 7376 19071
rect 7428 19019 7484 19071
rect 7536 19019 7592 19071
rect 7644 19019 7700 19071
rect 7752 19019 7808 19071
rect 7860 19019 7916 19071
rect 7968 19019 8024 19071
rect 8076 19019 8132 19071
rect 8184 19019 8240 19071
rect 8292 19019 8348 19071
rect 8400 19019 8456 19071
rect 8508 19019 8564 19071
rect 8616 19019 8672 19071
rect 8724 19019 8780 19071
rect 8832 19019 8859 19071
rect 6809 18629 8859 19019
rect 6809 18577 6836 18629
rect 6888 18577 6944 18629
rect 6996 18577 7052 18629
rect 7104 18577 7160 18629
rect 7212 18577 7268 18629
rect 7320 18577 7376 18629
rect 7428 18577 7484 18629
rect 7536 18577 7592 18629
rect 7644 18577 7700 18629
rect 7752 18577 7808 18629
rect 7860 18577 7916 18629
rect 7968 18577 8024 18629
rect 8076 18577 8132 18629
rect 8184 18577 8240 18629
rect 8292 18577 8348 18629
rect 8400 18577 8456 18629
rect 8508 18577 8564 18629
rect 8616 18577 8672 18629
rect 8724 18577 8780 18629
rect 8832 18577 8859 18629
rect 6809 18521 8859 18577
rect 6809 18469 6836 18521
rect 6888 18469 6944 18521
rect 6996 18469 7052 18521
rect 7104 18469 7160 18521
rect 7212 18469 7268 18521
rect 7320 18469 7376 18521
rect 7428 18469 7484 18521
rect 7536 18469 7592 18521
rect 7644 18469 7700 18521
rect 7752 18469 7808 18521
rect 7860 18469 7916 18521
rect 7968 18469 8024 18521
rect 8076 18469 8132 18521
rect 8184 18469 8240 18521
rect 8292 18469 8348 18521
rect 8400 18469 8456 18521
rect 8508 18469 8564 18521
rect 8616 18469 8672 18521
rect 8724 18469 8780 18521
rect 8832 18469 8859 18521
rect 6809 18079 8859 18469
rect 6809 18027 6836 18079
rect 6888 18027 6944 18079
rect 6996 18027 7052 18079
rect 7104 18027 7160 18079
rect 7212 18027 7268 18079
rect 7320 18027 7376 18079
rect 7428 18027 7484 18079
rect 7536 18027 7592 18079
rect 7644 18027 7700 18079
rect 7752 18027 7808 18079
rect 7860 18027 7916 18079
rect 7968 18027 8024 18079
rect 8076 18027 8132 18079
rect 8184 18027 8240 18079
rect 8292 18027 8348 18079
rect 8400 18027 8456 18079
rect 8508 18027 8564 18079
rect 8616 18027 8672 18079
rect 8724 18027 8780 18079
rect 8832 18027 8859 18079
rect 6809 17591 8859 18027
rect 6809 17539 6836 17591
rect 6888 17539 6944 17591
rect 6996 17539 7052 17591
rect 7104 17539 7160 17591
rect 7212 17539 7268 17591
rect 7320 17539 7376 17591
rect 7428 17539 7484 17591
rect 7536 17539 7592 17591
rect 7644 17539 7700 17591
rect 7752 17539 7808 17591
rect 7860 17539 7916 17591
rect 7968 17539 8024 17591
rect 8076 17539 8132 17591
rect 8184 17539 8240 17591
rect 8292 17539 8348 17591
rect 8400 17539 8456 17591
rect 8508 17539 8564 17591
rect 8616 17539 8672 17591
rect 8724 17539 8780 17591
rect 8832 17539 8859 17591
rect 6809 17103 8859 17539
rect 6809 17051 6836 17103
rect 6888 17051 6944 17103
rect 6996 17051 7052 17103
rect 7104 17051 7160 17103
rect 7212 17051 7268 17103
rect 7320 17051 7376 17103
rect 7428 17051 7484 17103
rect 7536 17051 7592 17103
rect 7644 17051 7700 17103
rect 7752 17051 7808 17103
rect 7860 17051 7916 17103
rect 7968 17051 8024 17103
rect 8076 17051 8132 17103
rect 8184 17051 8240 17103
rect 8292 17051 8348 17103
rect 8400 17051 8456 17103
rect 8508 17051 8564 17103
rect 8616 17051 8672 17103
rect 8724 17051 8780 17103
rect 8832 17051 8859 17103
rect 6809 16615 8859 17051
rect 6809 16563 6836 16615
rect 6888 16563 6944 16615
rect 6996 16563 7052 16615
rect 7104 16563 7160 16615
rect 7212 16563 7268 16615
rect 7320 16563 7376 16615
rect 7428 16563 7484 16615
rect 7536 16563 7592 16615
rect 7644 16563 7700 16615
rect 7752 16563 7808 16615
rect 7860 16563 7916 16615
rect 7968 16563 8024 16615
rect 8076 16563 8132 16615
rect 8184 16563 8240 16615
rect 8292 16563 8348 16615
rect 8400 16563 8456 16615
rect 8508 16563 8564 16615
rect 8616 16563 8672 16615
rect 8724 16563 8780 16615
rect 8832 16563 8859 16615
rect 6809 16127 8859 16563
rect 6809 16075 6836 16127
rect 6888 16075 6944 16127
rect 6996 16075 7052 16127
rect 7104 16075 7160 16127
rect 7212 16075 7268 16127
rect 7320 16075 7376 16127
rect 7428 16075 7484 16127
rect 7536 16075 7592 16127
rect 7644 16075 7700 16127
rect 7752 16075 7808 16127
rect 7860 16075 7916 16127
rect 7968 16075 8024 16127
rect 8076 16075 8132 16127
rect 8184 16075 8240 16127
rect 8292 16075 8348 16127
rect 8400 16075 8456 16127
rect 8508 16075 8564 16127
rect 8616 16075 8672 16127
rect 8724 16075 8780 16127
rect 8832 16075 8859 16127
rect 6809 15639 8859 16075
rect 6809 15587 6836 15639
rect 6888 15587 6944 15639
rect 6996 15587 7052 15639
rect 7104 15587 7160 15639
rect 7212 15587 7268 15639
rect 7320 15587 7376 15639
rect 7428 15587 7484 15639
rect 7536 15587 7592 15639
rect 7644 15587 7700 15639
rect 7752 15587 7808 15639
rect 7860 15587 7916 15639
rect 7968 15587 8024 15639
rect 8076 15587 8132 15639
rect 8184 15587 8240 15639
rect 8292 15587 8348 15639
rect 8400 15587 8456 15639
rect 8508 15587 8564 15639
rect 8616 15587 8672 15639
rect 8724 15587 8780 15639
rect 8832 15587 8859 15639
rect 6809 15151 8859 15587
rect 6809 15099 6836 15151
rect 6888 15099 6944 15151
rect 6996 15099 7052 15151
rect 7104 15099 7160 15151
rect 7212 15099 7268 15151
rect 7320 15099 7376 15151
rect 7428 15099 7484 15151
rect 7536 15099 7592 15151
rect 7644 15099 7700 15151
rect 7752 15099 7808 15151
rect 7860 15099 7916 15151
rect 7968 15099 8024 15151
rect 8076 15099 8132 15151
rect 8184 15099 8240 15151
rect 8292 15099 8348 15151
rect 8400 15099 8456 15151
rect 8508 15099 8564 15151
rect 8616 15099 8672 15151
rect 8724 15099 8780 15151
rect 8832 15099 8859 15151
rect 6809 14663 8859 15099
rect 6809 14611 6836 14663
rect 6888 14611 6944 14663
rect 6996 14611 7052 14663
rect 7104 14611 7160 14663
rect 7212 14611 7268 14663
rect 7320 14611 7376 14663
rect 7428 14611 7484 14663
rect 7536 14611 7592 14663
rect 7644 14611 7700 14663
rect 7752 14611 7808 14663
rect 7860 14611 7916 14663
rect 7968 14611 8024 14663
rect 8076 14611 8132 14663
rect 8184 14611 8240 14663
rect 8292 14611 8348 14663
rect 8400 14611 8456 14663
rect 8508 14611 8564 14663
rect 8616 14611 8672 14663
rect 8724 14611 8780 14663
rect 8832 14611 8859 14663
rect 6809 14175 8859 14611
rect 6809 14123 6836 14175
rect 6888 14123 6944 14175
rect 6996 14123 7052 14175
rect 7104 14123 7160 14175
rect 7212 14123 7268 14175
rect 7320 14123 7376 14175
rect 7428 14123 7484 14175
rect 7536 14123 7592 14175
rect 7644 14123 7700 14175
rect 7752 14123 7808 14175
rect 7860 14123 7916 14175
rect 7968 14123 8024 14175
rect 8076 14123 8132 14175
rect 8184 14123 8240 14175
rect 8292 14123 8348 14175
rect 8400 14123 8456 14175
rect 8508 14123 8564 14175
rect 8616 14123 8672 14175
rect 8724 14123 8780 14175
rect 8832 14123 8859 14175
rect 6809 13687 8859 14123
rect 6809 13635 6836 13687
rect 6888 13635 6944 13687
rect 6996 13635 7052 13687
rect 7104 13635 7160 13687
rect 7212 13635 7268 13687
rect 7320 13635 7376 13687
rect 7428 13635 7484 13687
rect 7536 13635 7592 13687
rect 7644 13635 7700 13687
rect 7752 13635 7808 13687
rect 7860 13635 7916 13687
rect 7968 13635 8024 13687
rect 8076 13635 8132 13687
rect 8184 13635 8240 13687
rect 8292 13635 8348 13687
rect 8400 13635 8456 13687
rect 8508 13635 8564 13687
rect 8616 13635 8672 13687
rect 8724 13635 8780 13687
rect 8832 13635 8859 13687
rect 6809 13199 8859 13635
rect 6809 13147 6836 13199
rect 6888 13147 6944 13199
rect 6996 13147 7052 13199
rect 7104 13147 7160 13199
rect 7212 13147 7268 13199
rect 7320 13147 7376 13199
rect 7428 13147 7484 13199
rect 7536 13147 7592 13199
rect 7644 13147 7700 13199
rect 7752 13147 7808 13199
rect 7860 13147 7916 13199
rect 7968 13147 8024 13199
rect 8076 13147 8132 13199
rect 8184 13147 8240 13199
rect 8292 13147 8348 13199
rect 8400 13147 8456 13199
rect 8508 13147 8564 13199
rect 8616 13147 8672 13199
rect 8724 13147 8780 13199
rect 8832 13147 8859 13199
rect 6809 12757 8859 13147
rect 6809 12705 6836 12757
rect 6888 12705 6944 12757
rect 6996 12705 7052 12757
rect 7104 12705 7160 12757
rect 7212 12705 7268 12757
rect 7320 12705 7376 12757
rect 7428 12705 7484 12757
rect 7536 12705 7592 12757
rect 7644 12705 7700 12757
rect 7752 12705 7808 12757
rect 7860 12705 7916 12757
rect 7968 12705 8024 12757
rect 8076 12705 8132 12757
rect 8184 12705 8240 12757
rect 8292 12705 8348 12757
rect 8400 12705 8456 12757
rect 8508 12705 8564 12757
rect 8616 12705 8672 12757
rect 8724 12705 8780 12757
rect 8832 12705 8859 12757
rect 6809 12649 8859 12705
rect 6809 12597 6836 12649
rect 6888 12597 6944 12649
rect 6996 12597 7052 12649
rect 7104 12597 7160 12649
rect 7212 12597 7268 12649
rect 7320 12597 7376 12649
rect 7428 12597 7484 12649
rect 7536 12597 7592 12649
rect 7644 12597 7700 12649
rect 7752 12597 7808 12649
rect 7860 12597 7916 12649
rect 7968 12597 8024 12649
rect 8076 12597 8132 12649
rect 8184 12597 8240 12649
rect 8292 12597 8348 12649
rect 8400 12597 8456 12649
rect 8508 12597 8564 12649
rect 8616 12597 8672 12649
rect 8724 12597 8780 12649
rect 8832 12597 8859 12649
rect 6809 12207 8859 12597
rect 6809 12155 6836 12207
rect 6888 12155 6944 12207
rect 6996 12155 7052 12207
rect 7104 12155 7160 12207
rect 7212 12155 7268 12207
rect 7320 12155 7376 12207
rect 7428 12155 7484 12207
rect 7536 12155 7592 12207
rect 7644 12155 7700 12207
rect 7752 12155 7808 12207
rect 7860 12155 7916 12207
rect 7968 12155 8024 12207
rect 8076 12155 8132 12207
rect 8184 12155 8240 12207
rect 8292 12155 8348 12207
rect 8400 12155 8456 12207
rect 8508 12155 8564 12207
rect 8616 12155 8672 12207
rect 8724 12155 8780 12207
rect 8832 12155 8859 12207
rect 6809 11719 8859 12155
rect 6809 11667 6836 11719
rect 6888 11667 6944 11719
rect 6996 11667 7052 11719
rect 7104 11667 7160 11719
rect 7212 11667 7268 11719
rect 7320 11667 7376 11719
rect 7428 11667 7484 11719
rect 7536 11667 7592 11719
rect 7644 11667 7700 11719
rect 7752 11667 7808 11719
rect 7860 11667 7916 11719
rect 7968 11667 8024 11719
rect 8076 11667 8132 11719
rect 8184 11667 8240 11719
rect 8292 11667 8348 11719
rect 8400 11667 8456 11719
rect 8508 11667 8564 11719
rect 8616 11667 8672 11719
rect 8724 11667 8780 11719
rect 8832 11667 8859 11719
rect 6809 11231 8859 11667
rect 6809 11179 6836 11231
rect 6888 11179 6944 11231
rect 6996 11179 7052 11231
rect 7104 11179 7160 11231
rect 7212 11179 7268 11231
rect 7320 11179 7376 11231
rect 7428 11179 7484 11231
rect 7536 11179 7592 11231
rect 7644 11179 7700 11231
rect 7752 11179 7808 11231
rect 7860 11179 7916 11231
rect 7968 11179 8024 11231
rect 8076 11179 8132 11231
rect 8184 11179 8240 11231
rect 8292 11179 8348 11231
rect 8400 11179 8456 11231
rect 8508 11179 8564 11231
rect 8616 11179 8672 11231
rect 8724 11179 8780 11231
rect 8832 11179 8859 11231
rect 6809 10743 8859 11179
rect 6809 10691 6836 10743
rect 6888 10691 6944 10743
rect 6996 10691 7052 10743
rect 7104 10691 7160 10743
rect 7212 10691 7268 10743
rect 7320 10691 7376 10743
rect 7428 10691 7484 10743
rect 7536 10691 7592 10743
rect 7644 10691 7700 10743
rect 7752 10691 7808 10743
rect 7860 10691 7916 10743
rect 7968 10691 8024 10743
rect 8076 10691 8132 10743
rect 8184 10691 8240 10743
rect 8292 10691 8348 10743
rect 8400 10691 8456 10743
rect 8508 10691 8564 10743
rect 8616 10691 8672 10743
rect 8724 10691 8780 10743
rect 8832 10691 8859 10743
rect 6809 10255 8859 10691
rect 6809 10203 6836 10255
rect 6888 10203 6944 10255
rect 6996 10203 7052 10255
rect 7104 10203 7160 10255
rect 7212 10203 7268 10255
rect 7320 10203 7376 10255
rect 7428 10203 7484 10255
rect 7536 10203 7592 10255
rect 7644 10203 7700 10255
rect 7752 10203 7808 10255
rect 7860 10203 7916 10255
rect 7968 10203 8024 10255
rect 8076 10203 8132 10255
rect 8184 10203 8240 10255
rect 8292 10203 8348 10255
rect 8400 10203 8456 10255
rect 8508 10203 8564 10255
rect 8616 10203 8672 10255
rect 8724 10203 8780 10255
rect 8832 10203 8859 10255
rect 6809 9767 8859 10203
rect 6809 9715 6836 9767
rect 6888 9715 6944 9767
rect 6996 9715 7052 9767
rect 7104 9715 7160 9767
rect 7212 9715 7268 9767
rect 7320 9715 7376 9767
rect 7428 9715 7484 9767
rect 7536 9715 7592 9767
rect 7644 9715 7700 9767
rect 7752 9715 7808 9767
rect 7860 9715 7916 9767
rect 7968 9715 8024 9767
rect 8076 9715 8132 9767
rect 8184 9715 8240 9767
rect 8292 9715 8348 9767
rect 8400 9715 8456 9767
rect 8508 9715 8564 9767
rect 8616 9715 8672 9767
rect 8724 9715 8780 9767
rect 8832 9715 8859 9767
rect 6809 9279 8859 9715
rect 6809 9227 6836 9279
rect 6888 9227 6944 9279
rect 6996 9227 7052 9279
rect 7104 9227 7160 9279
rect 7212 9227 7268 9279
rect 7320 9227 7376 9279
rect 7428 9227 7484 9279
rect 7536 9227 7592 9279
rect 7644 9227 7700 9279
rect 7752 9227 7808 9279
rect 7860 9227 7916 9279
rect 7968 9227 8024 9279
rect 8076 9227 8132 9279
rect 8184 9227 8240 9279
rect 8292 9227 8348 9279
rect 8400 9227 8456 9279
rect 8508 9227 8564 9279
rect 8616 9227 8672 9279
rect 8724 9227 8780 9279
rect 8832 9227 8859 9279
rect 6809 8791 8859 9227
rect 6809 8739 6836 8791
rect 6888 8739 6944 8791
rect 6996 8739 7052 8791
rect 7104 8739 7160 8791
rect 7212 8739 7268 8791
rect 7320 8739 7376 8791
rect 7428 8739 7484 8791
rect 7536 8739 7592 8791
rect 7644 8739 7700 8791
rect 7752 8739 7808 8791
rect 7860 8739 7916 8791
rect 7968 8739 8024 8791
rect 8076 8739 8132 8791
rect 8184 8739 8240 8791
rect 8292 8739 8348 8791
rect 8400 8739 8456 8791
rect 8508 8739 8564 8791
rect 8616 8739 8672 8791
rect 8724 8739 8780 8791
rect 8832 8739 8859 8791
rect 6809 8303 8859 8739
rect 6809 8251 6836 8303
rect 6888 8251 6944 8303
rect 6996 8251 7052 8303
rect 7104 8251 7160 8303
rect 7212 8251 7268 8303
rect 7320 8251 7376 8303
rect 7428 8251 7484 8303
rect 7536 8251 7592 8303
rect 7644 8251 7700 8303
rect 7752 8251 7808 8303
rect 7860 8251 7916 8303
rect 7968 8251 8024 8303
rect 8076 8251 8132 8303
rect 8184 8251 8240 8303
rect 8292 8251 8348 8303
rect 8400 8251 8456 8303
rect 8508 8251 8564 8303
rect 8616 8251 8672 8303
rect 8724 8251 8780 8303
rect 8832 8251 8859 8303
rect 6809 7815 8859 8251
rect 6809 7763 6836 7815
rect 6888 7763 6944 7815
rect 6996 7763 7052 7815
rect 7104 7763 7160 7815
rect 7212 7763 7268 7815
rect 7320 7763 7376 7815
rect 7428 7763 7484 7815
rect 7536 7763 7592 7815
rect 7644 7763 7700 7815
rect 7752 7763 7808 7815
rect 7860 7763 7916 7815
rect 7968 7763 8024 7815
rect 8076 7763 8132 7815
rect 8184 7763 8240 7815
rect 8292 7763 8348 7815
rect 8400 7763 8456 7815
rect 8508 7763 8564 7815
rect 8616 7763 8672 7815
rect 8724 7763 8780 7815
rect 8832 7763 8859 7815
rect 6809 7327 8859 7763
rect 6809 7275 6836 7327
rect 6888 7275 6944 7327
rect 6996 7275 7052 7327
rect 7104 7275 7160 7327
rect 7212 7275 7268 7327
rect 7320 7275 7376 7327
rect 7428 7275 7484 7327
rect 7536 7275 7592 7327
rect 7644 7275 7700 7327
rect 7752 7275 7808 7327
rect 7860 7275 7916 7327
rect 7968 7275 8024 7327
rect 8076 7275 8132 7327
rect 8184 7275 8240 7327
rect 8292 7275 8348 7327
rect 8400 7275 8456 7327
rect 8508 7275 8564 7327
rect 8616 7275 8672 7327
rect 8724 7275 8780 7327
rect 8832 7275 8859 7327
rect 6809 6885 8859 7275
rect 6809 6833 6836 6885
rect 6888 6833 6944 6885
rect 6996 6833 7052 6885
rect 7104 6833 7160 6885
rect 7212 6833 7268 6885
rect 7320 6833 7376 6885
rect 7428 6833 7484 6885
rect 7536 6833 7592 6885
rect 7644 6833 7700 6885
rect 7752 6833 7808 6885
rect 7860 6833 7916 6885
rect 7968 6833 8024 6885
rect 8076 6833 8132 6885
rect 8184 6833 8240 6885
rect 8292 6833 8348 6885
rect 8400 6833 8456 6885
rect 8508 6833 8564 6885
rect 8616 6833 8672 6885
rect 8724 6833 8780 6885
rect 8832 6833 8859 6885
rect 6809 6777 8859 6833
rect 6809 6725 6836 6777
rect 6888 6725 6944 6777
rect 6996 6725 7052 6777
rect 7104 6725 7160 6777
rect 7212 6725 7268 6777
rect 7320 6725 7376 6777
rect 7428 6725 7484 6777
rect 7536 6725 7592 6777
rect 7644 6725 7700 6777
rect 7752 6725 7808 6777
rect 7860 6725 7916 6777
rect 7968 6725 8024 6777
rect 8076 6725 8132 6777
rect 8184 6725 8240 6777
rect 8292 6725 8348 6777
rect 8400 6725 8456 6777
rect 8508 6725 8564 6777
rect 8616 6725 8672 6777
rect 8724 6725 8780 6777
rect 8832 6725 8859 6777
rect 6809 6335 8859 6725
rect 6809 6283 6836 6335
rect 6888 6283 6944 6335
rect 6996 6283 7052 6335
rect 7104 6283 7160 6335
rect 7212 6283 7268 6335
rect 7320 6283 7376 6335
rect 7428 6283 7484 6335
rect 7536 6283 7592 6335
rect 7644 6283 7700 6335
rect 7752 6283 7808 6335
rect 7860 6283 7916 6335
rect 7968 6283 8024 6335
rect 8076 6283 8132 6335
rect 8184 6283 8240 6335
rect 8292 6283 8348 6335
rect 8400 6283 8456 6335
rect 8508 6283 8564 6335
rect 8616 6283 8672 6335
rect 8724 6283 8780 6335
rect 8832 6283 8859 6335
rect 6809 5847 8859 6283
rect 6809 5795 6836 5847
rect 6888 5795 6944 5847
rect 6996 5795 7052 5847
rect 7104 5795 7160 5847
rect 7212 5795 7268 5847
rect 7320 5795 7376 5847
rect 7428 5795 7484 5847
rect 7536 5795 7592 5847
rect 7644 5795 7700 5847
rect 7752 5795 7808 5847
rect 7860 5795 7916 5847
rect 7968 5795 8024 5847
rect 8076 5795 8132 5847
rect 8184 5795 8240 5847
rect 8292 5795 8348 5847
rect 8400 5795 8456 5847
rect 8508 5795 8564 5847
rect 8616 5795 8672 5847
rect 8724 5795 8780 5847
rect 8832 5795 8859 5847
rect 6809 5359 8859 5795
rect 6809 5307 6836 5359
rect 6888 5307 6944 5359
rect 6996 5307 7052 5359
rect 7104 5307 7160 5359
rect 7212 5307 7268 5359
rect 7320 5307 7376 5359
rect 7428 5307 7484 5359
rect 7536 5307 7592 5359
rect 7644 5307 7700 5359
rect 7752 5307 7808 5359
rect 7860 5307 7916 5359
rect 7968 5307 8024 5359
rect 8076 5307 8132 5359
rect 8184 5307 8240 5359
rect 8292 5307 8348 5359
rect 8400 5307 8456 5359
rect 8508 5307 8564 5359
rect 8616 5307 8672 5359
rect 8724 5307 8780 5359
rect 8832 5307 8859 5359
rect 6809 4871 8859 5307
rect 6809 4819 6836 4871
rect 6888 4819 6944 4871
rect 6996 4819 7052 4871
rect 7104 4819 7160 4871
rect 7212 4819 7268 4871
rect 7320 4819 7376 4871
rect 7428 4819 7484 4871
rect 7536 4819 7592 4871
rect 7644 4819 7700 4871
rect 7752 4819 7808 4871
rect 7860 4819 7916 4871
rect 7968 4819 8024 4871
rect 8076 4819 8132 4871
rect 8184 4819 8240 4871
rect 8292 4819 8348 4871
rect 8400 4819 8456 4871
rect 8508 4819 8564 4871
rect 8616 4819 8672 4871
rect 8724 4819 8780 4871
rect 8832 4819 8859 4871
rect 6809 4383 8859 4819
rect 6809 4331 6836 4383
rect 6888 4331 6944 4383
rect 6996 4331 7052 4383
rect 7104 4331 7160 4383
rect 7212 4331 7268 4383
rect 7320 4331 7376 4383
rect 7428 4331 7484 4383
rect 7536 4331 7592 4383
rect 7644 4331 7700 4383
rect 7752 4331 7808 4383
rect 7860 4331 7916 4383
rect 7968 4331 8024 4383
rect 8076 4331 8132 4383
rect 8184 4331 8240 4383
rect 8292 4331 8348 4383
rect 8400 4331 8456 4383
rect 8508 4331 8564 4383
rect 8616 4331 8672 4383
rect 8724 4331 8780 4383
rect 8832 4331 8859 4383
rect 6809 3895 8859 4331
rect 6809 3843 6836 3895
rect 6888 3843 6944 3895
rect 6996 3843 7052 3895
rect 7104 3843 7160 3895
rect 7212 3843 7268 3895
rect 7320 3843 7376 3895
rect 7428 3843 7484 3895
rect 7536 3843 7592 3895
rect 7644 3843 7700 3895
rect 7752 3843 7808 3895
rect 7860 3843 7916 3895
rect 7968 3843 8024 3895
rect 8076 3843 8132 3895
rect 8184 3843 8240 3895
rect 8292 3843 8348 3895
rect 8400 3843 8456 3895
rect 8508 3843 8564 3895
rect 8616 3843 8672 3895
rect 8724 3843 8780 3895
rect 8832 3843 8859 3895
rect 6809 3407 8859 3843
rect 6809 3355 6836 3407
rect 6888 3355 6944 3407
rect 6996 3355 7052 3407
rect 7104 3355 7160 3407
rect 7212 3355 7268 3407
rect 7320 3355 7376 3407
rect 7428 3355 7484 3407
rect 7536 3355 7592 3407
rect 7644 3355 7700 3407
rect 7752 3355 7808 3407
rect 7860 3355 7916 3407
rect 7968 3355 8024 3407
rect 8076 3355 8132 3407
rect 8184 3355 8240 3407
rect 8292 3355 8348 3407
rect 8400 3355 8456 3407
rect 8508 3355 8564 3407
rect 8616 3355 8672 3407
rect 8724 3355 8780 3407
rect 8832 3355 8859 3407
rect 6809 2919 8859 3355
rect 6809 2867 6836 2919
rect 6888 2867 6944 2919
rect 6996 2867 7052 2919
rect 7104 2867 7160 2919
rect 7212 2867 7268 2919
rect 7320 2867 7376 2919
rect 7428 2867 7484 2919
rect 7536 2867 7592 2919
rect 7644 2867 7700 2919
rect 7752 2867 7808 2919
rect 7860 2867 7916 2919
rect 7968 2867 8024 2919
rect 8076 2867 8132 2919
rect 8184 2867 8240 2919
rect 8292 2867 8348 2919
rect 8400 2867 8456 2919
rect 8508 2867 8564 2919
rect 8616 2867 8672 2919
rect 8724 2867 8780 2919
rect 8832 2867 8859 2919
rect 6809 2431 8859 2867
rect 6809 2379 6836 2431
rect 6888 2379 6944 2431
rect 6996 2379 7052 2431
rect 7104 2379 7160 2431
rect 7212 2379 7268 2431
rect 7320 2379 7376 2431
rect 7428 2379 7484 2431
rect 7536 2379 7592 2431
rect 7644 2379 7700 2431
rect 7752 2379 7808 2431
rect 7860 2379 7916 2431
rect 7968 2379 8024 2431
rect 8076 2379 8132 2431
rect 8184 2379 8240 2431
rect 8292 2379 8348 2431
rect 8400 2379 8456 2431
rect 8508 2379 8564 2431
rect 8616 2379 8672 2431
rect 8724 2379 8780 2431
rect 8832 2379 8859 2431
rect 6809 1943 8859 2379
rect 6809 1891 6836 1943
rect 6888 1891 6944 1943
rect 6996 1891 7052 1943
rect 7104 1891 7160 1943
rect 7212 1891 7268 1943
rect 7320 1891 7376 1943
rect 7428 1891 7484 1943
rect 7536 1891 7592 1943
rect 7644 1891 7700 1943
rect 7752 1891 7808 1943
rect 7860 1891 7916 1943
rect 7968 1891 8024 1943
rect 8076 1891 8132 1943
rect 8184 1891 8240 1943
rect 8292 1891 8348 1943
rect 8400 1891 8456 1943
rect 8508 1891 8564 1943
rect 8616 1891 8672 1943
rect 8724 1891 8780 1943
rect 8832 1891 8859 1943
rect 6809 1455 8859 1891
rect 6809 1403 6836 1455
rect 6888 1403 6944 1455
rect 6996 1403 7052 1455
rect 7104 1403 7160 1455
rect 7212 1403 7268 1455
rect 7320 1403 7376 1455
rect 7428 1403 7484 1455
rect 7536 1403 7592 1455
rect 7644 1403 7700 1455
rect 7752 1403 7808 1455
rect 7860 1403 7916 1455
rect 7968 1403 8024 1455
rect 8076 1403 8132 1455
rect 8184 1403 8240 1455
rect 8292 1403 8348 1455
rect 8400 1403 8456 1455
rect 8508 1403 8564 1455
rect 8616 1403 8672 1455
rect 8724 1403 8780 1455
rect 8832 1403 8859 1455
rect 6809 961 8859 1403
rect 6809 909 6836 961
rect 6888 909 6944 961
rect 6996 909 7052 961
rect 7104 909 7160 961
rect 7212 909 7268 961
rect 7320 909 7376 961
rect 7428 909 7484 961
rect 7536 909 7592 961
rect 7644 909 7700 961
rect 7752 909 7808 961
rect 7860 909 7916 961
rect 7968 909 8024 961
rect 8076 909 8132 961
rect 8184 909 8240 961
rect 8292 909 8348 961
rect 8400 909 8456 961
rect 8508 909 8564 961
rect 8616 909 8672 961
rect 8724 909 8780 961
rect 8832 909 8859 961
rect 6809 853 8859 909
rect 6809 801 6836 853
rect 6888 801 6944 853
rect 6996 801 7052 853
rect 7104 801 7160 853
rect 7212 801 7268 853
rect 7320 801 7376 853
rect 7428 801 7484 853
rect 7536 801 7592 853
rect 7644 801 7700 853
rect 7752 801 7808 853
rect 7860 801 7916 853
rect 7968 801 8024 853
rect 8076 801 8132 853
rect 8184 801 8240 853
rect 8292 801 8348 853
rect 8400 801 8456 853
rect 8508 801 8564 853
rect 8616 801 8672 853
rect 8724 801 8780 853
rect 8832 801 8859 853
rect 6809 745 8859 801
rect 6809 693 6836 745
rect 6888 693 6944 745
rect 6996 693 7052 745
rect 7104 693 7160 745
rect 7212 693 7268 745
rect 7320 693 7376 745
rect 7428 693 7484 745
rect 7536 693 7592 745
rect 7644 693 7700 745
rect 7752 693 7808 745
rect 7860 693 7916 745
rect 7968 693 8024 745
rect 8076 693 8132 745
rect 8184 693 8240 745
rect 8292 693 8348 745
rect 8400 693 8456 745
rect 8508 693 8564 745
rect 8616 693 8672 745
rect 8724 693 8780 745
rect 8832 693 8859 745
rect 6809 43 8859 693
rect 8919 25261 9119 25617
rect 8919 25209 8939 25261
rect 8991 25209 9047 25261
rect 9099 25209 9119 25261
rect 8919 25153 9119 25209
rect 8919 25101 8939 25153
rect 8991 25101 9047 25153
rect 9099 25101 9119 25153
rect 8919 25045 9119 25101
rect 8919 24993 8939 25045
rect 8991 24993 9047 25045
rect 9099 24993 9119 25045
rect 8919 23707 9119 24993
rect 8919 23655 8939 23707
rect 8991 23655 9047 23707
rect 9099 23655 9119 23707
rect 8919 23219 9119 23655
rect 8919 23167 8939 23219
rect 8991 23167 9047 23219
rect 9099 23167 9119 23219
rect 8919 22731 9119 23167
rect 8919 22679 8939 22731
rect 8991 22679 9047 22731
rect 9099 22679 9119 22731
rect 8919 22243 9119 22679
rect 8919 22191 8939 22243
rect 8991 22191 9047 22243
rect 9099 22191 9119 22243
rect 8919 21755 9119 22191
rect 8919 21703 8939 21755
rect 8991 21703 9047 21755
rect 9099 21703 9119 21755
rect 8919 21267 9119 21703
rect 8919 21215 8939 21267
rect 8991 21215 9047 21267
rect 9099 21215 9119 21267
rect 8919 20779 9119 21215
rect 8919 20727 8939 20779
rect 8991 20727 9047 20779
rect 9099 20727 9119 20779
rect 8919 20291 9119 20727
rect 8919 20239 8939 20291
rect 8991 20239 9047 20291
rect 9099 20239 9119 20291
rect 8919 19803 9119 20239
rect 8919 19751 8939 19803
rect 8991 19751 9047 19803
rect 9099 19751 9119 19803
rect 8919 19315 9119 19751
rect 8919 19263 8939 19315
rect 8991 19263 9047 19315
rect 9099 19263 9119 19315
rect 8919 17835 9119 19263
rect 8919 17783 8939 17835
rect 8991 17783 9047 17835
rect 9099 17783 9119 17835
rect 8919 17347 9119 17783
rect 8919 17295 8939 17347
rect 8991 17295 9047 17347
rect 9099 17295 9119 17347
rect 8919 16859 9119 17295
rect 8919 16807 8939 16859
rect 8991 16807 9047 16859
rect 9099 16807 9119 16859
rect 8919 16371 9119 16807
rect 8919 16319 8939 16371
rect 8991 16319 9047 16371
rect 9099 16319 9119 16371
rect 8919 15883 9119 16319
rect 8919 15831 8939 15883
rect 8991 15831 9047 15883
rect 9099 15831 9119 15883
rect 8919 15395 9119 15831
rect 8919 15343 8939 15395
rect 8991 15343 9047 15395
rect 9099 15343 9119 15395
rect 8919 14907 9119 15343
rect 8919 14855 8939 14907
rect 8991 14855 9047 14907
rect 9099 14855 9119 14907
rect 8919 14419 9119 14855
rect 8919 14367 8939 14419
rect 8991 14367 9047 14419
rect 9099 14367 9119 14419
rect 8919 13931 9119 14367
rect 8919 13879 8939 13931
rect 8991 13879 9047 13931
rect 9099 13879 9119 13931
rect 8919 13443 9119 13879
rect 8919 13391 8939 13443
rect 8991 13391 9047 13443
rect 9099 13391 9119 13443
rect 8919 11963 9119 13391
rect 8919 11911 8939 11963
rect 8991 11911 9047 11963
rect 9099 11911 9119 11963
rect 8919 11475 9119 11911
rect 8919 11423 8939 11475
rect 8991 11423 9047 11475
rect 9099 11423 9119 11475
rect 8919 10987 9119 11423
rect 8919 10935 8939 10987
rect 8991 10935 9047 10987
rect 9099 10935 9119 10987
rect 8919 10499 9119 10935
rect 8919 10447 8939 10499
rect 8991 10447 9047 10499
rect 9099 10447 9119 10499
rect 8919 10011 9119 10447
rect 8919 9959 8939 10011
rect 8991 9959 9047 10011
rect 9099 9959 9119 10011
rect 8919 9523 9119 9959
rect 8919 9471 8939 9523
rect 8991 9471 9047 9523
rect 9099 9471 9119 9523
rect 8919 9035 9119 9471
rect 8919 8983 8939 9035
rect 8991 8983 9047 9035
rect 9099 8983 9119 9035
rect 8919 8547 9119 8983
rect 8919 8495 8939 8547
rect 8991 8495 9047 8547
rect 9099 8495 9119 8547
rect 8919 8059 9119 8495
rect 8919 8007 8939 8059
rect 8991 8007 9047 8059
rect 9099 8007 9119 8059
rect 8919 7571 9119 8007
rect 8919 7519 8939 7571
rect 8991 7519 9047 7571
rect 9099 7519 9119 7571
rect 8919 6091 9119 7519
rect 8919 6039 8939 6091
rect 8991 6039 9047 6091
rect 9099 6039 9119 6091
rect 8919 5603 9119 6039
rect 8919 5551 8939 5603
rect 8991 5551 9047 5603
rect 9099 5551 9119 5603
rect 8919 5115 9119 5551
rect 8919 5063 8939 5115
rect 8991 5063 9047 5115
rect 9099 5063 9119 5115
rect 8919 4627 9119 5063
rect 8919 4575 8939 4627
rect 8991 4575 9047 4627
rect 9099 4575 9119 4627
rect 8919 4139 9119 4575
rect 8919 4087 8939 4139
rect 8991 4087 9047 4139
rect 9099 4087 9119 4139
rect 8919 3651 9119 4087
rect 8919 3599 8939 3651
rect 8991 3599 9047 3651
rect 9099 3599 9119 3651
rect 8919 3163 9119 3599
rect 8919 3111 8939 3163
rect 8991 3111 9047 3163
rect 9099 3111 9119 3163
rect 8919 2675 9119 3111
rect 8919 2623 8939 2675
rect 8991 2623 9047 2675
rect 9099 2623 9119 2675
rect 8919 2187 9119 2623
rect 8919 2135 8939 2187
rect 8991 2135 9047 2187
rect 9099 2135 9119 2187
rect 8919 1699 9119 2135
rect 8919 1647 8939 1699
rect 8991 1647 9047 1699
rect 9099 1647 9119 1699
rect 8919 361 9119 1647
rect 8919 309 8939 361
rect 8991 309 9047 361
rect 9099 309 9119 361
rect 8919 253 9119 309
rect 8919 201 8939 253
rect 8991 201 9047 253
rect 9099 201 9119 253
rect 8919 145 9119 201
rect 8919 93 8939 145
rect 8991 93 9047 145
rect 9099 93 9119 145
rect 8919 43 9119 93
rect 9179 24661 11229 25617
rect 9179 24609 9206 24661
rect 9258 24609 9314 24661
rect 9366 24609 9422 24661
rect 9474 24609 9530 24661
rect 9582 24609 9638 24661
rect 9690 24609 9746 24661
rect 9798 24609 9854 24661
rect 9906 24609 9962 24661
rect 10014 24609 10070 24661
rect 10122 24609 10178 24661
rect 10230 24609 10286 24661
rect 10338 24609 10394 24661
rect 10446 24609 10502 24661
rect 10554 24609 10610 24661
rect 10662 24609 10718 24661
rect 10770 24609 10826 24661
rect 10878 24609 10934 24661
rect 10986 24609 11042 24661
rect 11094 24609 11150 24661
rect 11202 24609 11229 24661
rect 9179 24553 11229 24609
rect 9179 24501 9206 24553
rect 9258 24501 9314 24553
rect 9366 24501 9422 24553
rect 9474 24501 9530 24553
rect 9582 24501 9638 24553
rect 9690 24501 9746 24553
rect 9798 24501 9854 24553
rect 9906 24501 9962 24553
rect 10014 24501 10070 24553
rect 10122 24501 10178 24553
rect 10230 24501 10286 24553
rect 10338 24501 10394 24553
rect 10446 24501 10502 24553
rect 10554 24501 10610 24553
rect 10662 24501 10718 24553
rect 10770 24501 10826 24553
rect 10878 24501 10934 24553
rect 10986 24501 11042 24553
rect 11094 24501 11150 24553
rect 11202 24501 11229 24553
rect 9179 24445 11229 24501
rect 9179 24393 9206 24445
rect 9258 24393 9314 24445
rect 9366 24393 9422 24445
rect 9474 24393 9530 24445
rect 9582 24393 9638 24445
rect 9690 24393 9746 24445
rect 9798 24393 9854 24445
rect 9906 24393 9962 24445
rect 10014 24393 10070 24445
rect 10122 24393 10178 24445
rect 10230 24393 10286 24445
rect 10338 24393 10394 24445
rect 10446 24393 10502 24445
rect 10554 24393 10610 24445
rect 10662 24393 10718 24445
rect 10770 24393 10826 24445
rect 10878 24393 10934 24445
rect 10986 24393 11042 24445
rect 11094 24393 11150 24445
rect 11202 24393 11229 24445
rect 9179 23951 11229 24393
rect 9179 23899 9206 23951
rect 9258 23899 9314 23951
rect 9366 23899 9422 23951
rect 9474 23899 9530 23951
rect 9582 23899 9638 23951
rect 9690 23899 9746 23951
rect 9798 23899 9854 23951
rect 9906 23899 9962 23951
rect 10014 23899 10070 23951
rect 10122 23899 10178 23951
rect 10230 23899 10286 23951
rect 10338 23899 10394 23951
rect 10446 23899 10502 23951
rect 10554 23899 10610 23951
rect 10662 23899 10718 23951
rect 10770 23899 10826 23951
rect 10878 23899 10934 23951
rect 10986 23899 11042 23951
rect 11094 23899 11150 23951
rect 11202 23899 11229 23951
rect 9179 23463 11229 23899
rect 9179 23411 9206 23463
rect 9258 23411 9314 23463
rect 9366 23411 9422 23463
rect 9474 23411 9530 23463
rect 9582 23411 9638 23463
rect 9690 23411 9746 23463
rect 9798 23411 9854 23463
rect 9906 23411 9962 23463
rect 10014 23411 10070 23463
rect 10122 23411 10178 23463
rect 10230 23411 10286 23463
rect 10338 23411 10394 23463
rect 10446 23411 10502 23463
rect 10554 23411 10610 23463
rect 10662 23411 10718 23463
rect 10770 23411 10826 23463
rect 10878 23411 10934 23463
rect 10986 23411 11042 23463
rect 11094 23411 11150 23463
rect 11202 23411 11229 23463
rect 9179 22975 11229 23411
rect 9179 22923 9206 22975
rect 9258 22923 9314 22975
rect 9366 22923 9422 22975
rect 9474 22923 9530 22975
rect 9582 22923 9638 22975
rect 9690 22923 9746 22975
rect 9798 22923 9854 22975
rect 9906 22923 9962 22975
rect 10014 22923 10070 22975
rect 10122 22923 10178 22975
rect 10230 22923 10286 22975
rect 10338 22923 10394 22975
rect 10446 22923 10502 22975
rect 10554 22923 10610 22975
rect 10662 22923 10718 22975
rect 10770 22923 10826 22975
rect 10878 22923 10934 22975
rect 10986 22923 11042 22975
rect 11094 22923 11150 22975
rect 11202 22923 11229 22975
rect 9179 22487 11229 22923
rect 9179 22435 9206 22487
rect 9258 22435 9314 22487
rect 9366 22435 9422 22487
rect 9474 22435 9530 22487
rect 9582 22435 9638 22487
rect 9690 22435 9746 22487
rect 9798 22435 9854 22487
rect 9906 22435 9962 22487
rect 10014 22435 10070 22487
rect 10122 22435 10178 22487
rect 10230 22435 10286 22487
rect 10338 22435 10394 22487
rect 10446 22435 10502 22487
rect 10554 22435 10610 22487
rect 10662 22435 10718 22487
rect 10770 22435 10826 22487
rect 10878 22435 10934 22487
rect 10986 22435 11042 22487
rect 11094 22435 11150 22487
rect 11202 22435 11229 22487
rect 9179 21999 11229 22435
rect 9179 21947 9206 21999
rect 9258 21947 9314 21999
rect 9366 21947 9422 21999
rect 9474 21947 9530 21999
rect 9582 21947 9638 21999
rect 9690 21947 9746 21999
rect 9798 21947 9854 21999
rect 9906 21947 9962 21999
rect 10014 21947 10070 21999
rect 10122 21947 10178 21999
rect 10230 21947 10286 21999
rect 10338 21947 10394 21999
rect 10446 21947 10502 21999
rect 10554 21947 10610 21999
rect 10662 21947 10718 21999
rect 10770 21947 10826 21999
rect 10878 21947 10934 21999
rect 10986 21947 11042 21999
rect 11094 21947 11150 21999
rect 11202 21947 11229 21999
rect 9179 21511 11229 21947
rect 9179 21459 9206 21511
rect 9258 21459 9314 21511
rect 9366 21459 9422 21511
rect 9474 21459 9530 21511
rect 9582 21459 9638 21511
rect 9690 21459 9746 21511
rect 9798 21459 9854 21511
rect 9906 21459 9962 21511
rect 10014 21459 10070 21511
rect 10122 21459 10178 21511
rect 10230 21459 10286 21511
rect 10338 21459 10394 21511
rect 10446 21459 10502 21511
rect 10554 21459 10610 21511
rect 10662 21459 10718 21511
rect 10770 21459 10826 21511
rect 10878 21459 10934 21511
rect 10986 21459 11042 21511
rect 11094 21459 11150 21511
rect 11202 21459 11229 21511
rect 9179 21023 11229 21459
rect 9179 20971 9206 21023
rect 9258 20971 9314 21023
rect 9366 20971 9422 21023
rect 9474 20971 9530 21023
rect 9582 20971 9638 21023
rect 9690 20971 9746 21023
rect 9798 20971 9854 21023
rect 9906 20971 9962 21023
rect 10014 20971 10070 21023
rect 10122 20971 10178 21023
rect 10230 20971 10286 21023
rect 10338 20971 10394 21023
rect 10446 20971 10502 21023
rect 10554 20971 10610 21023
rect 10662 20971 10718 21023
rect 10770 20971 10826 21023
rect 10878 20971 10934 21023
rect 10986 20971 11042 21023
rect 11094 20971 11150 21023
rect 11202 20971 11229 21023
rect 9179 20535 11229 20971
rect 9179 20483 9206 20535
rect 9258 20483 9314 20535
rect 9366 20483 9422 20535
rect 9474 20483 9530 20535
rect 9582 20483 9638 20535
rect 9690 20483 9746 20535
rect 9798 20483 9854 20535
rect 9906 20483 9962 20535
rect 10014 20483 10070 20535
rect 10122 20483 10178 20535
rect 10230 20483 10286 20535
rect 10338 20483 10394 20535
rect 10446 20483 10502 20535
rect 10554 20483 10610 20535
rect 10662 20483 10718 20535
rect 10770 20483 10826 20535
rect 10878 20483 10934 20535
rect 10986 20483 11042 20535
rect 11094 20483 11150 20535
rect 11202 20483 11229 20535
rect 9179 20047 11229 20483
rect 9179 19995 9206 20047
rect 9258 19995 9314 20047
rect 9366 19995 9422 20047
rect 9474 19995 9530 20047
rect 9582 19995 9638 20047
rect 9690 19995 9746 20047
rect 9798 19995 9854 20047
rect 9906 19995 9962 20047
rect 10014 19995 10070 20047
rect 10122 19995 10178 20047
rect 10230 19995 10286 20047
rect 10338 19995 10394 20047
rect 10446 19995 10502 20047
rect 10554 19995 10610 20047
rect 10662 19995 10718 20047
rect 10770 19995 10826 20047
rect 10878 19995 10934 20047
rect 10986 19995 11042 20047
rect 11094 19995 11150 20047
rect 11202 19995 11229 20047
rect 9179 19559 11229 19995
rect 9179 19507 9206 19559
rect 9258 19507 9314 19559
rect 9366 19507 9422 19559
rect 9474 19507 9530 19559
rect 9582 19507 9638 19559
rect 9690 19507 9746 19559
rect 9798 19507 9854 19559
rect 9906 19507 9962 19559
rect 10014 19507 10070 19559
rect 10122 19507 10178 19559
rect 10230 19507 10286 19559
rect 10338 19507 10394 19559
rect 10446 19507 10502 19559
rect 10554 19507 10610 19559
rect 10662 19507 10718 19559
rect 10770 19507 10826 19559
rect 10878 19507 10934 19559
rect 10986 19507 11042 19559
rect 11094 19507 11150 19559
rect 11202 19507 11229 19559
rect 9179 19071 11229 19507
rect 9179 19019 9206 19071
rect 9258 19019 9314 19071
rect 9366 19019 9422 19071
rect 9474 19019 9530 19071
rect 9582 19019 9638 19071
rect 9690 19019 9746 19071
rect 9798 19019 9854 19071
rect 9906 19019 9962 19071
rect 10014 19019 10070 19071
rect 10122 19019 10178 19071
rect 10230 19019 10286 19071
rect 10338 19019 10394 19071
rect 10446 19019 10502 19071
rect 10554 19019 10610 19071
rect 10662 19019 10718 19071
rect 10770 19019 10826 19071
rect 10878 19019 10934 19071
rect 10986 19019 11042 19071
rect 11094 19019 11150 19071
rect 11202 19019 11229 19071
rect 9179 18629 11229 19019
rect 9179 18577 9206 18629
rect 9258 18577 9314 18629
rect 9366 18577 9422 18629
rect 9474 18577 9530 18629
rect 9582 18577 9638 18629
rect 9690 18577 9746 18629
rect 9798 18577 9854 18629
rect 9906 18577 9962 18629
rect 10014 18577 10070 18629
rect 10122 18577 10178 18629
rect 10230 18577 10286 18629
rect 10338 18577 10394 18629
rect 10446 18577 10502 18629
rect 10554 18577 10610 18629
rect 10662 18577 10718 18629
rect 10770 18577 10826 18629
rect 10878 18577 10934 18629
rect 10986 18577 11042 18629
rect 11094 18577 11150 18629
rect 11202 18577 11229 18629
rect 9179 18521 11229 18577
rect 9179 18469 9206 18521
rect 9258 18469 9314 18521
rect 9366 18469 9422 18521
rect 9474 18469 9530 18521
rect 9582 18469 9638 18521
rect 9690 18469 9746 18521
rect 9798 18469 9854 18521
rect 9906 18469 9962 18521
rect 10014 18469 10070 18521
rect 10122 18469 10178 18521
rect 10230 18469 10286 18521
rect 10338 18469 10394 18521
rect 10446 18469 10502 18521
rect 10554 18469 10610 18521
rect 10662 18469 10718 18521
rect 10770 18469 10826 18521
rect 10878 18469 10934 18521
rect 10986 18469 11042 18521
rect 11094 18469 11150 18521
rect 11202 18469 11229 18521
rect 9179 18079 11229 18469
rect 9179 18027 9206 18079
rect 9258 18027 9314 18079
rect 9366 18027 9422 18079
rect 9474 18027 9530 18079
rect 9582 18027 9638 18079
rect 9690 18027 9746 18079
rect 9798 18027 9854 18079
rect 9906 18027 9962 18079
rect 10014 18027 10070 18079
rect 10122 18027 10178 18079
rect 10230 18027 10286 18079
rect 10338 18027 10394 18079
rect 10446 18027 10502 18079
rect 10554 18027 10610 18079
rect 10662 18027 10718 18079
rect 10770 18027 10826 18079
rect 10878 18027 10934 18079
rect 10986 18027 11042 18079
rect 11094 18027 11150 18079
rect 11202 18027 11229 18079
rect 9179 17591 11229 18027
rect 9179 17539 9206 17591
rect 9258 17539 9314 17591
rect 9366 17539 9422 17591
rect 9474 17539 9530 17591
rect 9582 17539 9638 17591
rect 9690 17539 9746 17591
rect 9798 17539 9854 17591
rect 9906 17539 9962 17591
rect 10014 17539 10070 17591
rect 10122 17539 10178 17591
rect 10230 17539 10286 17591
rect 10338 17539 10394 17591
rect 10446 17539 10502 17591
rect 10554 17539 10610 17591
rect 10662 17539 10718 17591
rect 10770 17539 10826 17591
rect 10878 17539 10934 17591
rect 10986 17539 11042 17591
rect 11094 17539 11150 17591
rect 11202 17539 11229 17591
rect 9179 17103 11229 17539
rect 9179 17051 9206 17103
rect 9258 17051 9314 17103
rect 9366 17051 9422 17103
rect 9474 17051 9530 17103
rect 9582 17051 9638 17103
rect 9690 17051 9746 17103
rect 9798 17051 9854 17103
rect 9906 17051 9962 17103
rect 10014 17051 10070 17103
rect 10122 17051 10178 17103
rect 10230 17051 10286 17103
rect 10338 17051 10394 17103
rect 10446 17051 10502 17103
rect 10554 17051 10610 17103
rect 10662 17051 10718 17103
rect 10770 17051 10826 17103
rect 10878 17051 10934 17103
rect 10986 17051 11042 17103
rect 11094 17051 11150 17103
rect 11202 17051 11229 17103
rect 9179 16615 11229 17051
rect 9179 16563 9206 16615
rect 9258 16563 9314 16615
rect 9366 16563 9422 16615
rect 9474 16563 9530 16615
rect 9582 16563 9638 16615
rect 9690 16563 9746 16615
rect 9798 16563 9854 16615
rect 9906 16563 9962 16615
rect 10014 16563 10070 16615
rect 10122 16563 10178 16615
rect 10230 16563 10286 16615
rect 10338 16563 10394 16615
rect 10446 16563 10502 16615
rect 10554 16563 10610 16615
rect 10662 16563 10718 16615
rect 10770 16563 10826 16615
rect 10878 16563 10934 16615
rect 10986 16563 11042 16615
rect 11094 16563 11150 16615
rect 11202 16563 11229 16615
rect 9179 16127 11229 16563
rect 9179 16075 9206 16127
rect 9258 16075 9314 16127
rect 9366 16075 9422 16127
rect 9474 16075 9530 16127
rect 9582 16075 9638 16127
rect 9690 16075 9746 16127
rect 9798 16075 9854 16127
rect 9906 16075 9962 16127
rect 10014 16075 10070 16127
rect 10122 16075 10178 16127
rect 10230 16075 10286 16127
rect 10338 16075 10394 16127
rect 10446 16075 10502 16127
rect 10554 16075 10610 16127
rect 10662 16075 10718 16127
rect 10770 16075 10826 16127
rect 10878 16075 10934 16127
rect 10986 16075 11042 16127
rect 11094 16075 11150 16127
rect 11202 16075 11229 16127
rect 9179 15639 11229 16075
rect 9179 15587 9206 15639
rect 9258 15587 9314 15639
rect 9366 15587 9422 15639
rect 9474 15587 9530 15639
rect 9582 15587 9638 15639
rect 9690 15587 9746 15639
rect 9798 15587 9854 15639
rect 9906 15587 9962 15639
rect 10014 15587 10070 15639
rect 10122 15587 10178 15639
rect 10230 15587 10286 15639
rect 10338 15587 10394 15639
rect 10446 15587 10502 15639
rect 10554 15587 10610 15639
rect 10662 15587 10718 15639
rect 10770 15587 10826 15639
rect 10878 15587 10934 15639
rect 10986 15587 11042 15639
rect 11094 15587 11150 15639
rect 11202 15587 11229 15639
rect 9179 15151 11229 15587
rect 9179 15099 9206 15151
rect 9258 15099 9314 15151
rect 9366 15099 9422 15151
rect 9474 15099 9530 15151
rect 9582 15099 9638 15151
rect 9690 15099 9746 15151
rect 9798 15099 9854 15151
rect 9906 15099 9962 15151
rect 10014 15099 10070 15151
rect 10122 15099 10178 15151
rect 10230 15099 10286 15151
rect 10338 15099 10394 15151
rect 10446 15099 10502 15151
rect 10554 15099 10610 15151
rect 10662 15099 10718 15151
rect 10770 15099 10826 15151
rect 10878 15099 10934 15151
rect 10986 15099 11042 15151
rect 11094 15099 11150 15151
rect 11202 15099 11229 15151
rect 9179 14663 11229 15099
rect 9179 14611 9206 14663
rect 9258 14611 9314 14663
rect 9366 14611 9422 14663
rect 9474 14611 9530 14663
rect 9582 14611 9638 14663
rect 9690 14611 9746 14663
rect 9798 14611 9854 14663
rect 9906 14611 9962 14663
rect 10014 14611 10070 14663
rect 10122 14611 10178 14663
rect 10230 14611 10286 14663
rect 10338 14611 10394 14663
rect 10446 14611 10502 14663
rect 10554 14611 10610 14663
rect 10662 14611 10718 14663
rect 10770 14611 10826 14663
rect 10878 14611 10934 14663
rect 10986 14611 11042 14663
rect 11094 14611 11150 14663
rect 11202 14611 11229 14663
rect 9179 14175 11229 14611
rect 9179 14123 9206 14175
rect 9258 14123 9314 14175
rect 9366 14123 9422 14175
rect 9474 14123 9530 14175
rect 9582 14123 9638 14175
rect 9690 14123 9746 14175
rect 9798 14123 9854 14175
rect 9906 14123 9962 14175
rect 10014 14123 10070 14175
rect 10122 14123 10178 14175
rect 10230 14123 10286 14175
rect 10338 14123 10394 14175
rect 10446 14123 10502 14175
rect 10554 14123 10610 14175
rect 10662 14123 10718 14175
rect 10770 14123 10826 14175
rect 10878 14123 10934 14175
rect 10986 14123 11042 14175
rect 11094 14123 11150 14175
rect 11202 14123 11229 14175
rect 9179 13687 11229 14123
rect 9179 13635 9206 13687
rect 9258 13635 9314 13687
rect 9366 13635 9422 13687
rect 9474 13635 9530 13687
rect 9582 13635 9638 13687
rect 9690 13635 9746 13687
rect 9798 13635 9854 13687
rect 9906 13635 9962 13687
rect 10014 13635 10070 13687
rect 10122 13635 10178 13687
rect 10230 13635 10286 13687
rect 10338 13635 10394 13687
rect 10446 13635 10502 13687
rect 10554 13635 10610 13687
rect 10662 13635 10718 13687
rect 10770 13635 10826 13687
rect 10878 13635 10934 13687
rect 10986 13635 11042 13687
rect 11094 13635 11150 13687
rect 11202 13635 11229 13687
rect 9179 13199 11229 13635
rect 9179 13147 9206 13199
rect 9258 13147 9314 13199
rect 9366 13147 9422 13199
rect 9474 13147 9530 13199
rect 9582 13147 9638 13199
rect 9690 13147 9746 13199
rect 9798 13147 9854 13199
rect 9906 13147 9962 13199
rect 10014 13147 10070 13199
rect 10122 13147 10178 13199
rect 10230 13147 10286 13199
rect 10338 13147 10394 13199
rect 10446 13147 10502 13199
rect 10554 13147 10610 13199
rect 10662 13147 10718 13199
rect 10770 13147 10826 13199
rect 10878 13147 10934 13199
rect 10986 13147 11042 13199
rect 11094 13147 11150 13199
rect 11202 13147 11229 13199
rect 9179 12757 11229 13147
rect 9179 12705 9206 12757
rect 9258 12705 9314 12757
rect 9366 12705 9422 12757
rect 9474 12705 9530 12757
rect 9582 12705 9638 12757
rect 9690 12705 9746 12757
rect 9798 12705 9854 12757
rect 9906 12705 9962 12757
rect 10014 12705 10070 12757
rect 10122 12705 10178 12757
rect 10230 12705 10286 12757
rect 10338 12705 10394 12757
rect 10446 12705 10502 12757
rect 10554 12705 10610 12757
rect 10662 12705 10718 12757
rect 10770 12705 10826 12757
rect 10878 12705 10934 12757
rect 10986 12705 11042 12757
rect 11094 12705 11150 12757
rect 11202 12705 11229 12757
rect 9179 12649 11229 12705
rect 9179 12597 9206 12649
rect 9258 12597 9314 12649
rect 9366 12597 9422 12649
rect 9474 12597 9530 12649
rect 9582 12597 9638 12649
rect 9690 12597 9746 12649
rect 9798 12597 9854 12649
rect 9906 12597 9962 12649
rect 10014 12597 10070 12649
rect 10122 12597 10178 12649
rect 10230 12597 10286 12649
rect 10338 12597 10394 12649
rect 10446 12597 10502 12649
rect 10554 12597 10610 12649
rect 10662 12597 10718 12649
rect 10770 12597 10826 12649
rect 10878 12597 10934 12649
rect 10986 12597 11042 12649
rect 11094 12597 11150 12649
rect 11202 12597 11229 12649
rect 9179 12207 11229 12597
rect 9179 12155 9206 12207
rect 9258 12155 9314 12207
rect 9366 12155 9422 12207
rect 9474 12155 9530 12207
rect 9582 12155 9638 12207
rect 9690 12155 9746 12207
rect 9798 12155 9854 12207
rect 9906 12155 9962 12207
rect 10014 12155 10070 12207
rect 10122 12155 10178 12207
rect 10230 12155 10286 12207
rect 10338 12155 10394 12207
rect 10446 12155 10502 12207
rect 10554 12155 10610 12207
rect 10662 12155 10718 12207
rect 10770 12155 10826 12207
rect 10878 12155 10934 12207
rect 10986 12155 11042 12207
rect 11094 12155 11150 12207
rect 11202 12155 11229 12207
rect 9179 11719 11229 12155
rect 9179 11667 9206 11719
rect 9258 11667 9314 11719
rect 9366 11667 9422 11719
rect 9474 11667 9530 11719
rect 9582 11667 9638 11719
rect 9690 11667 9746 11719
rect 9798 11667 9854 11719
rect 9906 11667 9962 11719
rect 10014 11667 10070 11719
rect 10122 11667 10178 11719
rect 10230 11667 10286 11719
rect 10338 11667 10394 11719
rect 10446 11667 10502 11719
rect 10554 11667 10610 11719
rect 10662 11667 10718 11719
rect 10770 11667 10826 11719
rect 10878 11667 10934 11719
rect 10986 11667 11042 11719
rect 11094 11667 11150 11719
rect 11202 11667 11229 11719
rect 9179 11231 11229 11667
rect 9179 11179 9206 11231
rect 9258 11179 9314 11231
rect 9366 11179 9422 11231
rect 9474 11179 9530 11231
rect 9582 11179 9638 11231
rect 9690 11179 9746 11231
rect 9798 11179 9854 11231
rect 9906 11179 9962 11231
rect 10014 11179 10070 11231
rect 10122 11179 10178 11231
rect 10230 11179 10286 11231
rect 10338 11179 10394 11231
rect 10446 11179 10502 11231
rect 10554 11179 10610 11231
rect 10662 11179 10718 11231
rect 10770 11179 10826 11231
rect 10878 11179 10934 11231
rect 10986 11179 11042 11231
rect 11094 11179 11150 11231
rect 11202 11179 11229 11231
rect 9179 10743 11229 11179
rect 9179 10691 9206 10743
rect 9258 10691 9314 10743
rect 9366 10691 9422 10743
rect 9474 10691 9530 10743
rect 9582 10691 9638 10743
rect 9690 10691 9746 10743
rect 9798 10691 9854 10743
rect 9906 10691 9962 10743
rect 10014 10691 10070 10743
rect 10122 10691 10178 10743
rect 10230 10691 10286 10743
rect 10338 10691 10394 10743
rect 10446 10691 10502 10743
rect 10554 10691 10610 10743
rect 10662 10691 10718 10743
rect 10770 10691 10826 10743
rect 10878 10691 10934 10743
rect 10986 10691 11042 10743
rect 11094 10691 11150 10743
rect 11202 10691 11229 10743
rect 9179 10255 11229 10691
rect 9179 10203 9206 10255
rect 9258 10203 9314 10255
rect 9366 10203 9422 10255
rect 9474 10203 9530 10255
rect 9582 10203 9638 10255
rect 9690 10203 9746 10255
rect 9798 10203 9854 10255
rect 9906 10203 9962 10255
rect 10014 10203 10070 10255
rect 10122 10203 10178 10255
rect 10230 10203 10286 10255
rect 10338 10203 10394 10255
rect 10446 10203 10502 10255
rect 10554 10203 10610 10255
rect 10662 10203 10718 10255
rect 10770 10203 10826 10255
rect 10878 10203 10934 10255
rect 10986 10203 11042 10255
rect 11094 10203 11150 10255
rect 11202 10203 11229 10255
rect 9179 9767 11229 10203
rect 9179 9715 9206 9767
rect 9258 9715 9314 9767
rect 9366 9715 9422 9767
rect 9474 9715 9530 9767
rect 9582 9715 9638 9767
rect 9690 9715 9746 9767
rect 9798 9715 9854 9767
rect 9906 9715 9962 9767
rect 10014 9715 10070 9767
rect 10122 9715 10178 9767
rect 10230 9715 10286 9767
rect 10338 9715 10394 9767
rect 10446 9715 10502 9767
rect 10554 9715 10610 9767
rect 10662 9715 10718 9767
rect 10770 9715 10826 9767
rect 10878 9715 10934 9767
rect 10986 9715 11042 9767
rect 11094 9715 11150 9767
rect 11202 9715 11229 9767
rect 9179 9279 11229 9715
rect 9179 9227 9206 9279
rect 9258 9227 9314 9279
rect 9366 9227 9422 9279
rect 9474 9227 9530 9279
rect 9582 9227 9638 9279
rect 9690 9227 9746 9279
rect 9798 9227 9854 9279
rect 9906 9227 9962 9279
rect 10014 9227 10070 9279
rect 10122 9227 10178 9279
rect 10230 9227 10286 9279
rect 10338 9227 10394 9279
rect 10446 9227 10502 9279
rect 10554 9227 10610 9279
rect 10662 9227 10718 9279
rect 10770 9227 10826 9279
rect 10878 9227 10934 9279
rect 10986 9227 11042 9279
rect 11094 9227 11150 9279
rect 11202 9227 11229 9279
rect 9179 8791 11229 9227
rect 9179 8739 9206 8791
rect 9258 8739 9314 8791
rect 9366 8739 9422 8791
rect 9474 8739 9530 8791
rect 9582 8739 9638 8791
rect 9690 8739 9746 8791
rect 9798 8739 9854 8791
rect 9906 8739 9962 8791
rect 10014 8739 10070 8791
rect 10122 8739 10178 8791
rect 10230 8739 10286 8791
rect 10338 8739 10394 8791
rect 10446 8739 10502 8791
rect 10554 8739 10610 8791
rect 10662 8739 10718 8791
rect 10770 8739 10826 8791
rect 10878 8739 10934 8791
rect 10986 8739 11042 8791
rect 11094 8739 11150 8791
rect 11202 8739 11229 8791
rect 9179 8303 11229 8739
rect 9179 8251 9206 8303
rect 9258 8251 9314 8303
rect 9366 8251 9422 8303
rect 9474 8251 9530 8303
rect 9582 8251 9638 8303
rect 9690 8251 9746 8303
rect 9798 8251 9854 8303
rect 9906 8251 9962 8303
rect 10014 8251 10070 8303
rect 10122 8251 10178 8303
rect 10230 8251 10286 8303
rect 10338 8251 10394 8303
rect 10446 8251 10502 8303
rect 10554 8251 10610 8303
rect 10662 8251 10718 8303
rect 10770 8251 10826 8303
rect 10878 8251 10934 8303
rect 10986 8251 11042 8303
rect 11094 8251 11150 8303
rect 11202 8251 11229 8303
rect 9179 7815 11229 8251
rect 9179 7763 9206 7815
rect 9258 7763 9314 7815
rect 9366 7763 9422 7815
rect 9474 7763 9530 7815
rect 9582 7763 9638 7815
rect 9690 7763 9746 7815
rect 9798 7763 9854 7815
rect 9906 7763 9962 7815
rect 10014 7763 10070 7815
rect 10122 7763 10178 7815
rect 10230 7763 10286 7815
rect 10338 7763 10394 7815
rect 10446 7763 10502 7815
rect 10554 7763 10610 7815
rect 10662 7763 10718 7815
rect 10770 7763 10826 7815
rect 10878 7763 10934 7815
rect 10986 7763 11042 7815
rect 11094 7763 11150 7815
rect 11202 7763 11229 7815
rect 9179 7327 11229 7763
rect 9179 7275 9206 7327
rect 9258 7275 9314 7327
rect 9366 7275 9422 7327
rect 9474 7275 9530 7327
rect 9582 7275 9638 7327
rect 9690 7275 9746 7327
rect 9798 7275 9854 7327
rect 9906 7275 9962 7327
rect 10014 7275 10070 7327
rect 10122 7275 10178 7327
rect 10230 7275 10286 7327
rect 10338 7275 10394 7327
rect 10446 7275 10502 7327
rect 10554 7275 10610 7327
rect 10662 7275 10718 7327
rect 10770 7275 10826 7327
rect 10878 7275 10934 7327
rect 10986 7275 11042 7327
rect 11094 7275 11150 7327
rect 11202 7275 11229 7327
rect 9179 6885 11229 7275
rect 9179 6833 9206 6885
rect 9258 6833 9314 6885
rect 9366 6833 9422 6885
rect 9474 6833 9530 6885
rect 9582 6833 9638 6885
rect 9690 6833 9746 6885
rect 9798 6833 9854 6885
rect 9906 6833 9962 6885
rect 10014 6833 10070 6885
rect 10122 6833 10178 6885
rect 10230 6833 10286 6885
rect 10338 6833 10394 6885
rect 10446 6833 10502 6885
rect 10554 6833 10610 6885
rect 10662 6833 10718 6885
rect 10770 6833 10826 6885
rect 10878 6833 10934 6885
rect 10986 6833 11042 6885
rect 11094 6833 11150 6885
rect 11202 6833 11229 6885
rect 9179 6777 11229 6833
rect 9179 6725 9206 6777
rect 9258 6725 9314 6777
rect 9366 6725 9422 6777
rect 9474 6725 9530 6777
rect 9582 6725 9638 6777
rect 9690 6725 9746 6777
rect 9798 6725 9854 6777
rect 9906 6725 9962 6777
rect 10014 6725 10070 6777
rect 10122 6725 10178 6777
rect 10230 6725 10286 6777
rect 10338 6725 10394 6777
rect 10446 6725 10502 6777
rect 10554 6725 10610 6777
rect 10662 6725 10718 6777
rect 10770 6725 10826 6777
rect 10878 6725 10934 6777
rect 10986 6725 11042 6777
rect 11094 6725 11150 6777
rect 11202 6725 11229 6777
rect 9179 6335 11229 6725
rect 9179 6283 9206 6335
rect 9258 6283 9314 6335
rect 9366 6283 9422 6335
rect 9474 6283 9530 6335
rect 9582 6283 9638 6335
rect 9690 6283 9746 6335
rect 9798 6283 9854 6335
rect 9906 6283 9962 6335
rect 10014 6283 10070 6335
rect 10122 6283 10178 6335
rect 10230 6283 10286 6335
rect 10338 6283 10394 6335
rect 10446 6283 10502 6335
rect 10554 6283 10610 6335
rect 10662 6283 10718 6335
rect 10770 6283 10826 6335
rect 10878 6283 10934 6335
rect 10986 6283 11042 6335
rect 11094 6283 11150 6335
rect 11202 6283 11229 6335
rect 9179 5847 11229 6283
rect 9179 5795 9206 5847
rect 9258 5795 9314 5847
rect 9366 5795 9422 5847
rect 9474 5795 9530 5847
rect 9582 5795 9638 5847
rect 9690 5795 9746 5847
rect 9798 5795 9854 5847
rect 9906 5795 9962 5847
rect 10014 5795 10070 5847
rect 10122 5795 10178 5847
rect 10230 5795 10286 5847
rect 10338 5795 10394 5847
rect 10446 5795 10502 5847
rect 10554 5795 10610 5847
rect 10662 5795 10718 5847
rect 10770 5795 10826 5847
rect 10878 5795 10934 5847
rect 10986 5795 11042 5847
rect 11094 5795 11150 5847
rect 11202 5795 11229 5847
rect 9179 5359 11229 5795
rect 9179 5307 9206 5359
rect 9258 5307 9314 5359
rect 9366 5307 9422 5359
rect 9474 5307 9530 5359
rect 9582 5307 9638 5359
rect 9690 5307 9746 5359
rect 9798 5307 9854 5359
rect 9906 5307 9962 5359
rect 10014 5307 10070 5359
rect 10122 5307 10178 5359
rect 10230 5307 10286 5359
rect 10338 5307 10394 5359
rect 10446 5307 10502 5359
rect 10554 5307 10610 5359
rect 10662 5307 10718 5359
rect 10770 5307 10826 5359
rect 10878 5307 10934 5359
rect 10986 5307 11042 5359
rect 11094 5307 11150 5359
rect 11202 5307 11229 5359
rect 9179 4871 11229 5307
rect 9179 4819 9206 4871
rect 9258 4819 9314 4871
rect 9366 4819 9422 4871
rect 9474 4819 9530 4871
rect 9582 4819 9638 4871
rect 9690 4819 9746 4871
rect 9798 4819 9854 4871
rect 9906 4819 9962 4871
rect 10014 4819 10070 4871
rect 10122 4819 10178 4871
rect 10230 4819 10286 4871
rect 10338 4819 10394 4871
rect 10446 4819 10502 4871
rect 10554 4819 10610 4871
rect 10662 4819 10718 4871
rect 10770 4819 10826 4871
rect 10878 4819 10934 4871
rect 10986 4819 11042 4871
rect 11094 4819 11150 4871
rect 11202 4819 11229 4871
rect 9179 4383 11229 4819
rect 9179 4331 9206 4383
rect 9258 4331 9314 4383
rect 9366 4331 9422 4383
rect 9474 4331 9530 4383
rect 9582 4331 9638 4383
rect 9690 4331 9746 4383
rect 9798 4331 9854 4383
rect 9906 4331 9962 4383
rect 10014 4331 10070 4383
rect 10122 4331 10178 4383
rect 10230 4331 10286 4383
rect 10338 4331 10394 4383
rect 10446 4331 10502 4383
rect 10554 4331 10610 4383
rect 10662 4331 10718 4383
rect 10770 4331 10826 4383
rect 10878 4331 10934 4383
rect 10986 4331 11042 4383
rect 11094 4331 11150 4383
rect 11202 4331 11229 4383
rect 9179 3895 11229 4331
rect 9179 3843 9206 3895
rect 9258 3843 9314 3895
rect 9366 3843 9422 3895
rect 9474 3843 9530 3895
rect 9582 3843 9638 3895
rect 9690 3843 9746 3895
rect 9798 3843 9854 3895
rect 9906 3843 9962 3895
rect 10014 3843 10070 3895
rect 10122 3843 10178 3895
rect 10230 3843 10286 3895
rect 10338 3843 10394 3895
rect 10446 3843 10502 3895
rect 10554 3843 10610 3895
rect 10662 3843 10718 3895
rect 10770 3843 10826 3895
rect 10878 3843 10934 3895
rect 10986 3843 11042 3895
rect 11094 3843 11150 3895
rect 11202 3843 11229 3895
rect 9179 3407 11229 3843
rect 9179 3355 9206 3407
rect 9258 3355 9314 3407
rect 9366 3355 9422 3407
rect 9474 3355 9530 3407
rect 9582 3355 9638 3407
rect 9690 3355 9746 3407
rect 9798 3355 9854 3407
rect 9906 3355 9962 3407
rect 10014 3355 10070 3407
rect 10122 3355 10178 3407
rect 10230 3355 10286 3407
rect 10338 3355 10394 3407
rect 10446 3355 10502 3407
rect 10554 3355 10610 3407
rect 10662 3355 10718 3407
rect 10770 3355 10826 3407
rect 10878 3355 10934 3407
rect 10986 3355 11042 3407
rect 11094 3355 11150 3407
rect 11202 3355 11229 3407
rect 9179 2919 11229 3355
rect 9179 2867 9206 2919
rect 9258 2867 9314 2919
rect 9366 2867 9422 2919
rect 9474 2867 9530 2919
rect 9582 2867 9638 2919
rect 9690 2867 9746 2919
rect 9798 2867 9854 2919
rect 9906 2867 9962 2919
rect 10014 2867 10070 2919
rect 10122 2867 10178 2919
rect 10230 2867 10286 2919
rect 10338 2867 10394 2919
rect 10446 2867 10502 2919
rect 10554 2867 10610 2919
rect 10662 2867 10718 2919
rect 10770 2867 10826 2919
rect 10878 2867 10934 2919
rect 10986 2867 11042 2919
rect 11094 2867 11150 2919
rect 11202 2867 11229 2919
rect 9179 2431 11229 2867
rect 9179 2379 9206 2431
rect 9258 2379 9314 2431
rect 9366 2379 9422 2431
rect 9474 2379 9530 2431
rect 9582 2379 9638 2431
rect 9690 2379 9746 2431
rect 9798 2379 9854 2431
rect 9906 2379 9962 2431
rect 10014 2379 10070 2431
rect 10122 2379 10178 2431
rect 10230 2379 10286 2431
rect 10338 2379 10394 2431
rect 10446 2379 10502 2431
rect 10554 2379 10610 2431
rect 10662 2379 10718 2431
rect 10770 2379 10826 2431
rect 10878 2379 10934 2431
rect 10986 2379 11042 2431
rect 11094 2379 11150 2431
rect 11202 2379 11229 2431
rect 9179 1943 11229 2379
rect 9179 1891 9206 1943
rect 9258 1891 9314 1943
rect 9366 1891 9422 1943
rect 9474 1891 9530 1943
rect 9582 1891 9638 1943
rect 9690 1891 9746 1943
rect 9798 1891 9854 1943
rect 9906 1891 9962 1943
rect 10014 1891 10070 1943
rect 10122 1891 10178 1943
rect 10230 1891 10286 1943
rect 10338 1891 10394 1943
rect 10446 1891 10502 1943
rect 10554 1891 10610 1943
rect 10662 1891 10718 1943
rect 10770 1891 10826 1943
rect 10878 1891 10934 1943
rect 10986 1891 11042 1943
rect 11094 1891 11150 1943
rect 11202 1891 11229 1943
rect 9179 1455 11229 1891
rect 9179 1403 9206 1455
rect 9258 1403 9314 1455
rect 9366 1403 9422 1455
rect 9474 1403 9530 1455
rect 9582 1403 9638 1455
rect 9690 1403 9746 1455
rect 9798 1403 9854 1455
rect 9906 1403 9962 1455
rect 10014 1403 10070 1455
rect 10122 1403 10178 1455
rect 10230 1403 10286 1455
rect 10338 1403 10394 1455
rect 10446 1403 10502 1455
rect 10554 1403 10610 1455
rect 10662 1403 10718 1455
rect 10770 1403 10826 1455
rect 10878 1403 10934 1455
rect 10986 1403 11042 1455
rect 11094 1403 11150 1455
rect 11202 1403 11229 1455
rect 9179 961 11229 1403
rect 9179 909 9206 961
rect 9258 909 9314 961
rect 9366 909 9422 961
rect 9474 909 9530 961
rect 9582 909 9638 961
rect 9690 909 9746 961
rect 9798 909 9854 961
rect 9906 909 9962 961
rect 10014 909 10070 961
rect 10122 909 10178 961
rect 10230 909 10286 961
rect 10338 909 10394 961
rect 10446 909 10502 961
rect 10554 909 10610 961
rect 10662 909 10718 961
rect 10770 909 10826 961
rect 10878 909 10934 961
rect 10986 909 11042 961
rect 11094 909 11150 961
rect 11202 909 11229 961
rect 9179 853 11229 909
rect 9179 801 9206 853
rect 9258 801 9314 853
rect 9366 801 9422 853
rect 9474 801 9530 853
rect 9582 801 9638 853
rect 9690 801 9746 853
rect 9798 801 9854 853
rect 9906 801 9962 853
rect 10014 801 10070 853
rect 10122 801 10178 853
rect 10230 801 10286 853
rect 10338 801 10394 853
rect 10446 801 10502 853
rect 10554 801 10610 853
rect 10662 801 10718 853
rect 10770 801 10826 853
rect 10878 801 10934 853
rect 10986 801 11042 853
rect 11094 801 11150 853
rect 11202 801 11229 853
rect 9179 745 11229 801
rect 9179 693 9206 745
rect 9258 693 9314 745
rect 9366 693 9422 745
rect 9474 693 9530 745
rect 9582 693 9638 745
rect 9690 693 9746 745
rect 9798 693 9854 745
rect 9906 693 9962 745
rect 10014 693 10070 745
rect 10122 693 10178 745
rect 10230 693 10286 745
rect 10338 693 10394 745
rect 10446 693 10502 745
rect 10554 693 10610 745
rect 10662 693 10718 745
rect 10770 693 10826 745
rect 10878 693 10934 745
rect 10986 693 11042 745
rect 11094 693 11150 745
rect 11202 693 11229 745
rect 9179 43 11229 693
rect 11289 25261 11489 25617
rect 11289 25209 11309 25261
rect 11361 25209 11417 25261
rect 11469 25209 11489 25261
rect 11289 25153 11489 25209
rect 11289 25101 11309 25153
rect 11361 25101 11417 25153
rect 11469 25101 11489 25153
rect 11289 25045 11489 25101
rect 11289 24993 11309 25045
rect 11361 24993 11417 25045
rect 11469 24993 11489 25045
rect 11289 23707 11489 24993
rect 11289 23655 11309 23707
rect 11361 23655 11417 23707
rect 11469 23655 11489 23707
rect 11289 23219 11489 23655
rect 11289 23167 11309 23219
rect 11361 23167 11417 23219
rect 11469 23167 11489 23219
rect 11289 22731 11489 23167
rect 11289 22679 11309 22731
rect 11361 22679 11417 22731
rect 11469 22679 11489 22731
rect 11289 22243 11489 22679
rect 11289 22191 11309 22243
rect 11361 22191 11417 22243
rect 11469 22191 11489 22243
rect 11289 21755 11489 22191
rect 11289 21703 11309 21755
rect 11361 21703 11417 21755
rect 11469 21703 11489 21755
rect 11289 21267 11489 21703
rect 11289 21215 11309 21267
rect 11361 21215 11417 21267
rect 11469 21215 11489 21267
rect 11289 20779 11489 21215
rect 11289 20727 11309 20779
rect 11361 20727 11417 20779
rect 11469 20727 11489 20779
rect 11289 20291 11489 20727
rect 11289 20239 11309 20291
rect 11361 20239 11417 20291
rect 11469 20239 11489 20291
rect 11289 19803 11489 20239
rect 11289 19751 11309 19803
rect 11361 19751 11417 19803
rect 11469 19751 11489 19803
rect 11289 19315 11489 19751
rect 11289 19263 11309 19315
rect 11361 19263 11417 19315
rect 11469 19263 11489 19315
rect 11289 17835 11489 19263
rect 11289 17783 11309 17835
rect 11361 17783 11417 17835
rect 11469 17783 11489 17835
rect 11289 17347 11489 17783
rect 11289 17295 11309 17347
rect 11361 17295 11417 17347
rect 11469 17295 11489 17347
rect 11289 16859 11489 17295
rect 11289 16807 11309 16859
rect 11361 16807 11417 16859
rect 11469 16807 11489 16859
rect 11289 16371 11489 16807
rect 11289 16319 11309 16371
rect 11361 16319 11417 16371
rect 11469 16319 11489 16371
rect 11289 15883 11489 16319
rect 11289 15831 11309 15883
rect 11361 15831 11417 15883
rect 11469 15831 11489 15883
rect 11289 15395 11489 15831
rect 11289 15343 11309 15395
rect 11361 15343 11417 15395
rect 11469 15343 11489 15395
rect 11289 14907 11489 15343
rect 11289 14855 11309 14907
rect 11361 14855 11417 14907
rect 11469 14855 11489 14907
rect 11289 14419 11489 14855
rect 11289 14367 11309 14419
rect 11361 14367 11417 14419
rect 11469 14367 11489 14419
rect 11289 13931 11489 14367
rect 11289 13879 11309 13931
rect 11361 13879 11417 13931
rect 11469 13879 11489 13931
rect 11289 13443 11489 13879
rect 11289 13391 11309 13443
rect 11361 13391 11417 13443
rect 11469 13391 11489 13443
rect 11289 11963 11489 13391
rect 11289 11911 11309 11963
rect 11361 11911 11417 11963
rect 11469 11911 11489 11963
rect 11289 11475 11489 11911
rect 11289 11423 11309 11475
rect 11361 11423 11417 11475
rect 11469 11423 11489 11475
rect 11289 10987 11489 11423
rect 11289 10935 11309 10987
rect 11361 10935 11417 10987
rect 11469 10935 11489 10987
rect 11289 10499 11489 10935
rect 11289 10447 11309 10499
rect 11361 10447 11417 10499
rect 11469 10447 11489 10499
rect 11289 10011 11489 10447
rect 11289 9959 11309 10011
rect 11361 9959 11417 10011
rect 11469 9959 11489 10011
rect 11289 9523 11489 9959
rect 11289 9471 11309 9523
rect 11361 9471 11417 9523
rect 11469 9471 11489 9523
rect 11289 9035 11489 9471
rect 11289 8983 11309 9035
rect 11361 8983 11417 9035
rect 11469 8983 11489 9035
rect 11289 8547 11489 8983
rect 11289 8495 11309 8547
rect 11361 8495 11417 8547
rect 11469 8495 11489 8547
rect 11289 8059 11489 8495
rect 11289 8007 11309 8059
rect 11361 8007 11417 8059
rect 11469 8007 11489 8059
rect 11289 7571 11489 8007
rect 11289 7519 11309 7571
rect 11361 7519 11417 7571
rect 11469 7519 11489 7571
rect 11289 6091 11489 7519
rect 11289 6039 11309 6091
rect 11361 6039 11417 6091
rect 11469 6039 11489 6091
rect 11289 5603 11489 6039
rect 11289 5551 11309 5603
rect 11361 5551 11417 5603
rect 11469 5551 11489 5603
rect 11289 5115 11489 5551
rect 11289 5063 11309 5115
rect 11361 5063 11417 5115
rect 11469 5063 11489 5115
rect 11289 4627 11489 5063
rect 11289 4575 11309 4627
rect 11361 4575 11417 4627
rect 11469 4575 11489 4627
rect 11289 4139 11489 4575
rect 11289 4087 11309 4139
rect 11361 4087 11417 4139
rect 11469 4087 11489 4139
rect 11289 3651 11489 4087
rect 11289 3599 11309 3651
rect 11361 3599 11417 3651
rect 11469 3599 11489 3651
rect 11289 3163 11489 3599
rect 11289 3111 11309 3163
rect 11361 3111 11417 3163
rect 11469 3111 11489 3163
rect 11289 2675 11489 3111
rect 11289 2623 11309 2675
rect 11361 2623 11417 2675
rect 11469 2623 11489 2675
rect 11289 2187 11489 2623
rect 11289 2135 11309 2187
rect 11361 2135 11417 2187
rect 11469 2135 11489 2187
rect 11289 1699 11489 2135
rect 11289 1647 11309 1699
rect 11361 1647 11417 1699
rect 11469 1647 11489 1699
rect 11289 361 11489 1647
rect 11549 23887 11749 25617
rect 11549 23835 11569 23887
rect 11621 23835 11677 23887
rect 11729 23835 11749 23887
rect 11549 23779 11749 23835
rect 11549 23727 11569 23779
rect 11621 23727 11677 23779
rect 11729 23727 11749 23779
rect 11549 23671 11749 23727
rect 11549 23619 11569 23671
rect 11621 23619 11677 23671
rect 11729 23619 11749 23671
rect 11549 23563 11749 23619
rect 11549 23511 11569 23563
rect 11621 23511 11677 23563
rect 11729 23511 11749 23563
rect 11549 23455 11749 23511
rect 11549 23403 11569 23455
rect 11621 23403 11677 23455
rect 11729 23403 11749 23455
rect 11549 23347 11749 23403
rect 11549 23295 11569 23347
rect 11621 23295 11677 23347
rect 11729 23295 11749 23347
rect 11549 23239 11749 23295
rect 11549 23187 11569 23239
rect 11621 23187 11677 23239
rect 11729 23187 11749 23239
rect 11549 23131 11749 23187
rect 11549 23079 11569 23131
rect 11621 23079 11677 23131
rect 11729 23079 11749 23131
rect 11549 23023 11749 23079
rect 11549 22971 11569 23023
rect 11621 22971 11677 23023
rect 11729 22971 11749 23023
rect 11549 22915 11749 22971
rect 11549 22863 11569 22915
rect 11621 22863 11677 22915
rect 11729 22863 11749 22915
rect 11549 22807 11749 22863
rect 11549 22755 11569 22807
rect 11621 22755 11677 22807
rect 11729 22755 11749 22807
rect 11549 22699 11749 22755
rect 11549 22647 11569 22699
rect 11621 22647 11677 22699
rect 11729 22647 11749 22699
rect 11549 22591 11749 22647
rect 11549 22539 11569 22591
rect 11621 22539 11677 22591
rect 11729 22539 11749 22591
rect 11549 22483 11749 22539
rect 11549 22431 11569 22483
rect 11621 22431 11677 22483
rect 11729 22431 11749 22483
rect 11549 22375 11749 22431
rect 11549 22323 11569 22375
rect 11621 22323 11677 22375
rect 11729 22323 11749 22375
rect 11549 22267 11749 22323
rect 11549 22215 11569 22267
rect 11621 22215 11677 22267
rect 11729 22215 11749 22267
rect 11549 22159 11749 22215
rect 11549 22107 11569 22159
rect 11621 22107 11677 22159
rect 11729 22107 11749 22159
rect 11549 22051 11749 22107
rect 11549 21999 11569 22051
rect 11621 21999 11677 22051
rect 11729 21999 11749 22051
rect 11549 21943 11749 21999
rect 11549 21891 11569 21943
rect 11621 21891 11677 21943
rect 11729 21891 11749 21943
rect 11549 21835 11749 21891
rect 11549 21783 11569 21835
rect 11621 21783 11677 21835
rect 11729 21783 11749 21835
rect 11549 21727 11749 21783
rect 11549 21675 11569 21727
rect 11621 21675 11677 21727
rect 11729 21675 11749 21727
rect 11549 21619 11749 21675
rect 11549 21567 11569 21619
rect 11621 21567 11677 21619
rect 11729 21567 11749 21619
rect 11549 21511 11749 21567
rect 11549 21459 11569 21511
rect 11621 21459 11677 21511
rect 11729 21459 11749 21511
rect 11549 21403 11749 21459
rect 11549 21351 11569 21403
rect 11621 21351 11677 21403
rect 11729 21351 11749 21403
rect 11549 21295 11749 21351
rect 11549 21243 11569 21295
rect 11621 21243 11677 21295
rect 11729 21243 11749 21295
rect 11549 21187 11749 21243
rect 11549 21135 11569 21187
rect 11621 21135 11677 21187
rect 11729 21135 11749 21187
rect 11549 21079 11749 21135
rect 11549 21027 11569 21079
rect 11621 21027 11677 21079
rect 11729 21027 11749 21079
rect 11549 20971 11749 21027
rect 11549 20919 11569 20971
rect 11621 20919 11677 20971
rect 11729 20919 11749 20971
rect 11549 20863 11749 20919
rect 11549 20811 11569 20863
rect 11621 20811 11677 20863
rect 11729 20811 11749 20863
rect 11549 20755 11749 20811
rect 11549 20703 11569 20755
rect 11621 20703 11677 20755
rect 11729 20703 11749 20755
rect 11549 20647 11749 20703
rect 11549 20595 11569 20647
rect 11621 20595 11677 20647
rect 11729 20595 11749 20647
rect 11549 20539 11749 20595
rect 11549 20487 11569 20539
rect 11621 20487 11677 20539
rect 11729 20487 11749 20539
rect 11549 20431 11749 20487
rect 11549 20379 11569 20431
rect 11621 20379 11677 20431
rect 11729 20379 11749 20431
rect 11549 20323 11749 20379
rect 11549 20271 11569 20323
rect 11621 20271 11677 20323
rect 11729 20271 11749 20323
rect 11549 20215 11749 20271
rect 11549 20163 11569 20215
rect 11621 20163 11677 20215
rect 11729 20163 11749 20215
rect 11549 20107 11749 20163
rect 11549 20055 11569 20107
rect 11621 20055 11677 20107
rect 11729 20055 11749 20107
rect 11549 19999 11749 20055
rect 11549 19947 11569 19999
rect 11621 19947 11677 19999
rect 11729 19947 11749 19999
rect 11549 19891 11749 19947
rect 11549 19839 11569 19891
rect 11621 19839 11677 19891
rect 11729 19839 11749 19891
rect 11549 19783 11749 19839
rect 11549 19731 11569 19783
rect 11621 19731 11677 19783
rect 11729 19731 11749 19783
rect 11549 19675 11749 19731
rect 11549 19623 11569 19675
rect 11621 19623 11677 19675
rect 11729 19623 11749 19675
rect 11549 19567 11749 19623
rect 11549 19515 11569 19567
rect 11621 19515 11677 19567
rect 11729 19515 11749 19567
rect 11549 19459 11749 19515
rect 11549 19407 11569 19459
rect 11621 19407 11677 19459
rect 11729 19407 11749 19459
rect 11549 19351 11749 19407
rect 11549 19299 11569 19351
rect 11621 19299 11677 19351
rect 11729 19299 11749 19351
rect 11549 19243 11749 19299
rect 11549 19191 11569 19243
rect 11621 19191 11677 19243
rect 11729 19191 11749 19243
rect 11549 19135 11749 19191
rect 11549 19083 11569 19135
rect 11621 19083 11677 19135
rect 11729 19083 11749 19135
rect 11549 18015 11749 19083
rect 11549 17963 11569 18015
rect 11621 17963 11677 18015
rect 11729 17963 11749 18015
rect 11549 17907 11749 17963
rect 11549 17855 11569 17907
rect 11621 17855 11677 17907
rect 11729 17855 11749 17907
rect 11549 17799 11749 17855
rect 11549 17747 11569 17799
rect 11621 17747 11677 17799
rect 11729 17747 11749 17799
rect 11549 17691 11749 17747
rect 11549 17639 11569 17691
rect 11621 17639 11677 17691
rect 11729 17639 11749 17691
rect 11549 17583 11749 17639
rect 11549 17531 11569 17583
rect 11621 17531 11677 17583
rect 11729 17531 11749 17583
rect 11549 17475 11749 17531
rect 11549 17423 11569 17475
rect 11621 17423 11677 17475
rect 11729 17423 11749 17475
rect 11549 17367 11749 17423
rect 11549 17315 11569 17367
rect 11621 17315 11677 17367
rect 11729 17315 11749 17367
rect 11549 17259 11749 17315
rect 11549 17207 11569 17259
rect 11621 17207 11677 17259
rect 11729 17207 11749 17259
rect 11549 17151 11749 17207
rect 11549 17099 11569 17151
rect 11621 17099 11677 17151
rect 11729 17099 11749 17151
rect 11549 17043 11749 17099
rect 11549 16991 11569 17043
rect 11621 16991 11677 17043
rect 11729 16991 11749 17043
rect 11549 16935 11749 16991
rect 11549 16883 11569 16935
rect 11621 16883 11677 16935
rect 11729 16883 11749 16935
rect 11549 16827 11749 16883
rect 11549 16775 11569 16827
rect 11621 16775 11677 16827
rect 11729 16775 11749 16827
rect 11549 16719 11749 16775
rect 11549 16667 11569 16719
rect 11621 16667 11677 16719
rect 11729 16667 11749 16719
rect 11549 16611 11749 16667
rect 11549 16559 11569 16611
rect 11621 16559 11677 16611
rect 11729 16559 11749 16611
rect 11549 16503 11749 16559
rect 11549 16451 11569 16503
rect 11621 16451 11677 16503
rect 11729 16451 11749 16503
rect 11549 16395 11749 16451
rect 11549 16343 11569 16395
rect 11621 16343 11677 16395
rect 11729 16343 11749 16395
rect 11549 16287 11749 16343
rect 11549 16235 11569 16287
rect 11621 16235 11677 16287
rect 11729 16235 11749 16287
rect 11549 16179 11749 16235
rect 11549 16127 11569 16179
rect 11621 16127 11677 16179
rect 11729 16127 11749 16179
rect 11549 16071 11749 16127
rect 11549 16019 11569 16071
rect 11621 16019 11677 16071
rect 11729 16019 11749 16071
rect 11549 15963 11749 16019
rect 11549 15911 11569 15963
rect 11621 15911 11677 15963
rect 11729 15911 11749 15963
rect 11549 15855 11749 15911
rect 11549 15803 11569 15855
rect 11621 15803 11677 15855
rect 11729 15803 11749 15855
rect 11549 15747 11749 15803
rect 11549 15695 11569 15747
rect 11621 15695 11677 15747
rect 11729 15695 11749 15747
rect 11549 15639 11749 15695
rect 11549 15587 11569 15639
rect 11621 15587 11677 15639
rect 11729 15587 11749 15639
rect 11549 15531 11749 15587
rect 11549 15479 11569 15531
rect 11621 15479 11677 15531
rect 11729 15479 11749 15531
rect 11549 15423 11749 15479
rect 11549 15371 11569 15423
rect 11621 15371 11677 15423
rect 11729 15371 11749 15423
rect 11549 15315 11749 15371
rect 11549 15263 11569 15315
rect 11621 15263 11677 15315
rect 11729 15263 11749 15315
rect 11549 15207 11749 15263
rect 11549 15155 11569 15207
rect 11621 15155 11677 15207
rect 11729 15155 11749 15207
rect 11549 15099 11749 15155
rect 11549 15047 11569 15099
rect 11621 15047 11677 15099
rect 11729 15047 11749 15099
rect 11549 14991 11749 15047
rect 11549 14939 11569 14991
rect 11621 14939 11677 14991
rect 11729 14939 11749 14991
rect 11549 14883 11749 14939
rect 11549 14831 11569 14883
rect 11621 14831 11677 14883
rect 11729 14831 11749 14883
rect 11549 14775 11749 14831
rect 11549 14723 11569 14775
rect 11621 14723 11677 14775
rect 11729 14723 11749 14775
rect 11549 14667 11749 14723
rect 11549 14615 11569 14667
rect 11621 14615 11677 14667
rect 11729 14615 11749 14667
rect 11549 14559 11749 14615
rect 11549 14507 11569 14559
rect 11621 14507 11677 14559
rect 11729 14507 11749 14559
rect 11549 14451 11749 14507
rect 11549 14399 11569 14451
rect 11621 14399 11677 14451
rect 11729 14399 11749 14451
rect 11549 14343 11749 14399
rect 11549 14291 11569 14343
rect 11621 14291 11677 14343
rect 11729 14291 11749 14343
rect 11549 14235 11749 14291
rect 11549 14183 11569 14235
rect 11621 14183 11677 14235
rect 11729 14183 11749 14235
rect 11549 14127 11749 14183
rect 11549 14075 11569 14127
rect 11621 14075 11677 14127
rect 11729 14075 11749 14127
rect 11549 14019 11749 14075
rect 11549 13967 11569 14019
rect 11621 13967 11677 14019
rect 11729 13967 11749 14019
rect 11549 13911 11749 13967
rect 11549 13859 11569 13911
rect 11621 13859 11677 13911
rect 11729 13859 11749 13911
rect 11549 13803 11749 13859
rect 11549 13751 11569 13803
rect 11621 13751 11677 13803
rect 11729 13751 11749 13803
rect 11549 13695 11749 13751
rect 11549 13643 11569 13695
rect 11621 13643 11677 13695
rect 11729 13643 11749 13695
rect 11549 13587 11749 13643
rect 11549 13535 11569 13587
rect 11621 13535 11677 13587
rect 11729 13535 11749 13587
rect 11549 13479 11749 13535
rect 11549 13427 11569 13479
rect 11621 13427 11677 13479
rect 11729 13427 11749 13479
rect 11549 13371 11749 13427
rect 11549 13319 11569 13371
rect 11621 13319 11677 13371
rect 11729 13319 11749 13371
rect 11549 13263 11749 13319
rect 11549 13211 11569 13263
rect 11621 13211 11677 13263
rect 11729 13211 11749 13263
rect 11549 12143 11749 13211
rect 11549 12091 11569 12143
rect 11621 12091 11677 12143
rect 11729 12091 11749 12143
rect 11549 12035 11749 12091
rect 11549 11983 11569 12035
rect 11621 11983 11677 12035
rect 11729 11983 11749 12035
rect 11549 11927 11749 11983
rect 11549 11875 11569 11927
rect 11621 11875 11677 11927
rect 11729 11875 11749 11927
rect 11549 11819 11749 11875
rect 11549 11767 11569 11819
rect 11621 11767 11677 11819
rect 11729 11767 11749 11819
rect 11549 11711 11749 11767
rect 11549 11659 11569 11711
rect 11621 11659 11677 11711
rect 11729 11659 11749 11711
rect 11549 11603 11749 11659
rect 11549 11551 11569 11603
rect 11621 11551 11677 11603
rect 11729 11551 11749 11603
rect 11549 11495 11749 11551
rect 11549 11443 11569 11495
rect 11621 11443 11677 11495
rect 11729 11443 11749 11495
rect 11549 11387 11749 11443
rect 11549 11335 11569 11387
rect 11621 11335 11677 11387
rect 11729 11335 11749 11387
rect 11549 11279 11749 11335
rect 11549 11227 11569 11279
rect 11621 11227 11677 11279
rect 11729 11227 11749 11279
rect 11549 11171 11749 11227
rect 11549 11119 11569 11171
rect 11621 11119 11677 11171
rect 11729 11119 11749 11171
rect 11549 11063 11749 11119
rect 11549 11011 11569 11063
rect 11621 11011 11677 11063
rect 11729 11011 11749 11063
rect 11549 10955 11749 11011
rect 11549 10903 11569 10955
rect 11621 10903 11677 10955
rect 11729 10903 11749 10955
rect 11549 10847 11749 10903
rect 11549 10795 11569 10847
rect 11621 10795 11677 10847
rect 11729 10795 11749 10847
rect 11549 10739 11749 10795
rect 11549 10687 11569 10739
rect 11621 10687 11677 10739
rect 11729 10687 11749 10739
rect 11549 10631 11749 10687
rect 11549 10579 11569 10631
rect 11621 10579 11677 10631
rect 11729 10579 11749 10631
rect 11549 10523 11749 10579
rect 11549 10471 11569 10523
rect 11621 10471 11677 10523
rect 11729 10471 11749 10523
rect 11549 10415 11749 10471
rect 11549 10363 11569 10415
rect 11621 10363 11677 10415
rect 11729 10363 11749 10415
rect 11549 10307 11749 10363
rect 11549 10255 11569 10307
rect 11621 10255 11677 10307
rect 11729 10255 11749 10307
rect 11549 10199 11749 10255
rect 11549 10147 11569 10199
rect 11621 10147 11677 10199
rect 11729 10147 11749 10199
rect 11549 10091 11749 10147
rect 11549 10039 11569 10091
rect 11621 10039 11677 10091
rect 11729 10039 11749 10091
rect 11549 9983 11749 10039
rect 11549 9931 11569 9983
rect 11621 9931 11677 9983
rect 11729 9931 11749 9983
rect 11549 9875 11749 9931
rect 11549 9823 11569 9875
rect 11621 9823 11677 9875
rect 11729 9823 11749 9875
rect 11549 9767 11749 9823
rect 11549 9715 11569 9767
rect 11621 9715 11677 9767
rect 11729 9715 11749 9767
rect 11549 9659 11749 9715
rect 11549 9607 11569 9659
rect 11621 9607 11677 9659
rect 11729 9607 11749 9659
rect 11549 9551 11749 9607
rect 11549 9499 11569 9551
rect 11621 9499 11677 9551
rect 11729 9499 11749 9551
rect 11549 9443 11749 9499
rect 11549 9391 11569 9443
rect 11621 9391 11677 9443
rect 11729 9391 11749 9443
rect 11549 9335 11749 9391
rect 11549 9283 11569 9335
rect 11621 9283 11677 9335
rect 11729 9283 11749 9335
rect 11549 9227 11749 9283
rect 11549 9175 11569 9227
rect 11621 9175 11677 9227
rect 11729 9175 11749 9227
rect 11549 9119 11749 9175
rect 11549 9067 11569 9119
rect 11621 9067 11677 9119
rect 11729 9067 11749 9119
rect 11549 9011 11749 9067
rect 11549 8959 11569 9011
rect 11621 8959 11677 9011
rect 11729 8959 11749 9011
rect 11549 8903 11749 8959
rect 11549 8851 11569 8903
rect 11621 8851 11677 8903
rect 11729 8851 11749 8903
rect 11549 8795 11749 8851
rect 11549 8743 11569 8795
rect 11621 8743 11677 8795
rect 11729 8743 11749 8795
rect 11549 8687 11749 8743
rect 11549 8635 11569 8687
rect 11621 8635 11677 8687
rect 11729 8635 11749 8687
rect 11549 8579 11749 8635
rect 11549 8527 11569 8579
rect 11621 8527 11677 8579
rect 11729 8527 11749 8579
rect 11549 8471 11749 8527
rect 11549 8419 11569 8471
rect 11621 8419 11677 8471
rect 11729 8419 11749 8471
rect 11549 8363 11749 8419
rect 11549 8311 11569 8363
rect 11621 8311 11677 8363
rect 11729 8311 11749 8363
rect 11549 8255 11749 8311
rect 11549 8203 11569 8255
rect 11621 8203 11677 8255
rect 11729 8203 11749 8255
rect 11549 8147 11749 8203
rect 11549 8095 11569 8147
rect 11621 8095 11677 8147
rect 11729 8095 11749 8147
rect 11549 8039 11749 8095
rect 11549 7987 11569 8039
rect 11621 7987 11677 8039
rect 11729 7987 11749 8039
rect 11549 7931 11749 7987
rect 11549 7879 11569 7931
rect 11621 7879 11677 7931
rect 11729 7879 11749 7931
rect 11549 7823 11749 7879
rect 11549 7771 11569 7823
rect 11621 7771 11677 7823
rect 11729 7771 11749 7823
rect 11549 7715 11749 7771
rect 11549 7663 11569 7715
rect 11621 7663 11677 7715
rect 11729 7663 11749 7715
rect 11549 7607 11749 7663
rect 11549 7555 11569 7607
rect 11621 7555 11677 7607
rect 11729 7555 11749 7607
rect 11549 7499 11749 7555
rect 11549 7447 11569 7499
rect 11621 7447 11677 7499
rect 11729 7447 11749 7499
rect 11549 7391 11749 7447
rect 11549 7339 11569 7391
rect 11621 7339 11677 7391
rect 11729 7339 11749 7391
rect 11549 6271 11749 7339
rect 11549 6219 11569 6271
rect 11621 6219 11677 6271
rect 11729 6219 11749 6271
rect 11549 6163 11749 6219
rect 11549 6111 11569 6163
rect 11621 6111 11677 6163
rect 11729 6111 11749 6163
rect 11549 6055 11749 6111
rect 11549 6003 11569 6055
rect 11621 6003 11677 6055
rect 11729 6003 11749 6055
rect 11549 5947 11749 6003
rect 11549 5895 11569 5947
rect 11621 5895 11677 5947
rect 11729 5895 11749 5947
rect 11549 5839 11749 5895
rect 11549 5787 11569 5839
rect 11621 5787 11677 5839
rect 11729 5787 11749 5839
rect 11549 5731 11749 5787
rect 11549 5679 11569 5731
rect 11621 5679 11677 5731
rect 11729 5679 11749 5731
rect 11549 5623 11749 5679
rect 11549 5571 11569 5623
rect 11621 5571 11677 5623
rect 11729 5571 11749 5623
rect 11549 5515 11749 5571
rect 11549 5463 11569 5515
rect 11621 5463 11677 5515
rect 11729 5463 11749 5515
rect 11549 5407 11749 5463
rect 11549 5355 11569 5407
rect 11621 5355 11677 5407
rect 11729 5355 11749 5407
rect 11549 5299 11749 5355
rect 11549 5247 11569 5299
rect 11621 5247 11677 5299
rect 11729 5247 11749 5299
rect 11549 5191 11749 5247
rect 11549 5139 11569 5191
rect 11621 5139 11677 5191
rect 11729 5139 11749 5191
rect 11549 5083 11749 5139
rect 11549 5031 11569 5083
rect 11621 5031 11677 5083
rect 11729 5031 11749 5083
rect 11549 4975 11749 5031
rect 11549 4923 11569 4975
rect 11621 4923 11677 4975
rect 11729 4923 11749 4975
rect 11549 4867 11749 4923
rect 11549 4815 11569 4867
rect 11621 4815 11677 4867
rect 11729 4815 11749 4867
rect 11549 4759 11749 4815
rect 11549 4707 11569 4759
rect 11621 4707 11677 4759
rect 11729 4707 11749 4759
rect 11549 4651 11749 4707
rect 11549 4599 11569 4651
rect 11621 4599 11677 4651
rect 11729 4599 11749 4651
rect 11549 4543 11749 4599
rect 11549 4491 11569 4543
rect 11621 4491 11677 4543
rect 11729 4491 11749 4543
rect 11549 4435 11749 4491
rect 11549 4383 11569 4435
rect 11621 4383 11677 4435
rect 11729 4383 11749 4435
rect 11549 4327 11749 4383
rect 11549 4275 11569 4327
rect 11621 4275 11677 4327
rect 11729 4275 11749 4327
rect 11549 4219 11749 4275
rect 11549 4167 11569 4219
rect 11621 4167 11677 4219
rect 11729 4167 11749 4219
rect 11549 4111 11749 4167
rect 11549 4059 11569 4111
rect 11621 4059 11677 4111
rect 11729 4059 11749 4111
rect 11549 4003 11749 4059
rect 11549 3951 11569 4003
rect 11621 3951 11677 4003
rect 11729 3951 11749 4003
rect 11549 3895 11749 3951
rect 11549 3843 11569 3895
rect 11621 3843 11677 3895
rect 11729 3843 11749 3895
rect 11549 3787 11749 3843
rect 11549 3735 11569 3787
rect 11621 3735 11677 3787
rect 11729 3735 11749 3787
rect 11549 3679 11749 3735
rect 11549 3627 11569 3679
rect 11621 3627 11677 3679
rect 11729 3627 11749 3679
rect 11549 3571 11749 3627
rect 11549 3519 11569 3571
rect 11621 3519 11677 3571
rect 11729 3519 11749 3571
rect 11549 3463 11749 3519
rect 11549 3411 11569 3463
rect 11621 3411 11677 3463
rect 11729 3411 11749 3463
rect 11549 3355 11749 3411
rect 11549 3303 11569 3355
rect 11621 3303 11677 3355
rect 11729 3303 11749 3355
rect 11549 3247 11749 3303
rect 11549 3195 11569 3247
rect 11621 3195 11677 3247
rect 11729 3195 11749 3247
rect 11549 3139 11749 3195
rect 11549 3087 11569 3139
rect 11621 3087 11677 3139
rect 11729 3087 11749 3139
rect 11549 3031 11749 3087
rect 11549 2979 11569 3031
rect 11621 2979 11677 3031
rect 11729 2979 11749 3031
rect 11549 2923 11749 2979
rect 11549 2871 11569 2923
rect 11621 2871 11677 2923
rect 11729 2871 11749 2923
rect 11549 2815 11749 2871
rect 11549 2763 11569 2815
rect 11621 2763 11677 2815
rect 11729 2763 11749 2815
rect 11549 2707 11749 2763
rect 11549 2655 11569 2707
rect 11621 2655 11677 2707
rect 11729 2655 11749 2707
rect 11549 2599 11749 2655
rect 11549 2547 11569 2599
rect 11621 2547 11677 2599
rect 11729 2547 11749 2599
rect 11549 2491 11749 2547
rect 11549 2439 11569 2491
rect 11621 2439 11677 2491
rect 11729 2439 11749 2491
rect 11549 2383 11749 2439
rect 11549 2331 11569 2383
rect 11621 2331 11677 2383
rect 11729 2331 11749 2383
rect 11549 2275 11749 2331
rect 11549 2223 11569 2275
rect 11621 2223 11677 2275
rect 11729 2223 11749 2275
rect 11549 2167 11749 2223
rect 11549 2115 11569 2167
rect 11621 2115 11677 2167
rect 11729 2115 11749 2167
rect 11549 2059 11749 2115
rect 11549 2007 11569 2059
rect 11621 2007 11677 2059
rect 11729 2007 11749 2059
rect 11549 1951 11749 2007
rect 11549 1899 11569 1951
rect 11621 1899 11677 1951
rect 11729 1899 11749 1951
rect 11549 1843 11749 1899
rect 11549 1791 11569 1843
rect 11621 1791 11677 1843
rect 11729 1791 11749 1843
rect 11549 1735 11749 1791
rect 11549 1683 11569 1735
rect 11621 1683 11677 1735
rect 11729 1683 11749 1735
rect 11549 1627 11749 1683
rect 11549 1575 11569 1627
rect 11621 1575 11677 1627
rect 11729 1575 11749 1627
rect 11549 1519 11749 1575
rect 11549 1467 11569 1519
rect 11621 1467 11677 1519
rect 11729 1467 11749 1519
rect 11549 1455 11749 1467
rect 11809 24691 13709 25617
rect 11809 24639 12051 24691
rect 12103 24639 12159 24691
rect 12211 24639 12267 24691
rect 12319 24639 13709 24691
rect 11809 24583 13709 24639
rect 11809 24531 12051 24583
rect 12103 24531 12159 24583
rect 12211 24531 12267 24583
rect 12319 24531 13709 24583
rect 11809 24475 13709 24531
rect 11809 24423 12051 24475
rect 12103 24423 12159 24475
rect 12211 24423 12267 24475
rect 12319 24423 13709 24475
rect 11809 24367 13709 24423
rect 11809 24315 12051 24367
rect 12103 24315 12159 24367
rect 12211 24315 12267 24367
rect 12319 24315 13709 24367
rect 11809 24259 13709 24315
rect 11809 24207 12051 24259
rect 12103 24207 12159 24259
rect 12211 24207 12267 24259
rect 12319 24207 13709 24259
rect 11809 24151 13709 24207
rect 11809 24099 12051 24151
rect 12103 24099 12159 24151
rect 12211 24099 12267 24151
rect 12319 24099 13709 24151
rect 11809 24043 13709 24099
rect 11809 23991 12051 24043
rect 12103 23991 12159 24043
rect 12211 23991 12267 24043
rect 12319 23991 13709 24043
rect 11809 23935 13709 23991
rect 11809 23883 12051 23935
rect 12103 23883 12159 23935
rect 12211 23883 12267 23935
rect 12319 23883 13709 23935
rect 11809 23827 13709 23883
rect 11809 23775 12051 23827
rect 12103 23775 12159 23827
rect 12211 23775 12267 23827
rect 12319 23775 13709 23827
rect 11809 23719 13709 23775
rect 11809 23667 12051 23719
rect 12103 23667 12159 23719
rect 12211 23667 12267 23719
rect 12319 23667 13709 23719
rect 11809 23611 13709 23667
rect 11809 23559 12051 23611
rect 12103 23559 12159 23611
rect 12211 23559 12267 23611
rect 12319 23559 13709 23611
rect 11809 23503 13709 23559
rect 11809 23451 12051 23503
rect 12103 23451 12159 23503
rect 12211 23451 12267 23503
rect 12319 23451 13709 23503
rect 11809 23395 13709 23451
rect 11809 23343 12051 23395
rect 12103 23343 12159 23395
rect 12211 23343 12267 23395
rect 12319 23343 13709 23395
rect 11809 23287 13709 23343
rect 11809 23235 12051 23287
rect 12103 23235 12159 23287
rect 12211 23235 12267 23287
rect 12319 23235 13709 23287
rect 11809 23179 13709 23235
rect 11809 23127 12051 23179
rect 12103 23127 12159 23179
rect 12211 23127 12267 23179
rect 12319 23127 13709 23179
rect 11809 23071 13709 23127
rect 11809 23019 12051 23071
rect 12103 23019 12159 23071
rect 12211 23019 12267 23071
rect 12319 23019 13709 23071
rect 11809 22963 13709 23019
rect 11809 22911 12051 22963
rect 12103 22911 12159 22963
rect 12211 22911 12267 22963
rect 12319 22911 13709 22963
rect 11809 22855 13709 22911
rect 11809 22803 12051 22855
rect 12103 22803 12159 22855
rect 12211 22803 12267 22855
rect 12319 22803 13709 22855
rect 11809 22747 13709 22803
rect 11809 22695 12051 22747
rect 12103 22695 12159 22747
rect 12211 22695 12267 22747
rect 12319 22695 13709 22747
rect 11809 22639 13709 22695
rect 11809 22587 12051 22639
rect 12103 22587 12159 22639
rect 12211 22587 12267 22639
rect 12319 22587 13709 22639
rect 11809 22531 13709 22587
rect 11809 22479 12051 22531
rect 12103 22479 12159 22531
rect 12211 22479 12267 22531
rect 12319 22479 13709 22531
rect 11809 22423 13709 22479
rect 11809 22371 12051 22423
rect 12103 22371 12159 22423
rect 12211 22371 12267 22423
rect 12319 22371 13709 22423
rect 11809 22315 13709 22371
rect 11809 22263 12051 22315
rect 12103 22263 12159 22315
rect 12211 22263 12267 22315
rect 12319 22263 13709 22315
rect 11809 22207 13709 22263
rect 11809 22155 12051 22207
rect 12103 22155 12159 22207
rect 12211 22155 12267 22207
rect 12319 22155 13709 22207
rect 11809 22099 13709 22155
rect 11809 22047 12051 22099
rect 12103 22047 12159 22099
rect 12211 22047 12267 22099
rect 12319 22047 13709 22099
rect 11809 21991 13709 22047
rect 11809 21939 12051 21991
rect 12103 21939 12159 21991
rect 12211 21939 12267 21991
rect 12319 21939 13709 21991
rect 11809 21883 13709 21939
rect 11809 21831 12051 21883
rect 12103 21831 12159 21883
rect 12211 21831 12267 21883
rect 12319 21831 13709 21883
rect 11809 21775 13709 21831
rect 11809 21723 12051 21775
rect 12103 21723 12159 21775
rect 12211 21723 12267 21775
rect 12319 21723 13709 21775
rect 11809 21667 13709 21723
rect 11809 21615 12051 21667
rect 12103 21615 12159 21667
rect 12211 21615 12267 21667
rect 12319 21615 13709 21667
rect 11809 21559 13709 21615
rect 11809 21507 12051 21559
rect 12103 21507 12159 21559
rect 12211 21507 12267 21559
rect 12319 21507 13709 21559
rect 11809 21451 13709 21507
rect 11809 21399 12051 21451
rect 12103 21399 12159 21451
rect 12211 21399 12267 21451
rect 12319 21399 13709 21451
rect 11809 21343 13709 21399
rect 11809 21291 12051 21343
rect 12103 21291 12159 21343
rect 12211 21291 12267 21343
rect 12319 21291 13709 21343
rect 11809 21235 13709 21291
rect 11809 21183 12051 21235
rect 12103 21183 12159 21235
rect 12211 21183 12267 21235
rect 12319 21183 13709 21235
rect 11809 21127 13709 21183
rect 11809 21075 12051 21127
rect 12103 21075 12159 21127
rect 12211 21075 12267 21127
rect 12319 21075 13709 21127
rect 11809 21019 13709 21075
rect 11809 20967 12051 21019
rect 12103 20967 12159 21019
rect 12211 20967 12267 21019
rect 12319 20967 13709 21019
rect 11809 20911 13709 20967
rect 11809 20859 12051 20911
rect 12103 20859 12159 20911
rect 12211 20859 12267 20911
rect 12319 20859 13709 20911
rect 11809 20803 13709 20859
rect 11809 20751 12051 20803
rect 12103 20751 12159 20803
rect 12211 20751 12267 20803
rect 12319 20751 13709 20803
rect 11809 20695 13709 20751
rect 11809 20643 12051 20695
rect 12103 20643 12159 20695
rect 12211 20643 12267 20695
rect 12319 20643 13709 20695
rect 11809 20587 13709 20643
rect 11809 20535 12051 20587
rect 12103 20535 12159 20587
rect 12211 20535 12267 20587
rect 12319 20535 13709 20587
rect 11809 20479 13709 20535
rect 11809 20427 12051 20479
rect 12103 20427 12159 20479
rect 12211 20427 12267 20479
rect 12319 20427 13709 20479
rect 11809 20371 13709 20427
rect 11809 20319 12051 20371
rect 12103 20319 12159 20371
rect 12211 20319 12267 20371
rect 12319 20319 13709 20371
rect 11809 20263 13709 20319
rect 11809 20211 12051 20263
rect 12103 20211 12159 20263
rect 12211 20211 12267 20263
rect 12319 20211 13709 20263
rect 11809 20155 13709 20211
rect 11809 20103 12051 20155
rect 12103 20103 12159 20155
rect 12211 20103 12267 20155
rect 12319 20103 13709 20155
rect 11809 20047 13709 20103
rect 11809 19995 12051 20047
rect 12103 19995 12159 20047
rect 12211 19995 12267 20047
rect 12319 19995 13709 20047
rect 11809 19939 13709 19995
rect 11809 19887 12051 19939
rect 12103 19887 12159 19939
rect 12211 19887 12267 19939
rect 12319 19887 13709 19939
rect 11809 19831 13709 19887
rect 11809 19779 12051 19831
rect 12103 19779 12159 19831
rect 12211 19779 12267 19831
rect 12319 19779 13709 19831
rect 11809 19723 13709 19779
rect 11809 19671 12051 19723
rect 12103 19671 12159 19723
rect 12211 19671 12267 19723
rect 12319 19671 13709 19723
rect 11809 19615 13709 19671
rect 11809 19563 12051 19615
rect 12103 19563 12159 19615
rect 12211 19563 12267 19615
rect 12319 19563 13709 19615
rect 11809 19507 13709 19563
rect 11809 19455 12051 19507
rect 12103 19455 12159 19507
rect 12211 19455 12267 19507
rect 12319 19455 13709 19507
rect 11809 19399 13709 19455
rect 11809 19347 12051 19399
rect 12103 19347 12159 19399
rect 12211 19347 12267 19399
rect 12319 19347 13709 19399
rect 11809 19291 13709 19347
rect 11809 19239 12051 19291
rect 12103 19239 12159 19291
rect 12211 19239 12267 19291
rect 12319 19239 13709 19291
rect 11809 19183 13709 19239
rect 11809 19131 12051 19183
rect 12103 19131 12159 19183
rect 12211 19131 12267 19183
rect 12319 19131 13709 19183
rect 11809 19075 13709 19131
rect 11809 19023 12051 19075
rect 12103 19023 12159 19075
rect 12211 19023 12267 19075
rect 12319 19023 13709 19075
rect 11809 18967 13709 19023
rect 11809 18915 12051 18967
rect 12103 18915 12159 18967
rect 12211 18915 12267 18967
rect 12319 18915 13709 18967
rect 11809 18859 13709 18915
rect 11809 18807 12051 18859
rect 12103 18807 12159 18859
rect 12211 18807 12267 18859
rect 12319 18807 13709 18859
rect 11809 18751 13709 18807
rect 11809 18699 12051 18751
rect 12103 18699 12159 18751
rect 12211 18699 12267 18751
rect 12319 18699 13709 18751
rect 11809 18643 13709 18699
rect 11809 18591 12051 18643
rect 12103 18591 12159 18643
rect 12211 18591 12267 18643
rect 12319 18591 13709 18643
rect 11809 18535 13709 18591
rect 11809 18483 12051 18535
rect 12103 18483 12159 18535
rect 12211 18483 12267 18535
rect 12319 18483 13709 18535
rect 11809 18427 13709 18483
rect 11809 18375 12051 18427
rect 12103 18375 12159 18427
rect 12211 18375 12267 18427
rect 12319 18375 13709 18427
rect 11809 18319 13709 18375
rect 11809 18267 12051 18319
rect 12103 18267 12159 18319
rect 12211 18267 12267 18319
rect 12319 18267 13709 18319
rect 11809 18211 13709 18267
rect 11809 18159 12051 18211
rect 12103 18159 12159 18211
rect 12211 18159 12267 18211
rect 12319 18159 13709 18211
rect 11809 18103 13709 18159
rect 11809 18051 12051 18103
rect 12103 18051 12159 18103
rect 12211 18051 12267 18103
rect 12319 18051 13709 18103
rect 11809 17995 13709 18051
rect 11809 17943 12051 17995
rect 12103 17943 12159 17995
rect 12211 17943 12267 17995
rect 12319 17943 13709 17995
rect 11809 17887 13709 17943
rect 11809 17835 12051 17887
rect 12103 17835 12159 17887
rect 12211 17835 12267 17887
rect 12319 17835 13709 17887
rect 11809 17779 13709 17835
rect 11809 17727 12051 17779
rect 12103 17727 12159 17779
rect 12211 17727 12267 17779
rect 12319 17727 13709 17779
rect 11809 17671 13709 17727
rect 11809 17619 12051 17671
rect 12103 17619 12159 17671
rect 12211 17619 12267 17671
rect 12319 17619 13709 17671
rect 11809 17563 13709 17619
rect 11809 17511 12051 17563
rect 12103 17511 12159 17563
rect 12211 17511 12267 17563
rect 12319 17511 13709 17563
rect 11809 17455 13709 17511
rect 11809 17403 12051 17455
rect 12103 17403 12159 17455
rect 12211 17403 12267 17455
rect 12319 17403 13709 17455
rect 11809 17347 13709 17403
rect 11809 17295 12051 17347
rect 12103 17295 12159 17347
rect 12211 17295 12267 17347
rect 12319 17295 13709 17347
rect 11809 17239 13709 17295
rect 11809 17187 12051 17239
rect 12103 17187 12159 17239
rect 12211 17187 12267 17239
rect 12319 17187 13709 17239
rect 11809 17131 13709 17187
rect 11809 17079 12051 17131
rect 12103 17079 12159 17131
rect 12211 17079 12267 17131
rect 12319 17079 13709 17131
rect 11809 17023 13709 17079
rect 11809 16971 12051 17023
rect 12103 16971 12159 17023
rect 12211 16971 12267 17023
rect 12319 16971 13709 17023
rect 11809 16915 13709 16971
rect 11809 16863 12051 16915
rect 12103 16863 12159 16915
rect 12211 16863 12267 16915
rect 12319 16863 13709 16915
rect 11809 16807 13709 16863
rect 11809 16755 12051 16807
rect 12103 16755 12159 16807
rect 12211 16755 12267 16807
rect 12319 16755 13709 16807
rect 11809 16699 13709 16755
rect 11809 16647 12051 16699
rect 12103 16647 12159 16699
rect 12211 16647 12267 16699
rect 12319 16647 13709 16699
rect 11809 16591 13709 16647
rect 11809 16539 12051 16591
rect 12103 16539 12159 16591
rect 12211 16539 12267 16591
rect 12319 16539 13709 16591
rect 11809 16483 13709 16539
rect 11809 16431 12051 16483
rect 12103 16431 12159 16483
rect 12211 16431 12267 16483
rect 12319 16431 13709 16483
rect 11809 16375 13709 16431
rect 11809 16323 12051 16375
rect 12103 16323 12159 16375
rect 12211 16323 12267 16375
rect 12319 16323 13709 16375
rect 11809 16267 13709 16323
rect 11809 16215 12051 16267
rect 12103 16215 12159 16267
rect 12211 16215 12267 16267
rect 12319 16215 13709 16267
rect 11809 16159 13709 16215
rect 11809 16107 12051 16159
rect 12103 16107 12159 16159
rect 12211 16107 12267 16159
rect 12319 16107 13709 16159
rect 11809 16051 13709 16107
rect 11809 15999 12051 16051
rect 12103 15999 12159 16051
rect 12211 15999 12267 16051
rect 12319 15999 13709 16051
rect 11809 15943 13709 15999
rect 11809 15891 12051 15943
rect 12103 15891 12159 15943
rect 12211 15891 12267 15943
rect 12319 15891 13709 15943
rect 11809 15835 13709 15891
rect 11809 15783 12051 15835
rect 12103 15783 12159 15835
rect 12211 15783 12267 15835
rect 12319 15783 13709 15835
rect 11809 15727 13709 15783
rect 11809 15675 12051 15727
rect 12103 15675 12159 15727
rect 12211 15675 12267 15727
rect 12319 15675 13709 15727
rect 11809 15619 13709 15675
rect 11809 15567 12051 15619
rect 12103 15567 12159 15619
rect 12211 15567 12267 15619
rect 12319 15567 13709 15619
rect 11809 15511 13709 15567
rect 11809 15459 12051 15511
rect 12103 15459 12159 15511
rect 12211 15459 12267 15511
rect 12319 15459 13709 15511
rect 11809 15403 13709 15459
rect 11809 15351 12051 15403
rect 12103 15351 12159 15403
rect 12211 15351 12267 15403
rect 12319 15351 13709 15403
rect 11809 15295 13709 15351
rect 11809 15243 12051 15295
rect 12103 15243 12159 15295
rect 12211 15243 12267 15295
rect 12319 15243 13709 15295
rect 11809 15187 13709 15243
rect 11809 15135 12051 15187
rect 12103 15135 12159 15187
rect 12211 15135 12267 15187
rect 12319 15135 13709 15187
rect 11809 15079 13709 15135
rect 11809 15027 12051 15079
rect 12103 15027 12159 15079
rect 12211 15027 12267 15079
rect 12319 15027 13709 15079
rect 11809 14971 13709 15027
rect 11809 14919 12051 14971
rect 12103 14919 12159 14971
rect 12211 14919 12267 14971
rect 12319 14919 13709 14971
rect 11809 14863 13709 14919
rect 11809 14811 12051 14863
rect 12103 14811 12159 14863
rect 12211 14811 12267 14863
rect 12319 14811 13709 14863
rect 11809 14755 13709 14811
rect 11809 14703 12051 14755
rect 12103 14703 12159 14755
rect 12211 14703 12267 14755
rect 12319 14703 13709 14755
rect 11809 14647 13709 14703
rect 11809 14595 12051 14647
rect 12103 14595 12159 14647
rect 12211 14595 12267 14647
rect 12319 14595 13709 14647
rect 11809 14539 13709 14595
rect 11809 14487 12051 14539
rect 12103 14487 12159 14539
rect 12211 14487 12267 14539
rect 12319 14487 13709 14539
rect 11809 14431 13709 14487
rect 11809 14379 12051 14431
rect 12103 14379 12159 14431
rect 12211 14379 12267 14431
rect 12319 14379 13709 14431
rect 11809 14323 13709 14379
rect 11809 14271 12051 14323
rect 12103 14271 12159 14323
rect 12211 14271 12267 14323
rect 12319 14271 13709 14323
rect 11809 14215 13709 14271
rect 11809 14163 12051 14215
rect 12103 14163 12159 14215
rect 12211 14163 12267 14215
rect 12319 14163 13709 14215
rect 11809 14107 13709 14163
rect 11809 14055 12051 14107
rect 12103 14055 12159 14107
rect 12211 14055 12267 14107
rect 12319 14055 13709 14107
rect 11809 13999 13709 14055
rect 11809 13947 12051 13999
rect 12103 13947 12159 13999
rect 12211 13947 12267 13999
rect 12319 13947 13709 13999
rect 11809 13891 13709 13947
rect 11809 13839 12051 13891
rect 12103 13839 12159 13891
rect 12211 13839 12267 13891
rect 12319 13839 13709 13891
rect 11809 13783 13709 13839
rect 11809 13731 12051 13783
rect 12103 13731 12159 13783
rect 12211 13731 12267 13783
rect 12319 13731 13709 13783
rect 11809 13675 13709 13731
rect 11809 13623 12051 13675
rect 12103 13623 12159 13675
rect 12211 13623 12267 13675
rect 12319 13623 13709 13675
rect 11809 13567 13709 13623
rect 11809 13515 12051 13567
rect 12103 13515 12159 13567
rect 12211 13515 12267 13567
rect 12319 13515 13709 13567
rect 11809 13459 13709 13515
rect 11809 13407 12051 13459
rect 12103 13407 12159 13459
rect 12211 13407 12267 13459
rect 12319 13407 13709 13459
rect 11809 13351 13709 13407
rect 11809 13299 12051 13351
rect 12103 13299 12159 13351
rect 12211 13299 12267 13351
rect 12319 13299 13709 13351
rect 11809 13243 13709 13299
rect 11809 13191 12051 13243
rect 12103 13191 12159 13243
rect 12211 13191 12267 13243
rect 12319 13191 13709 13243
rect 11809 13135 13709 13191
rect 11809 13083 12051 13135
rect 12103 13083 12159 13135
rect 12211 13083 12267 13135
rect 12319 13083 13709 13135
rect 11809 13027 13709 13083
rect 11809 12975 12051 13027
rect 12103 12975 12159 13027
rect 12211 12975 12267 13027
rect 12319 12975 13709 13027
rect 11809 12919 13709 12975
rect 11809 12867 12051 12919
rect 12103 12867 12159 12919
rect 12211 12867 12267 12919
rect 12319 12867 13709 12919
rect 11809 12811 13709 12867
rect 11809 12759 12051 12811
rect 12103 12759 12159 12811
rect 12211 12759 12267 12811
rect 12319 12759 13709 12811
rect 11809 12703 13709 12759
rect 11809 12651 12051 12703
rect 12103 12651 12159 12703
rect 12211 12651 12267 12703
rect 12319 12651 13709 12703
rect 11809 12595 13709 12651
rect 11809 12543 12051 12595
rect 12103 12543 12159 12595
rect 12211 12543 12267 12595
rect 12319 12543 13709 12595
rect 11809 12487 13709 12543
rect 11809 12435 12051 12487
rect 12103 12435 12159 12487
rect 12211 12435 12267 12487
rect 12319 12435 13709 12487
rect 11809 12379 13709 12435
rect 11809 12327 12051 12379
rect 12103 12327 12159 12379
rect 12211 12327 12267 12379
rect 12319 12327 13709 12379
rect 11809 12271 13709 12327
rect 11809 12219 12051 12271
rect 12103 12219 12159 12271
rect 12211 12219 12267 12271
rect 12319 12219 13709 12271
rect 11809 12163 13709 12219
rect 11809 12111 12051 12163
rect 12103 12111 12159 12163
rect 12211 12111 12267 12163
rect 12319 12111 13709 12163
rect 11809 12055 13709 12111
rect 11809 12003 12051 12055
rect 12103 12003 12159 12055
rect 12211 12003 12267 12055
rect 12319 12003 13709 12055
rect 11809 11947 13709 12003
rect 11809 11895 12051 11947
rect 12103 11895 12159 11947
rect 12211 11895 12267 11947
rect 12319 11895 13709 11947
rect 11809 11839 13709 11895
rect 11809 11787 12051 11839
rect 12103 11787 12159 11839
rect 12211 11787 12267 11839
rect 12319 11787 13709 11839
rect 11809 11731 13709 11787
rect 11809 11679 12051 11731
rect 12103 11679 12159 11731
rect 12211 11679 12267 11731
rect 12319 11679 13709 11731
rect 11809 11623 13709 11679
rect 11809 11571 12051 11623
rect 12103 11571 12159 11623
rect 12211 11571 12267 11623
rect 12319 11571 13709 11623
rect 11809 11515 13709 11571
rect 11809 11463 12051 11515
rect 12103 11463 12159 11515
rect 12211 11463 12267 11515
rect 12319 11463 13709 11515
rect 11809 11407 13709 11463
rect 11809 11355 12051 11407
rect 12103 11355 12159 11407
rect 12211 11355 12267 11407
rect 12319 11355 13709 11407
rect 11809 11299 13709 11355
rect 11809 11247 12051 11299
rect 12103 11247 12159 11299
rect 12211 11247 12267 11299
rect 12319 11247 13709 11299
rect 11809 11191 13709 11247
rect 11809 11139 12051 11191
rect 12103 11139 12159 11191
rect 12211 11139 12267 11191
rect 12319 11139 13709 11191
rect 11809 11083 13709 11139
rect 11809 11031 12051 11083
rect 12103 11031 12159 11083
rect 12211 11031 12267 11083
rect 12319 11031 13709 11083
rect 11809 10975 13709 11031
rect 11809 10923 12051 10975
rect 12103 10923 12159 10975
rect 12211 10923 12267 10975
rect 12319 10923 13709 10975
rect 11809 10867 13709 10923
rect 11809 10815 12051 10867
rect 12103 10815 12159 10867
rect 12211 10815 12267 10867
rect 12319 10815 13709 10867
rect 11809 10759 13709 10815
rect 11809 10707 12051 10759
rect 12103 10707 12159 10759
rect 12211 10707 12267 10759
rect 12319 10707 13709 10759
rect 11809 10651 13709 10707
rect 11809 10599 12051 10651
rect 12103 10599 12159 10651
rect 12211 10599 12267 10651
rect 12319 10599 13709 10651
rect 11809 10543 13709 10599
rect 11809 10491 12051 10543
rect 12103 10491 12159 10543
rect 12211 10491 12267 10543
rect 12319 10491 13709 10543
rect 11809 10435 13709 10491
rect 11809 10383 12051 10435
rect 12103 10383 12159 10435
rect 12211 10383 12267 10435
rect 12319 10383 13709 10435
rect 11809 10327 13709 10383
rect 11809 10275 12051 10327
rect 12103 10275 12159 10327
rect 12211 10275 12267 10327
rect 12319 10275 13709 10327
rect 11809 10219 13709 10275
rect 11809 10167 12051 10219
rect 12103 10167 12159 10219
rect 12211 10167 12267 10219
rect 12319 10167 13709 10219
rect 11809 10111 13709 10167
rect 11809 10059 12051 10111
rect 12103 10059 12159 10111
rect 12211 10059 12267 10111
rect 12319 10059 13709 10111
rect 11809 10003 13709 10059
rect 11809 9951 12051 10003
rect 12103 9951 12159 10003
rect 12211 9951 12267 10003
rect 12319 9951 13709 10003
rect 11809 9895 13709 9951
rect 11809 9843 12051 9895
rect 12103 9843 12159 9895
rect 12211 9843 12267 9895
rect 12319 9843 13709 9895
rect 11809 9787 13709 9843
rect 11809 9735 12051 9787
rect 12103 9735 12159 9787
rect 12211 9735 12267 9787
rect 12319 9735 13709 9787
rect 11809 9679 13709 9735
rect 11809 9627 12051 9679
rect 12103 9627 12159 9679
rect 12211 9627 12267 9679
rect 12319 9627 13709 9679
rect 11809 9571 13709 9627
rect 11809 9519 12051 9571
rect 12103 9519 12159 9571
rect 12211 9519 12267 9571
rect 12319 9519 13709 9571
rect 11809 9463 13709 9519
rect 11809 9411 12051 9463
rect 12103 9411 12159 9463
rect 12211 9411 12267 9463
rect 12319 9411 13709 9463
rect 11809 9355 13709 9411
rect 11809 9303 12051 9355
rect 12103 9303 12159 9355
rect 12211 9303 12267 9355
rect 12319 9303 13709 9355
rect 11809 9247 13709 9303
rect 11809 9195 12051 9247
rect 12103 9195 12159 9247
rect 12211 9195 12267 9247
rect 12319 9195 13709 9247
rect 11809 9139 13709 9195
rect 11809 9087 12051 9139
rect 12103 9087 12159 9139
rect 12211 9087 12267 9139
rect 12319 9087 13709 9139
rect 11809 9031 13709 9087
rect 11809 8979 12051 9031
rect 12103 8979 12159 9031
rect 12211 8979 12267 9031
rect 12319 8979 13709 9031
rect 11809 8923 13709 8979
rect 11809 8871 12051 8923
rect 12103 8871 12159 8923
rect 12211 8871 12267 8923
rect 12319 8871 13709 8923
rect 11809 8815 13709 8871
rect 11809 8763 12051 8815
rect 12103 8763 12159 8815
rect 12211 8763 12267 8815
rect 12319 8763 13709 8815
rect 11809 8707 13709 8763
rect 11809 8655 12051 8707
rect 12103 8655 12159 8707
rect 12211 8655 12267 8707
rect 12319 8655 13709 8707
rect 11809 8599 13709 8655
rect 11809 8547 12051 8599
rect 12103 8547 12159 8599
rect 12211 8547 12267 8599
rect 12319 8547 13709 8599
rect 11809 8491 13709 8547
rect 11809 8439 12051 8491
rect 12103 8439 12159 8491
rect 12211 8439 12267 8491
rect 12319 8439 13709 8491
rect 11809 8383 13709 8439
rect 11809 8331 12051 8383
rect 12103 8331 12159 8383
rect 12211 8331 12267 8383
rect 12319 8331 13709 8383
rect 11809 8275 13709 8331
rect 11809 8223 12051 8275
rect 12103 8223 12159 8275
rect 12211 8223 12267 8275
rect 12319 8223 13709 8275
rect 11809 8167 13709 8223
rect 11809 8115 12051 8167
rect 12103 8115 12159 8167
rect 12211 8115 12267 8167
rect 12319 8115 13709 8167
rect 11809 8059 13709 8115
rect 11809 8007 12051 8059
rect 12103 8007 12159 8059
rect 12211 8007 12267 8059
rect 12319 8007 13709 8059
rect 11809 7951 13709 8007
rect 11809 7899 12051 7951
rect 12103 7899 12159 7951
rect 12211 7899 12267 7951
rect 12319 7899 13709 7951
rect 11809 7843 13709 7899
rect 11809 7791 12051 7843
rect 12103 7791 12159 7843
rect 12211 7791 12267 7843
rect 12319 7791 13709 7843
rect 11809 7735 13709 7791
rect 11809 7683 12051 7735
rect 12103 7683 12159 7735
rect 12211 7683 12267 7735
rect 12319 7683 13709 7735
rect 11809 7627 13709 7683
rect 11809 7575 12051 7627
rect 12103 7575 12159 7627
rect 12211 7575 12267 7627
rect 12319 7575 13709 7627
rect 11809 7519 13709 7575
rect 11809 7467 12051 7519
rect 12103 7467 12159 7519
rect 12211 7467 12267 7519
rect 12319 7467 13709 7519
rect 11809 7411 13709 7467
rect 11809 7359 12051 7411
rect 12103 7359 12159 7411
rect 12211 7359 12267 7411
rect 12319 7359 13709 7411
rect 11809 7303 13709 7359
rect 11809 7251 12051 7303
rect 12103 7251 12159 7303
rect 12211 7251 12267 7303
rect 12319 7251 13709 7303
rect 11809 7195 13709 7251
rect 11809 7143 12051 7195
rect 12103 7143 12159 7195
rect 12211 7143 12267 7195
rect 12319 7143 13709 7195
rect 11809 7087 13709 7143
rect 11809 7035 12051 7087
rect 12103 7035 12159 7087
rect 12211 7035 12267 7087
rect 12319 7035 13709 7087
rect 11809 6979 13709 7035
rect 11809 6927 12051 6979
rect 12103 6927 12159 6979
rect 12211 6927 12267 6979
rect 12319 6927 13709 6979
rect 11809 6871 13709 6927
rect 11809 6819 12051 6871
rect 12103 6819 12159 6871
rect 12211 6819 12267 6871
rect 12319 6819 13709 6871
rect 11809 6763 13709 6819
rect 11809 6711 12051 6763
rect 12103 6711 12159 6763
rect 12211 6711 12267 6763
rect 12319 6711 13709 6763
rect 11809 6655 13709 6711
rect 11809 6603 12051 6655
rect 12103 6603 12159 6655
rect 12211 6603 12267 6655
rect 12319 6603 13709 6655
rect 11809 6547 13709 6603
rect 11809 6495 12051 6547
rect 12103 6495 12159 6547
rect 12211 6495 12267 6547
rect 12319 6495 13709 6547
rect 11809 6439 13709 6495
rect 11809 6387 12051 6439
rect 12103 6387 12159 6439
rect 12211 6387 12267 6439
rect 12319 6387 13709 6439
rect 11809 6331 13709 6387
rect 11809 6279 12051 6331
rect 12103 6279 12159 6331
rect 12211 6279 12267 6331
rect 12319 6279 13709 6331
rect 11809 6223 13709 6279
rect 11809 6171 12051 6223
rect 12103 6171 12159 6223
rect 12211 6171 12267 6223
rect 12319 6171 13709 6223
rect 11809 6115 13709 6171
rect 11809 6063 12051 6115
rect 12103 6063 12159 6115
rect 12211 6063 12267 6115
rect 12319 6063 13709 6115
rect 11809 6007 13709 6063
rect 11809 5955 12051 6007
rect 12103 5955 12159 6007
rect 12211 5955 12267 6007
rect 12319 5955 13709 6007
rect 11809 5899 13709 5955
rect 11809 5847 12051 5899
rect 12103 5847 12159 5899
rect 12211 5847 12267 5899
rect 12319 5847 13709 5899
rect 11809 5791 13709 5847
rect 11809 5739 12051 5791
rect 12103 5739 12159 5791
rect 12211 5739 12267 5791
rect 12319 5739 13709 5791
rect 11809 5683 13709 5739
rect 11809 5631 12051 5683
rect 12103 5631 12159 5683
rect 12211 5631 12267 5683
rect 12319 5631 13709 5683
rect 11809 5575 13709 5631
rect 11809 5523 12051 5575
rect 12103 5523 12159 5575
rect 12211 5523 12267 5575
rect 12319 5523 13709 5575
rect 11809 5467 13709 5523
rect 11809 5415 12051 5467
rect 12103 5415 12159 5467
rect 12211 5415 12267 5467
rect 12319 5415 13709 5467
rect 11809 5359 13709 5415
rect 11809 5307 12051 5359
rect 12103 5307 12159 5359
rect 12211 5307 12267 5359
rect 12319 5307 13709 5359
rect 11809 5251 13709 5307
rect 11809 5199 12051 5251
rect 12103 5199 12159 5251
rect 12211 5199 12267 5251
rect 12319 5199 13709 5251
rect 11809 5143 13709 5199
rect 11809 5091 12051 5143
rect 12103 5091 12159 5143
rect 12211 5091 12267 5143
rect 12319 5091 13709 5143
rect 11809 5035 13709 5091
rect 11809 4983 12051 5035
rect 12103 4983 12159 5035
rect 12211 4983 12267 5035
rect 12319 4983 13709 5035
rect 11809 4927 13709 4983
rect 11809 4875 12051 4927
rect 12103 4875 12159 4927
rect 12211 4875 12267 4927
rect 12319 4875 13709 4927
rect 11809 4819 13709 4875
rect 11809 4767 12051 4819
rect 12103 4767 12159 4819
rect 12211 4767 12267 4819
rect 12319 4767 13709 4819
rect 11809 4711 13709 4767
rect 11809 4659 12051 4711
rect 12103 4659 12159 4711
rect 12211 4659 12267 4711
rect 12319 4659 13709 4711
rect 11809 4603 13709 4659
rect 11809 4551 12051 4603
rect 12103 4551 12159 4603
rect 12211 4551 12267 4603
rect 12319 4551 13709 4603
rect 11809 4495 13709 4551
rect 11809 4443 12051 4495
rect 12103 4443 12159 4495
rect 12211 4443 12267 4495
rect 12319 4443 13709 4495
rect 11809 4387 13709 4443
rect 11809 4335 12051 4387
rect 12103 4335 12159 4387
rect 12211 4335 12267 4387
rect 12319 4335 13709 4387
rect 11809 4279 13709 4335
rect 11809 4227 12051 4279
rect 12103 4227 12159 4279
rect 12211 4227 12267 4279
rect 12319 4227 13709 4279
rect 11809 4171 13709 4227
rect 11809 4119 12051 4171
rect 12103 4119 12159 4171
rect 12211 4119 12267 4171
rect 12319 4119 13709 4171
rect 11809 4063 13709 4119
rect 11809 4011 12051 4063
rect 12103 4011 12159 4063
rect 12211 4011 12267 4063
rect 12319 4011 13709 4063
rect 11809 3955 13709 4011
rect 11809 3903 12051 3955
rect 12103 3903 12159 3955
rect 12211 3903 12267 3955
rect 12319 3903 13709 3955
rect 11809 3847 13709 3903
rect 11809 3795 12051 3847
rect 12103 3795 12159 3847
rect 12211 3795 12267 3847
rect 12319 3795 13709 3847
rect 11809 3739 13709 3795
rect 11809 3687 12051 3739
rect 12103 3687 12159 3739
rect 12211 3687 12267 3739
rect 12319 3687 13709 3739
rect 11809 3631 13709 3687
rect 11809 3579 12051 3631
rect 12103 3579 12159 3631
rect 12211 3579 12267 3631
rect 12319 3579 13709 3631
rect 11809 3523 13709 3579
rect 11809 3471 12051 3523
rect 12103 3471 12159 3523
rect 12211 3471 12267 3523
rect 12319 3471 13709 3523
rect 11809 3415 13709 3471
rect 11809 3363 12051 3415
rect 12103 3363 12159 3415
rect 12211 3363 12267 3415
rect 12319 3363 13709 3415
rect 11809 3307 13709 3363
rect 11809 3255 12051 3307
rect 12103 3255 12159 3307
rect 12211 3255 12267 3307
rect 12319 3255 13709 3307
rect 11809 3199 13709 3255
rect 11809 3147 12051 3199
rect 12103 3147 12159 3199
rect 12211 3147 12267 3199
rect 12319 3147 13709 3199
rect 11809 3091 13709 3147
rect 11809 3039 12051 3091
rect 12103 3039 12159 3091
rect 12211 3039 12267 3091
rect 12319 3039 13709 3091
rect 11809 2983 13709 3039
rect 11809 2931 12051 2983
rect 12103 2931 12159 2983
rect 12211 2931 12267 2983
rect 12319 2931 13709 2983
rect 11809 2875 13709 2931
rect 11809 2823 12051 2875
rect 12103 2823 12159 2875
rect 12211 2823 12267 2875
rect 12319 2823 13709 2875
rect 11809 2767 13709 2823
rect 11809 2715 12051 2767
rect 12103 2715 12159 2767
rect 12211 2715 12267 2767
rect 12319 2715 13709 2767
rect 11809 2659 13709 2715
rect 11809 2607 12051 2659
rect 12103 2607 12159 2659
rect 12211 2607 12267 2659
rect 12319 2607 13709 2659
rect 11809 2551 13709 2607
rect 11809 2499 12051 2551
rect 12103 2499 12159 2551
rect 12211 2499 12267 2551
rect 12319 2499 13709 2551
rect 11809 2443 13709 2499
rect 11809 2391 12051 2443
rect 12103 2391 12159 2443
rect 12211 2391 12267 2443
rect 12319 2391 13709 2443
rect 11809 2335 13709 2391
rect 11809 2283 12051 2335
rect 12103 2283 12159 2335
rect 12211 2283 12267 2335
rect 12319 2283 13709 2335
rect 11809 2227 13709 2283
rect 11809 2175 12051 2227
rect 12103 2175 12159 2227
rect 12211 2175 12267 2227
rect 12319 2175 13709 2227
rect 11809 2119 13709 2175
rect 11809 2067 12051 2119
rect 12103 2067 12159 2119
rect 12211 2067 12267 2119
rect 12319 2067 13709 2119
rect 11809 2011 13709 2067
rect 11809 1959 12051 2011
rect 12103 1959 12159 2011
rect 12211 1959 12267 2011
rect 12319 1959 13709 2011
rect 11809 1903 13709 1959
rect 11809 1851 12051 1903
rect 12103 1851 12159 1903
rect 12211 1851 12267 1903
rect 12319 1851 13709 1903
rect 11809 1795 13709 1851
rect 11809 1743 12051 1795
rect 12103 1743 12159 1795
rect 12211 1743 12267 1795
rect 12319 1743 13709 1795
rect 11809 1687 13709 1743
rect 11809 1635 12051 1687
rect 12103 1635 12159 1687
rect 12211 1635 12267 1687
rect 12319 1635 13709 1687
rect 11809 1579 13709 1635
rect 11809 1527 12051 1579
rect 12103 1527 12159 1579
rect 12211 1527 12267 1579
rect 12319 1527 13709 1579
rect 11809 1471 13709 1527
rect 11289 309 11309 361
rect 11361 309 11417 361
rect 11469 309 11489 361
rect 11289 253 11489 309
rect 11289 201 11309 253
rect 11361 201 11417 253
rect 11469 201 11489 253
rect 11289 145 11489 201
rect 11289 93 11309 145
rect 11361 93 11417 145
rect 11469 93 11489 145
rect 11289 43 11489 93
rect 11809 1419 12051 1471
rect 12103 1419 12159 1471
rect 12211 1419 12267 1471
rect 12319 1419 13709 1471
rect 11809 1363 13709 1419
rect 11809 1311 12051 1363
rect 12103 1311 12159 1363
rect 12211 1311 12267 1363
rect 12319 1311 13709 1363
rect 11809 1255 13709 1311
rect 11809 1203 12051 1255
rect 12103 1203 12159 1255
rect 12211 1203 12267 1255
rect 12319 1203 13709 1255
rect 11809 1147 13709 1203
rect 11809 1095 12051 1147
rect 12103 1095 12159 1147
rect 12211 1095 12267 1147
rect 12319 1095 13709 1147
rect 11809 1039 13709 1095
rect 11809 987 12051 1039
rect 12103 987 12159 1039
rect 12211 987 12267 1039
rect 12319 987 13709 1039
rect 11809 931 13709 987
rect 11809 879 12051 931
rect 12103 879 12159 931
rect 12211 879 12267 931
rect 12319 879 13709 931
rect 11809 823 13709 879
rect 11809 771 12051 823
rect 12103 771 12159 823
rect 12211 771 12267 823
rect 12319 771 13709 823
rect 11809 715 13709 771
rect 11809 663 12051 715
rect 12103 663 12159 715
rect 12211 663 12267 715
rect 12319 663 13709 715
rect 11809 43 13709 663
use M1_NWELL_CDNS_40661953145131  M1_NWELL_CDNS_40661953145131_0
timestamp 1749760379
transform 1 0 227 0 1 12677
box 0 0 1 1
use M1_NWELL_CDNS_40661953145131  M1_NWELL_CDNS_40661953145131_1
timestamp 1749760379
transform 1 0 12735 0 1 12677
box 0 0 1 1
use M1_NWELL_CDNS_40661953145135  M1_NWELL_CDNS_40661953145135_0
timestamp 1749760379
transform 1 0 6481 0 1 227
box 0 0 1 1
use M1_NWELL_CDNS_40661953145135  M1_NWELL_CDNS_40661953145135_1
timestamp 1749760379
transform 1 0 6481 0 1 25127
box 0 0 1 1
use M1_POLY2_CDNS_40661953145132  M1_POLY2_CDNS_40661953145132_0
timestamp 1749760379
transform -1 0 11633 0 1 3869
box 0 0 1 1
use M1_POLY2_CDNS_40661953145132  M1_POLY2_CDNS_40661953145132_1
timestamp 1749760379
transform -1 0 11633 0 1 9741
box 0 0 1 1
use M1_POLY2_CDNS_40661953145132  M1_POLY2_CDNS_40661953145132_2
timestamp 1749760379
transform 1 0 1329 0 1 3869
box 0 0 1 1
use M1_POLY2_CDNS_40661953145132  M1_POLY2_CDNS_40661953145132_3
timestamp 1749760379
transform 1 0 1329 0 1 9741
box 0 0 1 1
use M1_POLY2_CDNS_40661953145132  M1_POLY2_CDNS_40661953145132_4
timestamp 1749760379
transform 1 0 1329 0 1 15613
box 0 0 1 1
use M1_POLY2_CDNS_40661953145132  M1_POLY2_CDNS_40661953145132_5
timestamp 1749760379
transform 1 0 1329 0 1 21485
box 0 0 1 1
use M1_POLY2_CDNS_40661953145132  M1_POLY2_CDNS_40661953145132_6
timestamp 1749760379
transform -1 0 11633 0 1 15613
box 0 0 1 1
use M1_POLY2_CDNS_40661953145132  M1_POLY2_CDNS_40661953145132_7
timestamp 1749760379
transform -1 0 11633 0 1 21485
box 0 0 1 1
use M1_PSUB_CDNS_40661953145130  M1_PSUB_CDNS_40661953145130_0
timestamp 1749760379
transform 1 0 6481 0 1 6805
box 0 0 1 1
use M1_PSUB_CDNS_40661953145130  M1_PSUB_CDNS_40661953145130_1
timestamp 1749760379
transform 1 0 6481 0 1 12677
box 0 0 1 1
use M1_PSUB_CDNS_40661953145130  M1_PSUB_CDNS_40661953145130_2
timestamp 1749760379
transform 1 0 6481 0 1 18549
box 0 0 1 1
use M1_PSUB_CDNS_40661953145133  M1_PSUB_CDNS_40661953145133_0
timestamp 1749760379
transform 1 0 12185 0 1 12677
box 0 0 1 1
use M1_PSUB_CDNS_40661953145133  M1_PSUB_CDNS_40661953145133_1
timestamp 1749760379
transform 1 0 777 0 1 12677
box 0 0 1 1
use M1_PSUB_CDNS_40661953145134  M1_PSUB_CDNS_40661953145134_0
timestamp 1749760379
transform 1 0 6481 0 1 24527
box 0 0 1 1
use M1_PSUB_CDNS_40661953145134  M1_PSUB_CDNS_40661953145134_1
timestamp 1749760379
transform 1 0 6481 0 1 827
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_0
timestamp 1749760379
transform -1 0 11389 0 1 227
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_1
timestamp 1749760379
transform -1 0 9019 0 1 227
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_2
timestamp 1749760379
transform -1 0 3943 0 1 227
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_3
timestamp 1749760379
transform 1 0 1573 0 1 227
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_4
timestamp 1749760379
transform -1 0 3943 0 1 25127
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_5
timestamp 1749760379
transform 1 0 1573 0 1 25127
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_6
timestamp 1749760379
transform -1 0 9019 0 1 25127
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_7
timestamp 1749760379
transform -1 0 11389 0 1 25127
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_0
timestamp 1749760379
transform 1 0 6481 0 1 25127
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_1
timestamp 1749760379
transform 1 0 6481 0 1 227
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_0
timestamp 1749760379
transform 1 0 6481 0 1 6065
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_1
timestamp 1749760379
transform 1 0 6481 0 1 11449
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_2
timestamp 1749760379
transform 1 0 6481 0 1 10961
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_3
timestamp 1749760379
transform 1 0 6481 0 1 10473
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_4
timestamp 1749760379
transform 1 0 6481 0 1 9985
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_5
timestamp 1749760379
transform 1 0 6481 0 1 9497
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_6
timestamp 1749760379
transform 1 0 6481 0 1 9009
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_7
timestamp 1749760379
transform 1 0 6481 0 1 8033
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_8
timestamp 1749760379
transform 1 0 6481 0 1 7545
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_9
timestamp 1749760379
transform 1 0 6481 0 1 5577
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_10
timestamp 1749760379
transform 1 0 6481 0 1 5089
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_11
timestamp 1749760379
transform 1 0 6481 0 1 4601
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_12
timestamp 1749760379
transform 1 0 6481 0 1 4113
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_13
timestamp 1749760379
transform 1 0 6481 0 1 3625
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_14
timestamp 1749760379
transform 1 0 6481 0 1 3137
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_15
timestamp 1749760379
transform 1 0 6481 0 1 2649
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_16
timestamp 1749760379
transform 1 0 6481 0 1 2161
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_17
timestamp 1749760379
transform 1 0 6481 0 1 1673
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_18
timestamp 1749760379
transform 1 0 6481 0 1 13417
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_19
timestamp 1749760379
transform 1 0 6481 0 1 11937
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_20
timestamp 1749760379
transform 1 0 6481 0 1 23681
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_21
timestamp 1749760379
transform 1 0 6481 0 1 23193
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_22
timestamp 1749760379
transform 1 0 6481 0 1 22705
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_23
timestamp 1749760379
transform 1 0 6481 0 1 22217
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_24
timestamp 1749760379
transform 1 0 6481 0 1 21729
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_25
timestamp 1749760379
transform 1 0 6481 0 1 21241
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_26
timestamp 1749760379
transform 1 0 6481 0 1 20753
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_27
timestamp 1749760379
transform 1 0 6481 0 1 20265
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_28
timestamp 1749760379
transform 1 0 6481 0 1 19777
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_29
timestamp 1749760379
transform 1 0 6481 0 1 19289
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_30
timestamp 1749760379
transform 1 0 6481 0 1 17809
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_31
timestamp 1749760379
transform 1 0 6481 0 1 17321
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_32
timestamp 1749760379
transform 1 0 6481 0 1 8521
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_33
timestamp 1749760379
transform 1 0 6481 0 1 16833
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_34
timestamp 1749760379
transform 1 0 6481 0 1 16345
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_35
timestamp 1749760379
transform 1 0 6481 0 1 15857
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_36
timestamp 1749760379
transform 1 0 6481 0 1 15369
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_37
timestamp 1749760379
transform 1 0 6481 0 1 14881
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_38
timestamp 1749760379
transform 1 0 6481 0 1 14393
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_39
timestamp 1749760379
transform 1 0 6481 0 1 13905
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_0
timestamp 1749760379
transform -1 0 11389 0 1 5577
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_1
timestamp 1749760379
transform -1 0 11389 0 1 6065
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_2
timestamp 1749760379
transform -1 0 11389 0 1 7545
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_3
timestamp 1749760379
transform -1 0 11389 0 1 8033
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_4
timestamp 1749760379
transform -1 0 11389 0 1 8521
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_5
timestamp 1749760379
transform -1 0 11389 0 1 9009
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_6
timestamp 1749760379
transform -1 0 11389 0 1 9497
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_7
timestamp 1749760379
transform -1 0 11389 0 1 9985
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_8
timestamp 1749760379
transform -1 0 11389 0 1 10473
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_9
timestamp 1749760379
transform -1 0 11389 0 1 10961
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_10
timestamp 1749760379
transform -1 0 9019 0 1 7545
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_11
timestamp 1749760379
transform -1 0 11389 0 1 11937
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_12
timestamp 1749760379
transform -1 0 9019 0 1 3137
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_13
timestamp 1749760379
transform -1 0 9019 0 1 2649
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_14
timestamp 1749760379
transform -1 0 9019 0 1 2161
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_15
timestamp 1749760379
transform -1 0 9019 0 1 1673
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_16
timestamp 1749760379
transform -1 0 9019 0 1 6065
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_17
timestamp 1749760379
transform -1 0 9019 0 1 8033
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_18
timestamp 1749760379
transform -1 0 9019 0 1 8521
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_19
timestamp 1749760379
transform -1 0 9019 0 1 9009
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_20
timestamp 1749760379
transform -1 0 9019 0 1 9497
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_21
timestamp 1749760379
transform -1 0 9019 0 1 9985
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_22
timestamp 1749760379
transform -1 0 11389 0 1 2649
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_23
timestamp 1749760379
transform -1 0 11389 0 1 2161
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_24
timestamp 1749760379
transform -1 0 11389 0 1 1673
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_25
timestamp 1749760379
transform -1 0 9019 0 1 10473
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_26
timestamp 1749760379
transform -1 0 11389 0 1 11449
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_27
timestamp 1749760379
transform -1 0 9019 0 1 10961
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_28
timestamp 1749760379
transform -1 0 9019 0 1 11449
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_29
timestamp 1749760379
transform -1 0 9019 0 1 11937
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_30
timestamp 1749760379
transform -1 0 9019 0 1 5577
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_31
timestamp 1749760379
transform -1 0 9019 0 1 5089
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_32
timestamp 1749760379
transform -1 0 9019 0 1 4601
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_33
timestamp 1749760379
transform -1 0 9019 0 1 4113
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_34
timestamp 1749760379
transform -1 0 9019 0 1 3625
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_35
timestamp 1749760379
transform -1 0 11389 0 1 3137
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_36
timestamp 1749760379
transform -1 0 11389 0 1 3625
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_37
timestamp 1749760379
transform -1 0 11389 0 1 4113
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_38
timestamp 1749760379
transform -1 0 11389 0 1 4601
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_39
timestamp 1749760379
transform -1 0 11389 0 1 5089
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_40
timestamp 1749760379
transform 1 0 1573 0 1 9009
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_41
timestamp 1749760379
transform 1 0 1573 0 1 8033
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_42
timestamp 1749760379
transform 1 0 1573 0 1 6065
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_43
timestamp 1749760379
transform 1 0 1573 0 1 5577
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_44
timestamp 1749760379
transform 1 0 1573 0 1 5089
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_45
timestamp 1749760379
transform 1 0 1573 0 1 4601
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_46
timestamp 1749760379
transform 1 0 1573 0 1 4113
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_47
timestamp 1749760379
transform -1 0 3943 0 1 1673
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_48
timestamp 1749760379
transform 1 0 1573 0 1 3625
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_49
timestamp 1749760379
transform -1 0 3943 0 1 2161
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_50
timestamp 1749760379
transform -1 0 3943 0 1 2649
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_51
timestamp 1749760379
transform -1 0 3943 0 1 3137
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_52
timestamp 1749760379
transform -1 0 3943 0 1 3625
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_53
timestamp 1749760379
transform -1 0 3943 0 1 4113
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_54
timestamp 1749760379
transform -1 0 3943 0 1 4601
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_55
timestamp 1749760379
transform -1 0 3943 0 1 5089
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_56
timestamp 1749760379
transform -1 0 3943 0 1 5577
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_57
timestamp 1749760379
transform -1 0 3943 0 1 6065
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_58
timestamp 1749760379
transform -1 0 3943 0 1 7545
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_59
timestamp 1749760379
transform -1 0 3943 0 1 8033
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_60
timestamp 1749760379
transform -1 0 3943 0 1 8521
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_61
timestamp 1749760379
transform -1 0 3943 0 1 9009
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_62
timestamp 1749760379
transform -1 0 3943 0 1 9985
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_63
timestamp 1749760379
transform -1 0 3943 0 1 10473
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_64
timestamp 1749760379
transform -1 0 3943 0 1 10961
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_65
timestamp 1749760379
transform -1 0 3943 0 1 11449
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_66
timestamp 1749760379
transform -1 0 3943 0 1 11937
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_67
timestamp 1749760379
transform 1 0 1573 0 1 3137
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_68
timestamp 1749760379
transform 1 0 1573 0 1 2649
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_69
timestamp 1749760379
transform 1 0 1573 0 1 2161
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_70
timestamp 1749760379
transform 1 0 1573 0 1 1673
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_71
timestamp 1749760379
transform 1 0 1573 0 1 7545
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_72
timestamp 1749760379
transform 1 0 1573 0 1 8521
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_73
timestamp 1749760379
transform 1 0 1573 0 1 11937
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_74
timestamp 1749760379
transform 1 0 1573 0 1 11449
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_75
timestamp 1749760379
transform 1 0 1573 0 1 10961
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_76
timestamp 1749760379
transform -1 0 3943 0 1 9497
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_77
timestamp 1749760379
transform 1 0 1573 0 1 10473
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_78
timestamp 1749760379
transform 1 0 1573 0 1 9985
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_79
timestamp 1749760379
transform 1 0 1573 0 1 9497
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_80
timestamp 1749760379
transform -1 0 3943 0 1 22705
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_81
timestamp 1749760379
transform -1 0 3943 0 1 22217
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_82
timestamp 1749760379
transform -1 0 3943 0 1 21729
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_83
timestamp 1749760379
transform -1 0 3943 0 1 21241
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_84
timestamp 1749760379
transform -1 0 3943 0 1 20753
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_85
timestamp 1749760379
transform -1 0 3943 0 1 20265
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_86
timestamp 1749760379
transform -1 0 3943 0 1 19289
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_87
timestamp 1749760379
transform -1 0 3943 0 1 19777
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_88
timestamp 1749760379
transform -1 0 3943 0 1 13417
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_89
timestamp 1749760379
transform -1 0 3943 0 1 13905
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_90
timestamp 1749760379
transform -1 0 3943 0 1 14393
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_91
timestamp 1749760379
transform -1 0 3943 0 1 14881
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_92
timestamp 1749760379
transform -1 0 3943 0 1 15369
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_93
timestamp 1749760379
transform -1 0 3943 0 1 15857
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_94
timestamp 1749760379
transform -1 0 3943 0 1 16345
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_95
timestamp 1749760379
transform -1 0 3943 0 1 16833
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_96
timestamp 1749760379
transform -1 0 3943 0 1 17321
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_97
timestamp 1749760379
transform -1 0 3943 0 1 17809
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_98
timestamp 1749760379
transform 1 0 1573 0 1 22217
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_99
timestamp 1749760379
transform 1 0 1573 0 1 19777
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_100
timestamp 1749760379
transform 1 0 1573 0 1 20753
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_101
timestamp 1749760379
transform 1 0 1573 0 1 22705
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_102
timestamp 1749760379
transform 1 0 1573 0 1 19289
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_103
timestamp 1749760379
transform 1 0 1573 0 1 20265
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_104
timestamp 1749760379
transform 1 0 1573 0 1 13417
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_105
timestamp 1749760379
transform 1 0 1573 0 1 21241
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_106
timestamp 1749760379
transform 1 0 1573 0 1 21729
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_107
timestamp 1749760379
transform 1 0 1573 0 1 17809
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_108
timestamp 1749760379
transform 1 0 1573 0 1 17321
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_109
timestamp 1749760379
transform 1 0 1573 0 1 16833
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_110
timestamp 1749760379
transform 1 0 1573 0 1 16345
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_111
timestamp 1749760379
transform 1 0 1573 0 1 15857
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_112
timestamp 1749760379
transform 1 0 1573 0 1 15369
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_113
timestamp 1749760379
transform 1 0 1573 0 1 14881
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_114
timestamp 1749760379
transform 1 0 1573 0 1 14393
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_115
timestamp 1749760379
transform 1 0 1573 0 1 13905
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_116
timestamp 1749760379
transform 1 0 1573 0 1 23681
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_117
timestamp 1749760379
transform 1 0 1573 0 1 23193
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_118
timestamp 1749760379
transform -1 0 3943 0 1 23681
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_119
timestamp 1749760379
transform -1 0 3943 0 1 23193
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_120
timestamp 1749760379
transform -1 0 11389 0 1 15369
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_121
timestamp 1749760379
transform -1 0 11389 0 1 15857
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_122
timestamp 1749760379
transform -1 0 11389 0 1 16345
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_123
timestamp 1749760379
transform -1 0 11389 0 1 16833
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_124
timestamp 1749760379
transform -1 0 11389 0 1 17321
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_125
timestamp 1749760379
transform -1 0 11389 0 1 17809
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_126
timestamp 1749760379
transform -1 0 11389 0 1 19289
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_127
timestamp 1749760379
transform -1 0 11389 0 1 19777
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_128
timestamp 1749760379
transform -1 0 11389 0 1 20265
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_129
timestamp 1749760379
transform -1 0 11389 0 1 20753
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_130
timestamp 1749760379
transform -1 0 11389 0 1 23681
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_131
timestamp 1749760379
transform -1 0 11389 0 1 23193
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_132
timestamp 1749760379
transform -1 0 11389 0 1 22705
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_133
timestamp 1749760379
transform -1 0 11389 0 1 21729
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_134
timestamp 1749760379
transform -1 0 11389 0 1 21241
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_135
timestamp 1749760379
transform -1 0 9019 0 1 13417
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_136
timestamp 1749760379
transform -1 0 9019 0 1 13905
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_137
timestamp 1749760379
transform -1 0 9019 0 1 14393
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_138
timestamp 1749760379
transform -1 0 9019 0 1 14881
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_139
timestamp 1749760379
transform -1 0 9019 0 1 15369
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_140
timestamp 1749760379
transform -1 0 9019 0 1 16345
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_141
timestamp 1749760379
transform -1 0 9019 0 1 16833
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_142
timestamp 1749760379
transform -1 0 9019 0 1 17321
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_143
timestamp 1749760379
transform -1 0 9019 0 1 17809
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_144
timestamp 1749760379
transform -1 0 9019 0 1 19289
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_145
timestamp 1749760379
transform -1 0 9019 0 1 19777
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_146
timestamp 1749760379
transform -1 0 9019 0 1 20265
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_147
timestamp 1749760379
transform -1 0 9019 0 1 20753
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_148
timestamp 1749760379
transform -1 0 9019 0 1 21241
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_149
timestamp 1749760379
transform -1 0 9019 0 1 21729
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_150
timestamp 1749760379
transform -1 0 9019 0 1 22217
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_151
timestamp 1749760379
transform -1 0 9019 0 1 22705
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_152
timestamp 1749760379
transform -1 0 9019 0 1 23193
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_153
timestamp 1749760379
transform -1 0 9019 0 1 23681
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_154
timestamp 1749760379
transform -1 0 9019 0 1 15857
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_155
timestamp 1749760379
transform -1 0 11389 0 1 13417
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_156
timestamp 1749760379
transform -1 0 11389 0 1 22217
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_157
timestamp 1749760379
transform -1 0 11389 0 1 13905
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_158
timestamp 1749760379
transform -1 0 11389 0 1 14393
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_159
timestamp 1749760379
transform -1 0 11389 0 1 14881
box 0 0 1 1
use M2_M1_CDNS_40661953145136  M2_M1_CDNS_40661953145136_0
timestamp 1749760379
transform 1 0 11649 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661953145136  M2_M1_CDNS_40661953145136_1
timestamp 1749760379
transform 1 0 11649 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661953145136  M2_M1_CDNS_40661953145136_2
timestamp 1749760379
transform 1 0 1313 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661953145136  M2_M1_CDNS_40661953145136_3
timestamp 1749760379
transform 1 0 1313 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661953145136  M2_M1_CDNS_40661953145136_4
timestamp 1749760379
transform 1 0 1313 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661953145136  M2_M1_CDNS_40661953145136_5
timestamp 1749760379
transform 1 0 1313 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661953145136  M2_M1_CDNS_40661953145136_6
timestamp 1749760379
transform 1 0 11649 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661953145136  M2_M1_CDNS_40661953145136_7
timestamp 1749760379
transform 1 0 11649 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661953145138  M2_M1_CDNS_40661953145138_0
timestamp 1749760379
transform -1 0 10204 0 1 827
box 0 0 1 1
use M2_M1_CDNS_40661953145138  M2_M1_CDNS_40661953145138_1
timestamp 1749760379
transform -1 0 7834 0 1 827
box 0 0 1 1
use M2_M1_CDNS_40661953145138  M2_M1_CDNS_40661953145138_2
timestamp 1749760379
transform 1 0 2758 0 1 827
box 0 0 1 1
use M2_M1_CDNS_40661953145138  M2_M1_CDNS_40661953145138_3
timestamp 1749760379
transform 1 0 5128 0 1 827
box 0 0 1 1
use M2_M1_CDNS_40661953145138  M2_M1_CDNS_40661953145138_4
timestamp 1749760379
transform 1 0 5128 0 1 24527
box 0 0 1 1
use M2_M1_CDNS_40661953145138  M2_M1_CDNS_40661953145138_5
timestamp 1749760379
transform 1 0 2758 0 1 24527
box 0 0 1 1
use M2_M1_CDNS_40661953145138  M2_M1_CDNS_40661953145138_6
timestamp 1749760379
transform -1 0 7834 0 1 24527
box 0 0 1 1
use M2_M1_CDNS_40661953145138  M2_M1_CDNS_40661953145138_7
timestamp 1749760379
transform -1 0 10204 0 1 24527
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_0
timestamp 1749760379
transform -1 0 10204 0 1 10717
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_1
timestamp 1749760379
transform -1 0 10204 0 1 10229
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_2
timestamp 1749760379
transform -1 0 10204 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_3
timestamp 1749760379
transform -1 0 10204 0 1 9253
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_4
timestamp 1749760379
transform -1 0 10204 0 1 8765
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_5
timestamp 1749760379
transform -1 0 10204 0 1 8277
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_6
timestamp 1749760379
transform -1 0 10204 0 1 7789
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_7
timestamp 1749760379
transform -1 0 10204 0 1 7301
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_8
timestamp 1749760379
transform -1 0 10204 0 1 6309
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_9
timestamp 1749760379
transform -1 0 10204 0 1 5821
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_10
timestamp 1749760379
transform -1 0 10204 0 1 11205
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_11
timestamp 1749760379
transform -1 0 10204 0 1 4845
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_12
timestamp 1749760379
transform -1 0 10204 0 1 4357
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_13
timestamp 1749760379
transform -1 0 10204 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_14
timestamp 1749760379
transform -1 0 10204 0 1 3381
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_15
timestamp 1749760379
transform -1 0 10204 0 1 2893
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_16
timestamp 1749760379
transform -1 0 10204 0 1 2405
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_17
timestamp 1749760379
transform -1 0 10204 0 1 1917
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_18
timestamp 1749760379
transform -1 0 10204 0 1 1429
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_19
timestamp 1749760379
transform -1 0 7834 0 1 1917
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_20
timestamp 1749760379
transform -1 0 10204 0 1 5333
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_21
timestamp 1749760379
transform -1 0 10204 0 1 11693
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_22
timestamp 1749760379
transform -1 0 10204 0 1 12181
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_23
timestamp 1749760379
transform -1 0 7834 0 1 8277
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_24
timestamp 1749760379
transform -1 0 7834 0 1 8765
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_25
timestamp 1749760379
transform -1 0 7834 0 1 9253
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_26
timestamp 1749760379
transform -1 0 7834 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_27
timestamp 1749760379
transform -1 0 7834 0 1 10229
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_28
timestamp 1749760379
transform -1 0 7834 0 1 10717
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_29
timestamp 1749760379
transform -1 0 7834 0 1 11205
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_30
timestamp 1749760379
transform -1 0 7834 0 1 11693
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_31
timestamp 1749760379
transform -1 0 7834 0 1 12181
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_32
timestamp 1749760379
transform -1 0 7834 0 1 1429
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_33
timestamp 1749760379
transform -1 0 7834 0 1 2405
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_34
timestamp 1749760379
transform -1 0 7834 0 1 2893
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_35
timestamp 1749760379
transform -1 0 7834 0 1 3381
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_36
timestamp 1749760379
transform -1 0 7834 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_37
timestamp 1749760379
transform -1 0 7834 0 1 4357
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_38
timestamp 1749760379
transform -1 0 7834 0 1 4845
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_39
timestamp 1749760379
transform -1 0 7834 0 1 5333
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_40
timestamp 1749760379
transform -1 0 7834 0 1 5821
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_41
timestamp 1749760379
transform -1 0 7834 0 1 6309
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_42
timestamp 1749760379
transform -1 0 7834 0 1 7789
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_43
timestamp 1749760379
transform -1 0 7834 0 1 7301
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_44
timestamp 1749760379
transform 1 0 5128 0 1 4845
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_45
timestamp 1749760379
transform 1 0 2758 0 1 12181
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_46
timestamp 1749760379
transform 1 0 5128 0 1 1429
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_47
timestamp 1749760379
transform 1 0 2758 0 1 6309
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_48
timestamp 1749760379
transform 1 0 2758 0 1 7301
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_49
timestamp 1749760379
transform 1 0 2758 0 1 7789
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_50
timestamp 1749760379
transform 1 0 2758 0 1 8277
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_51
timestamp 1749760379
transform 1 0 2758 0 1 8765
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_52
timestamp 1749760379
transform 1 0 2758 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_53
timestamp 1749760379
transform 1 0 2758 0 1 10229
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_54
timestamp 1749760379
transform 1 0 2758 0 1 11205
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_55
timestamp 1749760379
transform 1 0 2758 0 1 11693
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_56
timestamp 1749760379
transform 1 0 2758 0 1 1429
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_57
timestamp 1749760379
transform 1 0 2758 0 1 1917
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_58
timestamp 1749760379
transform 1 0 2758 0 1 2405
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_59
timestamp 1749760379
transform 1 0 2758 0 1 2893
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_60
timestamp 1749760379
transform 1 0 2758 0 1 3381
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_61
timestamp 1749760379
transform 1 0 2758 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_62
timestamp 1749760379
transform 1 0 2758 0 1 4357
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_63
timestamp 1749760379
transform 1 0 2758 0 1 4845
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_64
timestamp 1749760379
transform 1 0 2758 0 1 5333
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_65
timestamp 1749760379
transform 1 0 2758 0 1 10717
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_66
timestamp 1749760379
transform 1 0 5128 0 1 8277
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_67
timestamp 1749760379
transform 1 0 5128 0 1 8765
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_68
timestamp 1749760379
transform 1 0 5128 0 1 9253
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_69
timestamp 1749760379
transform 1 0 5128 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_70
timestamp 1749760379
transform 1 0 5128 0 1 10229
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_71
timestamp 1749760379
transform 1 0 5128 0 1 10717
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_72
timestamp 1749760379
transform 1 0 5128 0 1 11205
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_73
timestamp 1749760379
transform 1 0 5128 0 1 11693
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_74
timestamp 1749760379
transform 1 0 5128 0 1 12181
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_75
timestamp 1749760379
transform 1 0 5128 0 1 7789
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_76
timestamp 1749760379
transform 1 0 2758 0 1 9253
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_77
timestamp 1749760379
transform 1 0 2758 0 1 5821
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_78
timestamp 1749760379
transform 1 0 5128 0 1 7301
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_79
timestamp 1749760379
transform 1 0 5128 0 1 6309
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_80
timestamp 1749760379
transform 1 0 5128 0 1 5821
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_81
timestamp 1749760379
transform 1 0 5128 0 1 5333
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_82
timestamp 1749760379
transform 1 0 5128 0 1 1917
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_83
timestamp 1749760379
transform 1 0 5128 0 1 2405
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_84
timestamp 1749760379
transform 1 0 5128 0 1 2893
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_85
timestamp 1749760379
transform 1 0 5128 0 1 3381
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_86
timestamp 1749760379
transform 1 0 5128 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_87
timestamp 1749760379
transform 1 0 5128 0 1 4357
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_88
timestamp 1749760379
transform 1 0 2758 0 1 19045
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_89
timestamp 1749760379
transform 1 0 5128 0 1 13173
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_90
timestamp 1749760379
transform 1 0 5128 0 1 14149
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_91
timestamp 1749760379
transform 1 0 5128 0 1 14637
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_92
timestamp 1749760379
transform 1 0 5128 0 1 15125
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_93
timestamp 1749760379
transform 1 0 5128 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_94
timestamp 1749760379
transform 1 0 5128 0 1 16101
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_95
timestamp 1749760379
transform 1 0 5128 0 1 22949
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_96
timestamp 1749760379
transform 1 0 2758 0 1 23437
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_97
timestamp 1749760379
transform 1 0 5128 0 1 22461
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_98
timestamp 1749760379
transform 1 0 5128 0 1 13661
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_99
timestamp 1749760379
transform 1 0 2758 0 1 20509
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_100
timestamp 1749760379
transform 1 0 2758 0 1 20997
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_101
timestamp 1749760379
transform 1 0 2758 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_102
timestamp 1749760379
transform 1 0 2758 0 1 21973
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_103
timestamp 1749760379
transform 1 0 2758 0 1 22461
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_104
timestamp 1749760379
transform 1 0 2758 0 1 22949
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_105
timestamp 1749760379
transform 1 0 5128 0 1 16589
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_106
timestamp 1749760379
transform 1 0 5128 0 1 17077
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_107
timestamp 1749760379
transform 1 0 5128 0 1 17565
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_108
timestamp 1749760379
transform 1 0 5128 0 1 18053
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_109
timestamp 1749760379
transform 1 0 5128 0 1 19045
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_110
timestamp 1749760379
transform 1 0 2758 0 1 20021
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_111
timestamp 1749760379
transform 1 0 5128 0 1 21973
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_112
timestamp 1749760379
transform 1 0 5128 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_113
timestamp 1749760379
transform 1 0 5128 0 1 20997
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_114
timestamp 1749760379
transform 1 0 5128 0 1 20509
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_115
timestamp 1749760379
transform 1 0 5128 0 1 20021
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_116
timestamp 1749760379
transform 1 0 5128 0 1 19533
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_117
timestamp 1749760379
transform 1 0 2758 0 1 13661
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_118
timestamp 1749760379
transform 1 0 2758 0 1 13173
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_119
timestamp 1749760379
transform 1 0 2758 0 1 14149
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_120
timestamp 1749760379
transform 1 0 2758 0 1 14637
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_121
timestamp 1749760379
transform 1 0 2758 0 1 15125
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_122
timestamp 1749760379
transform 1 0 2758 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_123
timestamp 1749760379
transform 1 0 2758 0 1 16101
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_124
timestamp 1749760379
transform 1 0 2758 0 1 16589
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_125
timestamp 1749760379
transform 1 0 2758 0 1 17077
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_126
timestamp 1749760379
transform 1 0 2758 0 1 17565
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_127
timestamp 1749760379
transform 1 0 2758 0 1 18053
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_128
timestamp 1749760379
transform 1 0 2758 0 1 23925
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_129
timestamp 1749760379
transform 1 0 2758 0 1 19533
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_130
timestamp 1749760379
transform 1 0 5128 0 1 23437
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_131
timestamp 1749760379
transform 1 0 5128 0 1 23925
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_132
timestamp 1749760379
transform -1 0 7834 0 1 19045
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_133
timestamp 1749760379
transform -1 0 10204 0 1 18053
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_134
timestamp 1749760379
transform -1 0 10204 0 1 23925
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_135
timestamp 1749760379
transform -1 0 10204 0 1 23437
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_136
timestamp 1749760379
transform -1 0 10204 0 1 22949
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_137
timestamp 1749760379
transform -1 0 10204 0 1 22461
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_138
timestamp 1749760379
transform -1 0 10204 0 1 21973
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_139
timestamp 1749760379
transform -1 0 10204 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_140
timestamp 1749760379
transform -1 0 10204 0 1 20997
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_141
timestamp 1749760379
transform -1 0 10204 0 1 20509
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_142
timestamp 1749760379
transform -1 0 10204 0 1 20021
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_143
timestamp 1749760379
transform -1 0 10204 0 1 19045
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_144
timestamp 1749760379
transform -1 0 7834 0 1 13661
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_145
timestamp 1749760379
transform -1 0 7834 0 1 14149
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_146
timestamp 1749760379
transform -1 0 7834 0 1 14637
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_147
timestamp 1749760379
transform -1 0 7834 0 1 15125
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_148
timestamp 1749760379
transform -1 0 7834 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_149
timestamp 1749760379
transform -1 0 7834 0 1 16101
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_150
timestamp 1749760379
transform -1 0 7834 0 1 16589
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_151
timestamp 1749760379
transform -1 0 7834 0 1 17077
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_152
timestamp 1749760379
transform -1 0 7834 0 1 17565
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_153
timestamp 1749760379
transform -1 0 7834 0 1 18053
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_154
timestamp 1749760379
transform -1 0 10204 0 1 19533
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_155
timestamp 1749760379
transform -1 0 7834 0 1 13173
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_156
timestamp 1749760379
transform -1 0 10204 0 1 16101
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_157
timestamp 1749760379
transform -1 0 10204 0 1 17077
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_158
timestamp 1749760379
transform -1 0 10204 0 1 16589
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_159
timestamp 1749760379
transform -1 0 10204 0 1 17565
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_160
timestamp 1749760379
transform -1 0 10204 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_161
timestamp 1749760379
transform -1 0 10204 0 1 15125
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_162
timestamp 1749760379
transform -1 0 10204 0 1 14637
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_163
timestamp 1749760379
transform -1 0 10204 0 1 14149
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_164
timestamp 1749760379
transform -1 0 10204 0 1 13661
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_165
timestamp 1749760379
transform -1 0 10204 0 1 13173
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_166
timestamp 1749760379
transform -1 0 7834 0 1 19533
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_167
timestamp 1749760379
transform -1 0 7834 0 1 23925
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_168
timestamp 1749760379
transform -1 0 7834 0 1 23437
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_169
timestamp 1749760379
transform -1 0 7834 0 1 22949
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_170
timestamp 1749760379
transform -1 0 7834 0 1 22461
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_171
timestamp 1749760379
transform -1 0 7834 0 1 21973
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_172
timestamp 1749760379
transform -1 0 7834 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_173
timestamp 1749760379
transform -1 0 7834 0 1 20997
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_174
timestamp 1749760379
transform -1 0 7834 0 1 20509
box 0 0 1 1
use M2_M1_CDNS_40661953145140  M2_M1_CDNS_40661953145140_175
timestamp 1749760379
transform -1 0 7834 0 1 20021
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_0
timestamp 1749760379
transform -1 0 10204 0 1 6805
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_1
timestamp 1749760379
transform -1 0 7834 0 1 6805
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_2
timestamp 1749760379
transform 1 0 2758 0 1 6805
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_3
timestamp 1749760379
transform 1 0 5128 0 1 6805
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_4
timestamp 1749760379
transform 1 0 2758 0 1 18549
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_5
timestamp 1749760379
transform 1 0 5128 0 1 18549
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_6
timestamp 1749760379
transform -1 0 10204 0 1 18549
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_7
timestamp 1749760379
transform -1 0 7834 0 1 18549
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_8
timestamp 1749760379
transform -1 0 7834 0 1 12677
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_9
timestamp 1749760379
transform -1 0 10204 0 1 12677
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_10
timestamp 1749760379
transform 1 0 5128 0 1 12677
box 0 0 1 1
use M2_M1_CDNS_40661953145146  M2_M1_CDNS_40661953145146_11
timestamp 1749760379
transform 1 0 2758 0 1 12677
box 0 0 1 1
use M2_M1_CDNS_40661953145162  M2_M1_CDNS_40661953145162_0
timestamp 1749760379
transform 1 0 12185 0 1 12677
box 0 0 1 1
use M2_M1_CDNS_40661953145162  M2_M1_CDNS_40661953145162_1
timestamp 1749760379
transform 1 0 777 0 1 12677
box 0 0 1 1
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_0
timestamp 1749760379
transform 0 -1 11481 1 0 7353
box 0 0 1 1
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_1
timestamp 1749760379
transform 0 -1 11481 1 0 13225
box 0 0 1 1
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_2
timestamp 1749760379
transform 0 -1 11481 1 0 1481
box 0 0 1 1
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_3
timestamp 1749760379
transform 0 -1 11481 1 0 19097
box 0 0 1 1
<< properties >>
string GDS_END 4937384
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4892910
string path 32.825 165.850 32.825 27.450 
<< end >>
