magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
use M1_NWELL$$46277676_64x8m81_0  M1_NWELL$$46277676_64x8m81_0_0
timestamp 1749760379
transform 1 0 310 0 1 12142
box 0 0 1 1
use M1_NWELL$$47121452_64x8m81_0  M1_NWELL$$47121452_64x8m81_0_0
timestamp 1749760379
transform 1 0 237 0 1 1392
box 0 0 1 1
use M1_PACTIVE4310589983248_64x8m81  M1_PACTIVE4310589983248_64x8m81_0
timestamp 1749760379
transform 1 0 244 0 1 141
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_0
timestamp 1749760379
transform 1 0 310 0 1 3446
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_1
timestamp 1749760379
transform 1 0 310 0 1 3169
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_2
timestamp 1749760379
transform 1 0 253 0 1 1202
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_3
timestamp 1749760379
transform 1 0 310 0 1 7144
box 0 0 1 1
use M1_POLY24310589983237_64x8m81  M1_POLY24310589983237_64x8m81_0
timestamp 1749760379
transform 1 0 304 0 1 10311
box 0 0 1 1
use M1_PSUB$$45111340_64x8m81_0  M1_PSUB$$45111340_64x8m81_0_0
timestamp 1749760379
transform 1 0 0 0 1 5237
box 0 0 1 1
use M2_M1$$46894124_64x8m81_0  M2_M1$$46894124_64x8m81_0_0
timestamp 1749760379
transform 1 0 140 0 1 5239
box 0 0 1 1
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_0
timestamp 1749760379
transform 0 1 310 -1 0 3199
box 0 0 1 1
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_1
timestamp 1749760379
transform 1 0 96 0 1 9568
box 0 0 1 1
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_2
timestamp 1749760379
transform 1 0 329 0 1 10756
box 0 0 1 1
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_3
timestamp 1749760379
transform 1 0 290 0 1 11535
box 0 0 1 1
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_4
timestamp 1749760379
transform 1 0 105 0 1 8520
box 0 0 1 1
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_5
timestamp 1749760379
transform 1 0 233 0 1 986
box 0 0 1 1
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_6
timestamp 1749760379
transform 1 0 327 0 1 7085
box 0 0 1 1
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_7
timestamp 1749760379
transform 1 0 520 0 1 9568
box 0 0 1 1
use M2_M14310589983228_64x8m81  M2_M14310589983228_64x8m81_0
timestamp 1749760379
transform 1 0 520 0 1 5035
box 0 0 1 1
use M3_M2$$43368492_64x8m81  M3_M2$$43368492_64x8m81_0
timestamp 1749760379
transform 1 0 140 0 1 5130
box 0 0 1 1
use nmos_5p0431058998320_64x8m81  nmos_5p0431058998320_64x8m81_0
timestamp 1749760379
transform 1 0 250 0 -1 6919
box 0 0 1 1
use nmos_5p0431058998320_64x8m81  nmos_5p0431058998320_64x8m81_1
timestamp 1749760379
transform 1 0 250 0 -1 4915
box 0 0 1 1
use nmos_5p0431058998322_64x8m81  nmos_5p0431058998322_64x8m81_0
timestamp 1749760379
transform 1 0 66 0 1 383
box 0 0 1 1
use pmos_5p0431058998321_64x8m81  pmos_5p0431058998321_64x8m81_0
timestamp 1749760379
transform 1 0 250 0 -1 3060
box 0 0 1 1
use pmos_5p0431058998321_64x8m81  pmos_5p0431058998321_64x8m81_1
timestamp 1749760379
transform 1 0 248 0 -1 10197
box 0 0 1 1
use pmos_5p0431058998321_64x8m81  pmos_5p0431058998321_64x8m81_2
timestamp 1749760379
transform 1 0 250 0 -1 8610
box 0 0 1 1
use via1_2_64x8m81_0  via1_2_64x8m81_0_0
timestamp 1749760379
transform 1 0 264 0 1 88
box 0 0 1 1
use via1_R90_64x8m81_0  via1_R90_64x8m81_0_0
timestamp 1749760379
transform 0 -1 378 1 0 3348
box 0 0 1 1
use via1_R90_64x8m81_0  via1_R90_64x8m81_0_1
timestamp 1749760379
transform 0 -1 373 1 0 12131
box 0 0 1 1
use via1_R90_64x8m81_0  via1_R90_64x8m81_0_2
timestamp 1749760379
transform 0 -1 373 1 0 11945
box 0 0 1 1
use via1_R270_64x8m81_0  via1_R270_64x8m81_0_0
timestamp 1749760379
transform 0 1 317 -1 0 1251
box 0 0 1 1
use via1_x2_R90_64x8m81_0  via1_x2_R90_64x8m81_0_0
timestamp 1749760379
transform 0 1 -154 1 0 5391
box 0 0 1 1
use via2_R90_64x8m81_0  via2_R90_64x8m81_0_0
timestamp 1749760379
transform 0 -1 373 1 0 11945
box 0 0 1 1
use via2_R90_64x8m81_0  via2_R90_64x8m81_0_1
timestamp 1749760379
transform 0 -1 373 1 0 12131
box 0 0 1 1
<< properties >>
string GDS_END 1041894
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1032530
string path 0.525 61.850 0.525 27.925 
<< end >>
