magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect 322 23861 5755 29123
rect 627 18373 5591 19955
rect 495 17401 5723 18373
rect 120 15330 750 15911
rect 1464 15330 2094 15663
rect 120 12907 2094 15330
rect 1449 9429 2303 9575
rect 1448 9398 2303 9429
rect 1448 9382 2930 9398
rect 621 9175 2930 9382
rect 100 8385 2930 9175
rect 620 8384 1475 8385
rect 2300 8384 2930 8385
rect 621 8303 1475 8384
rect 2301 7754 2930 8384
rect 3186 2694 3236 2701
<< mvnmos >>
rect 881 22310 1001 23672
rect 1501 22310 1621 23672
rect 2120 22310 2240 23672
rect 2740 22310 2860 23672
rect 3358 22310 3478 23672
rect 3978 22310 4098 23672
rect 4597 22310 4717 23672
rect 5217 22310 5337 23672
rect 881 20306 1001 21668
rect 1501 20306 1621 21668
rect 2120 20306 2240 21668
rect 2740 20306 2860 21668
rect 3358 20306 3478 21668
rect 3978 20306 4098 21668
rect 4597 20306 4717 21668
rect 5217 20306 5337 21668
rect 855 17136 975 17250
rect 1079 17136 1199 17250
rect 1303 17136 1423 17250
rect 1527 17136 1647 17250
rect 2094 17136 2214 17250
rect 2318 17136 2438 17250
rect 2542 17136 2662 17250
rect 2766 17136 2886 17250
rect 3332 17136 3452 17250
rect 3556 17136 3676 17250
rect 3780 17136 3900 17250
rect 4004 17136 4124 17250
rect 4571 17136 4691 17250
rect 4795 17136 4915 17250
rect 5019 17136 5139 17250
rect 5243 17136 5363 17250
rect 1043 15469 1163 15697
rect 375 9891 495 12613
rect 823 10344 943 12612
rect 1271 10344 1391 12612
rect 1719 10344 1839 12612
rect 986 9612 1106 9804
rect 1704 9712 1824 9904
rect 2556 9536 2676 9990
rect 876 7971 996 8163
rect 1100 7971 1220 8163
rect 1704 7950 1824 8142
rect 1928 7950 2048 8142
<< mvpmos >>
rect 769 27944 889 28626
rect 993 27944 1113 28626
rect 1389 27944 1509 28626
rect 1613 27944 1733 28626
rect 2008 27944 2128 28626
rect 2232 27944 2352 28626
rect 2628 27944 2748 28626
rect 2852 27944 2972 28626
rect 3246 27944 3366 28626
rect 3470 27944 3590 28626
rect 3866 27944 3986 28626
rect 4090 27944 4210 28626
rect 4485 27944 4605 28626
rect 4709 27944 4829 28626
rect 5069 27944 5189 28626
rect 5294 27944 5414 28626
rect 769 27169 889 27851
rect 993 27169 1113 27851
rect 1389 27169 1509 27851
rect 1613 27169 1733 27851
rect 2008 27169 2128 27851
rect 2232 27169 2352 27851
rect 2628 27169 2748 27851
rect 2852 27169 2972 27851
rect 3246 27169 3366 27851
rect 3470 27169 3590 27851
rect 3866 27169 3986 27851
rect 4090 27169 4210 27851
rect 4485 27169 4605 27851
rect 4709 27169 4829 27851
rect 5069 27169 5189 27851
rect 5294 27169 5414 27851
rect 883 25588 1003 26950
rect 1499 25588 1619 26950
rect 2122 25588 2242 26950
rect 2738 25588 2858 26950
rect 3360 25588 3480 26950
rect 3976 25588 4096 26950
rect 4599 25588 4719 26950
rect 5215 25588 5335 26950
rect 881 24001 1001 25363
rect 1501 24001 1621 25363
rect 2120 24001 2240 25363
rect 2740 24001 2860 25363
rect 3358 24001 3478 25363
rect 3978 24001 4098 25363
rect 4597 24001 4717 25363
rect 5217 24001 5337 25363
rect 881 18451 1001 19813
rect 1501 18451 1621 19813
rect 2120 18451 2240 19813
rect 2740 18451 2860 19813
rect 3358 18451 3478 19813
rect 3978 18451 4098 19813
rect 4597 18451 4717 19813
rect 5217 18451 5337 19813
rect 812 17541 932 17838
rect 1064 17541 1184 17838
rect 1318 17541 1438 17838
rect 1570 17541 1690 17838
rect 2051 17541 2171 17838
rect 2303 17541 2423 17838
rect 2557 17541 2677 17838
rect 2809 17541 2929 17838
rect 3289 17541 3409 17838
rect 3541 17541 3661 17838
rect 3795 17541 3915 17838
rect 4047 17541 4167 17838
rect 4528 17541 4648 17838
rect 4780 17541 4900 17838
rect 5034 17541 5154 17838
rect 5285 17541 5405 17838
rect 375 13049 495 15771
rect 928 14893 1048 15190
rect 1201 14893 1321 15190
rect 823 13049 943 14411
rect 1271 13049 1391 14411
rect 1719 13049 1839 15317
rect 876 9012 996 9240
rect 1100 9012 1220 9240
rect 1704 9205 1824 9433
rect 1928 9205 2048 9433
rect 876 8444 996 8636
rect 1100 8444 1220 8636
rect 1704 8526 1824 8718
rect 1928 8526 2048 8718
rect 2556 7896 2676 9258
<< mvndiff >>
rect 793 23659 881 23672
rect 793 23613 806 23659
rect 852 23613 881 23659
rect 793 23551 881 23613
rect 793 23505 806 23551
rect 852 23505 881 23551
rect 793 23443 881 23505
rect 793 23397 806 23443
rect 852 23397 881 23443
rect 793 23335 881 23397
rect 793 23289 806 23335
rect 852 23289 881 23335
rect 793 23227 881 23289
rect 793 23181 806 23227
rect 852 23181 881 23227
rect 793 23119 881 23181
rect 793 23073 806 23119
rect 852 23073 881 23119
rect 793 23011 881 23073
rect 793 22965 806 23011
rect 852 22965 881 23011
rect 793 22904 881 22965
rect 793 22858 806 22904
rect 852 22858 881 22904
rect 793 22797 881 22858
rect 793 22751 806 22797
rect 852 22751 881 22797
rect 793 22690 881 22751
rect 793 22644 806 22690
rect 852 22644 881 22690
rect 793 22583 881 22644
rect 793 22537 806 22583
rect 852 22537 881 22583
rect 793 22476 881 22537
rect 793 22430 806 22476
rect 852 22430 881 22476
rect 793 22369 881 22430
rect 793 22323 806 22369
rect 852 22323 881 22369
rect 793 22310 881 22323
rect 1001 23659 1089 23672
rect 1001 23613 1030 23659
rect 1076 23613 1089 23659
rect 1001 23551 1089 23613
rect 1001 23505 1030 23551
rect 1076 23505 1089 23551
rect 1001 23443 1089 23505
rect 1001 23397 1030 23443
rect 1076 23397 1089 23443
rect 1001 23335 1089 23397
rect 1001 23289 1030 23335
rect 1076 23289 1089 23335
rect 1001 23227 1089 23289
rect 1001 23181 1030 23227
rect 1076 23181 1089 23227
rect 1001 23119 1089 23181
rect 1001 23073 1030 23119
rect 1076 23073 1089 23119
rect 1001 23011 1089 23073
rect 1001 22965 1030 23011
rect 1076 22965 1089 23011
rect 1001 22904 1089 22965
rect 1001 22858 1030 22904
rect 1076 22858 1089 22904
rect 1001 22797 1089 22858
rect 1001 22751 1030 22797
rect 1076 22751 1089 22797
rect 1001 22690 1089 22751
rect 1001 22644 1030 22690
rect 1076 22644 1089 22690
rect 1001 22583 1089 22644
rect 1001 22537 1030 22583
rect 1076 22537 1089 22583
rect 1001 22476 1089 22537
rect 1001 22430 1030 22476
rect 1076 22430 1089 22476
rect 1001 22369 1089 22430
rect 1001 22323 1030 22369
rect 1076 22323 1089 22369
rect 1001 22310 1089 22323
rect 1413 23659 1501 23672
rect 1413 23613 1426 23659
rect 1472 23613 1501 23659
rect 1413 23551 1501 23613
rect 1413 23505 1426 23551
rect 1472 23505 1501 23551
rect 1413 23443 1501 23505
rect 1413 23397 1426 23443
rect 1472 23397 1501 23443
rect 1413 23335 1501 23397
rect 1413 23289 1426 23335
rect 1472 23289 1501 23335
rect 1413 23227 1501 23289
rect 1413 23181 1426 23227
rect 1472 23181 1501 23227
rect 1413 23119 1501 23181
rect 1413 23073 1426 23119
rect 1472 23073 1501 23119
rect 1413 23011 1501 23073
rect 1413 22965 1426 23011
rect 1472 22965 1501 23011
rect 1413 22904 1501 22965
rect 1413 22858 1426 22904
rect 1472 22858 1501 22904
rect 1413 22797 1501 22858
rect 1413 22751 1426 22797
rect 1472 22751 1501 22797
rect 1413 22690 1501 22751
rect 1413 22644 1426 22690
rect 1472 22644 1501 22690
rect 1413 22583 1501 22644
rect 1413 22537 1426 22583
rect 1472 22537 1501 22583
rect 1413 22476 1501 22537
rect 1413 22430 1426 22476
rect 1472 22430 1501 22476
rect 1413 22369 1501 22430
rect 1413 22323 1426 22369
rect 1472 22323 1501 22369
rect 1413 22310 1501 22323
rect 1621 23659 1709 23672
rect 1621 23613 1650 23659
rect 1696 23613 1709 23659
rect 1621 23551 1709 23613
rect 1621 23505 1650 23551
rect 1696 23505 1709 23551
rect 1621 23443 1709 23505
rect 1621 23397 1650 23443
rect 1696 23397 1709 23443
rect 1621 23335 1709 23397
rect 1621 23289 1650 23335
rect 1696 23289 1709 23335
rect 1621 23227 1709 23289
rect 1621 23181 1650 23227
rect 1696 23181 1709 23227
rect 1621 23119 1709 23181
rect 1621 23073 1650 23119
rect 1696 23073 1709 23119
rect 1621 23011 1709 23073
rect 1621 22965 1650 23011
rect 1696 22965 1709 23011
rect 1621 22904 1709 22965
rect 1621 22858 1650 22904
rect 1696 22858 1709 22904
rect 1621 22797 1709 22858
rect 1621 22751 1650 22797
rect 1696 22751 1709 22797
rect 1621 22690 1709 22751
rect 1621 22644 1650 22690
rect 1696 22644 1709 22690
rect 1621 22583 1709 22644
rect 1621 22537 1650 22583
rect 1696 22537 1709 22583
rect 1621 22476 1709 22537
rect 1621 22430 1650 22476
rect 1696 22430 1709 22476
rect 1621 22369 1709 22430
rect 1621 22323 1650 22369
rect 1696 22323 1709 22369
rect 1621 22310 1709 22323
rect 2032 23659 2120 23672
rect 2032 23613 2045 23659
rect 2091 23613 2120 23659
rect 2032 23551 2120 23613
rect 2032 23505 2045 23551
rect 2091 23505 2120 23551
rect 2032 23443 2120 23505
rect 2032 23397 2045 23443
rect 2091 23397 2120 23443
rect 2032 23335 2120 23397
rect 2032 23289 2045 23335
rect 2091 23289 2120 23335
rect 2032 23227 2120 23289
rect 2032 23181 2045 23227
rect 2091 23181 2120 23227
rect 2032 23119 2120 23181
rect 2032 23073 2045 23119
rect 2091 23073 2120 23119
rect 2032 23011 2120 23073
rect 2032 22965 2045 23011
rect 2091 22965 2120 23011
rect 2032 22904 2120 22965
rect 2032 22858 2045 22904
rect 2091 22858 2120 22904
rect 2032 22797 2120 22858
rect 2032 22751 2045 22797
rect 2091 22751 2120 22797
rect 2032 22690 2120 22751
rect 2032 22644 2045 22690
rect 2091 22644 2120 22690
rect 2032 22583 2120 22644
rect 2032 22537 2045 22583
rect 2091 22537 2120 22583
rect 2032 22476 2120 22537
rect 2032 22430 2045 22476
rect 2091 22430 2120 22476
rect 2032 22369 2120 22430
rect 2032 22323 2045 22369
rect 2091 22323 2120 22369
rect 2032 22310 2120 22323
rect 2240 23659 2328 23672
rect 2240 23613 2269 23659
rect 2315 23613 2328 23659
rect 2240 23551 2328 23613
rect 2240 23505 2269 23551
rect 2315 23505 2328 23551
rect 2240 23443 2328 23505
rect 2240 23397 2269 23443
rect 2315 23397 2328 23443
rect 2240 23335 2328 23397
rect 2240 23289 2269 23335
rect 2315 23289 2328 23335
rect 2240 23227 2328 23289
rect 2240 23181 2269 23227
rect 2315 23181 2328 23227
rect 2240 23119 2328 23181
rect 2240 23073 2269 23119
rect 2315 23073 2328 23119
rect 2240 23011 2328 23073
rect 2240 22965 2269 23011
rect 2315 22965 2328 23011
rect 2240 22904 2328 22965
rect 2240 22858 2269 22904
rect 2315 22858 2328 22904
rect 2240 22797 2328 22858
rect 2240 22751 2269 22797
rect 2315 22751 2328 22797
rect 2240 22690 2328 22751
rect 2240 22644 2269 22690
rect 2315 22644 2328 22690
rect 2240 22583 2328 22644
rect 2240 22537 2269 22583
rect 2315 22537 2328 22583
rect 2240 22476 2328 22537
rect 2240 22430 2269 22476
rect 2315 22430 2328 22476
rect 2240 22369 2328 22430
rect 2240 22323 2269 22369
rect 2315 22323 2328 22369
rect 2240 22310 2328 22323
rect 2652 23659 2740 23672
rect 2652 23613 2665 23659
rect 2711 23613 2740 23659
rect 2652 23551 2740 23613
rect 2652 23505 2665 23551
rect 2711 23505 2740 23551
rect 2652 23443 2740 23505
rect 2652 23397 2665 23443
rect 2711 23397 2740 23443
rect 2652 23335 2740 23397
rect 2652 23289 2665 23335
rect 2711 23289 2740 23335
rect 2652 23227 2740 23289
rect 2652 23181 2665 23227
rect 2711 23181 2740 23227
rect 2652 23119 2740 23181
rect 2652 23073 2665 23119
rect 2711 23073 2740 23119
rect 2652 23011 2740 23073
rect 2652 22965 2665 23011
rect 2711 22965 2740 23011
rect 2652 22904 2740 22965
rect 2652 22858 2665 22904
rect 2711 22858 2740 22904
rect 2652 22797 2740 22858
rect 2652 22751 2665 22797
rect 2711 22751 2740 22797
rect 2652 22690 2740 22751
rect 2652 22644 2665 22690
rect 2711 22644 2740 22690
rect 2652 22583 2740 22644
rect 2652 22537 2665 22583
rect 2711 22537 2740 22583
rect 2652 22476 2740 22537
rect 2652 22430 2665 22476
rect 2711 22430 2740 22476
rect 2652 22369 2740 22430
rect 2652 22323 2665 22369
rect 2711 22323 2740 22369
rect 2652 22310 2740 22323
rect 2860 23659 2948 23672
rect 2860 23613 2889 23659
rect 2935 23613 2948 23659
rect 2860 23551 2948 23613
rect 2860 23505 2889 23551
rect 2935 23505 2948 23551
rect 2860 23443 2948 23505
rect 2860 23397 2889 23443
rect 2935 23397 2948 23443
rect 2860 23335 2948 23397
rect 2860 23289 2889 23335
rect 2935 23289 2948 23335
rect 2860 23227 2948 23289
rect 2860 23181 2889 23227
rect 2935 23181 2948 23227
rect 2860 23119 2948 23181
rect 2860 23073 2889 23119
rect 2935 23073 2948 23119
rect 2860 23011 2948 23073
rect 2860 22965 2889 23011
rect 2935 22965 2948 23011
rect 2860 22904 2948 22965
rect 2860 22858 2889 22904
rect 2935 22858 2948 22904
rect 2860 22797 2948 22858
rect 2860 22751 2889 22797
rect 2935 22751 2948 22797
rect 2860 22690 2948 22751
rect 2860 22644 2889 22690
rect 2935 22644 2948 22690
rect 2860 22583 2948 22644
rect 2860 22537 2889 22583
rect 2935 22537 2948 22583
rect 2860 22476 2948 22537
rect 2860 22430 2889 22476
rect 2935 22430 2948 22476
rect 2860 22369 2948 22430
rect 2860 22323 2889 22369
rect 2935 22323 2948 22369
rect 2860 22310 2948 22323
rect 3270 23659 3358 23672
rect 3270 23613 3283 23659
rect 3329 23613 3358 23659
rect 3270 23551 3358 23613
rect 3270 23505 3283 23551
rect 3329 23505 3358 23551
rect 3270 23443 3358 23505
rect 3270 23397 3283 23443
rect 3329 23397 3358 23443
rect 3270 23335 3358 23397
rect 3270 23289 3283 23335
rect 3329 23289 3358 23335
rect 3270 23227 3358 23289
rect 3270 23181 3283 23227
rect 3329 23181 3358 23227
rect 3270 23119 3358 23181
rect 3270 23073 3283 23119
rect 3329 23073 3358 23119
rect 3270 23011 3358 23073
rect 3270 22965 3283 23011
rect 3329 22965 3358 23011
rect 3270 22904 3358 22965
rect 3270 22858 3283 22904
rect 3329 22858 3358 22904
rect 3270 22797 3358 22858
rect 3270 22751 3283 22797
rect 3329 22751 3358 22797
rect 3270 22690 3358 22751
rect 3270 22644 3283 22690
rect 3329 22644 3358 22690
rect 3270 22583 3358 22644
rect 3270 22537 3283 22583
rect 3329 22537 3358 22583
rect 3270 22476 3358 22537
rect 3270 22430 3283 22476
rect 3329 22430 3358 22476
rect 3270 22369 3358 22430
rect 3270 22323 3283 22369
rect 3329 22323 3358 22369
rect 3270 22310 3358 22323
rect 3478 23659 3566 23672
rect 3478 23613 3507 23659
rect 3553 23613 3566 23659
rect 3478 23551 3566 23613
rect 3478 23505 3507 23551
rect 3553 23505 3566 23551
rect 3478 23443 3566 23505
rect 3478 23397 3507 23443
rect 3553 23397 3566 23443
rect 3478 23335 3566 23397
rect 3478 23289 3507 23335
rect 3553 23289 3566 23335
rect 3478 23227 3566 23289
rect 3478 23181 3507 23227
rect 3553 23181 3566 23227
rect 3478 23119 3566 23181
rect 3478 23073 3507 23119
rect 3553 23073 3566 23119
rect 3478 23011 3566 23073
rect 3478 22965 3507 23011
rect 3553 22965 3566 23011
rect 3478 22904 3566 22965
rect 3478 22858 3507 22904
rect 3553 22858 3566 22904
rect 3478 22797 3566 22858
rect 3478 22751 3507 22797
rect 3553 22751 3566 22797
rect 3478 22690 3566 22751
rect 3478 22644 3507 22690
rect 3553 22644 3566 22690
rect 3478 22583 3566 22644
rect 3478 22537 3507 22583
rect 3553 22537 3566 22583
rect 3478 22476 3566 22537
rect 3478 22430 3507 22476
rect 3553 22430 3566 22476
rect 3478 22369 3566 22430
rect 3478 22323 3507 22369
rect 3553 22323 3566 22369
rect 3478 22310 3566 22323
rect 3890 23659 3978 23672
rect 3890 23613 3903 23659
rect 3949 23613 3978 23659
rect 3890 23551 3978 23613
rect 3890 23505 3903 23551
rect 3949 23505 3978 23551
rect 3890 23443 3978 23505
rect 3890 23397 3903 23443
rect 3949 23397 3978 23443
rect 3890 23335 3978 23397
rect 3890 23289 3903 23335
rect 3949 23289 3978 23335
rect 3890 23227 3978 23289
rect 3890 23181 3903 23227
rect 3949 23181 3978 23227
rect 3890 23119 3978 23181
rect 3890 23073 3903 23119
rect 3949 23073 3978 23119
rect 3890 23011 3978 23073
rect 3890 22965 3903 23011
rect 3949 22965 3978 23011
rect 3890 22904 3978 22965
rect 3890 22858 3903 22904
rect 3949 22858 3978 22904
rect 3890 22797 3978 22858
rect 3890 22751 3903 22797
rect 3949 22751 3978 22797
rect 3890 22690 3978 22751
rect 3890 22644 3903 22690
rect 3949 22644 3978 22690
rect 3890 22583 3978 22644
rect 3890 22537 3903 22583
rect 3949 22537 3978 22583
rect 3890 22476 3978 22537
rect 3890 22430 3903 22476
rect 3949 22430 3978 22476
rect 3890 22369 3978 22430
rect 3890 22323 3903 22369
rect 3949 22323 3978 22369
rect 3890 22310 3978 22323
rect 4098 23659 4186 23672
rect 4098 23613 4127 23659
rect 4173 23613 4186 23659
rect 4098 23551 4186 23613
rect 4098 23505 4127 23551
rect 4173 23505 4186 23551
rect 4098 23443 4186 23505
rect 4098 23397 4127 23443
rect 4173 23397 4186 23443
rect 4098 23335 4186 23397
rect 4098 23289 4127 23335
rect 4173 23289 4186 23335
rect 4098 23227 4186 23289
rect 4098 23181 4127 23227
rect 4173 23181 4186 23227
rect 4098 23119 4186 23181
rect 4098 23073 4127 23119
rect 4173 23073 4186 23119
rect 4098 23011 4186 23073
rect 4098 22965 4127 23011
rect 4173 22965 4186 23011
rect 4098 22904 4186 22965
rect 4098 22858 4127 22904
rect 4173 22858 4186 22904
rect 4098 22797 4186 22858
rect 4098 22751 4127 22797
rect 4173 22751 4186 22797
rect 4098 22690 4186 22751
rect 4098 22644 4127 22690
rect 4173 22644 4186 22690
rect 4098 22583 4186 22644
rect 4098 22537 4127 22583
rect 4173 22537 4186 22583
rect 4098 22476 4186 22537
rect 4098 22430 4127 22476
rect 4173 22430 4186 22476
rect 4098 22369 4186 22430
rect 4098 22323 4127 22369
rect 4173 22323 4186 22369
rect 4098 22310 4186 22323
rect 4509 23659 4597 23672
rect 4509 23613 4522 23659
rect 4568 23613 4597 23659
rect 4509 23551 4597 23613
rect 4509 23505 4522 23551
rect 4568 23505 4597 23551
rect 4509 23443 4597 23505
rect 4509 23397 4522 23443
rect 4568 23397 4597 23443
rect 4509 23335 4597 23397
rect 4509 23289 4522 23335
rect 4568 23289 4597 23335
rect 4509 23227 4597 23289
rect 4509 23181 4522 23227
rect 4568 23181 4597 23227
rect 4509 23119 4597 23181
rect 4509 23073 4522 23119
rect 4568 23073 4597 23119
rect 4509 23011 4597 23073
rect 4509 22965 4522 23011
rect 4568 22965 4597 23011
rect 4509 22904 4597 22965
rect 4509 22858 4522 22904
rect 4568 22858 4597 22904
rect 4509 22797 4597 22858
rect 4509 22751 4522 22797
rect 4568 22751 4597 22797
rect 4509 22690 4597 22751
rect 4509 22644 4522 22690
rect 4568 22644 4597 22690
rect 4509 22583 4597 22644
rect 4509 22537 4522 22583
rect 4568 22537 4597 22583
rect 4509 22476 4597 22537
rect 4509 22430 4522 22476
rect 4568 22430 4597 22476
rect 4509 22369 4597 22430
rect 4509 22323 4522 22369
rect 4568 22323 4597 22369
rect 4509 22310 4597 22323
rect 4717 23659 4805 23672
rect 4717 23613 4746 23659
rect 4792 23613 4805 23659
rect 4717 23551 4805 23613
rect 4717 23505 4746 23551
rect 4792 23505 4805 23551
rect 4717 23443 4805 23505
rect 4717 23397 4746 23443
rect 4792 23397 4805 23443
rect 4717 23335 4805 23397
rect 4717 23289 4746 23335
rect 4792 23289 4805 23335
rect 4717 23227 4805 23289
rect 4717 23181 4746 23227
rect 4792 23181 4805 23227
rect 4717 23119 4805 23181
rect 4717 23073 4746 23119
rect 4792 23073 4805 23119
rect 4717 23011 4805 23073
rect 4717 22965 4746 23011
rect 4792 22965 4805 23011
rect 4717 22904 4805 22965
rect 4717 22858 4746 22904
rect 4792 22858 4805 22904
rect 4717 22797 4805 22858
rect 4717 22751 4746 22797
rect 4792 22751 4805 22797
rect 4717 22690 4805 22751
rect 4717 22644 4746 22690
rect 4792 22644 4805 22690
rect 4717 22583 4805 22644
rect 4717 22537 4746 22583
rect 4792 22537 4805 22583
rect 4717 22476 4805 22537
rect 4717 22430 4746 22476
rect 4792 22430 4805 22476
rect 4717 22369 4805 22430
rect 4717 22323 4746 22369
rect 4792 22323 4805 22369
rect 4717 22310 4805 22323
rect 5129 23659 5217 23672
rect 5129 23613 5142 23659
rect 5188 23613 5217 23659
rect 5129 23551 5217 23613
rect 5129 23505 5142 23551
rect 5188 23505 5217 23551
rect 5129 23443 5217 23505
rect 5129 23397 5142 23443
rect 5188 23397 5217 23443
rect 5129 23335 5217 23397
rect 5129 23289 5142 23335
rect 5188 23289 5217 23335
rect 5129 23227 5217 23289
rect 5129 23181 5142 23227
rect 5188 23181 5217 23227
rect 5129 23119 5217 23181
rect 5129 23073 5142 23119
rect 5188 23073 5217 23119
rect 5129 23011 5217 23073
rect 5129 22965 5142 23011
rect 5188 22965 5217 23011
rect 5129 22904 5217 22965
rect 5129 22858 5142 22904
rect 5188 22858 5217 22904
rect 5129 22797 5217 22858
rect 5129 22751 5142 22797
rect 5188 22751 5217 22797
rect 5129 22690 5217 22751
rect 5129 22644 5142 22690
rect 5188 22644 5217 22690
rect 5129 22583 5217 22644
rect 5129 22537 5142 22583
rect 5188 22537 5217 22583
rect 5129 22476 5217 22537
rect 5129 22430 5142 22476
rect 5188 22430 5217 22476
rect 5129 22369 5217 22430
rect 5129 22323 5142 22369
rect 5188 22323 5217 22369
rect 5129 22310 5217 22323
rect 5337 23659 5425 23672
rect 5337 23613 5366 23659
rect 5412 23613 5425 23659
rect 5337 23551 5425 23613
rect 5337 23505 5366 23551
rect 5412 23505 5425 23551
rect 5337 23443 5425 23505
rect 5337 23397 5366 23443
rect 5412 23397 5425 23443
rect 5337 23335 5425 23397
rect 5337 23289 5366 23335
rect 5412 23289 5425 23335
rect 5337 23227 5425 23289
rect 5337 23181 5366 23227
rect 5412 23181 5425 23227
rect 5337 23119 5425 23181
rect 5337 23073 5366 23119
rect 5412 23073 5425 23119
rect 5337 23011 5425 23073
rect 5337 22965 5366 23011
rect 5412 22965 5425 23011
rect 5337 22904 5425 22965
rect 5337 22858 5366 22904
rect 5412 22858 5425 22904
rect 5337 22797 5425 22858
rect 5337 22751 5366 22797
rect 5412 22751 5425 22797
rect 5337 22690 5425 22751
rect 5337 22644 5366 22690
rect 5412 22644 5425 22690
rect 5337 22583 5425 22644
rect 5337 22537 5366 22583
rect 5412 22537 5425 22583
rect 5337 22476 5425 22537
rect 5337 22430 5366 22476
rect 5412 22430 5425 22476
rect 5337 22369 5425 22430
rect 5337 22323 5366 22369
rect 5412 22323 5425 22369
rect 5337 22310 5425 22323
rect 793 21655 881 21668
rect 793 21609 806 21655
rect 852 21609 881 21655
rect 793 21547 881 21609
rect 793 21501 806 21547
rect 852 21501 881 21547
rect 793 21439 881 21501
rect 793 21393 806 21439
rect 852 21393 881 21439
rect 793 21331 881 21393
rect 793 21285 806 21331
rect 852 21285 881 21331
rect 793 21223 881 21285
rect 793 21177 806 21223
rect 852 21177 881 21223
rect 793 21115 881 21177
rect 793 21069 806 21115
rect 852 21069 881 21115
rect 793 21007 881 21069
rect 793 20961 806 21007
rect 852 20961 881 21007
rect 793 20900 881 20961
rect 793 20854 806 20900
rect 852 20854 881 20900
rect 793 20793 881 20854
rect 793 20747 806 20793
rect 852 20747 881 20793
rect 793 20686 881 20747
rect 793 20640 806 20686
rect 852 20640 881 20686
rect 793 20579 881 20640
rect 793 20533 806 20579
rect 852 20533 881 20579
rect 793 20472 881 20533
rect 793 20426 806 20472
rect 852 20426 881 20472
rect 793 20365 881 20426
rect 793 20319 806 20365
rect 852 20319 881 20365
rect 793 20306 881 20319
rect 1001 21655 1089 21668
rect 1001 21609 1030 21655
rect 1076 21609 1089 21655
rect 1001 21547 1089 21609
rect 1001 21501 1030 21547
rect 1076 21501 1089 21547
rect 1001 21439 1089 21501
rect 1001 21393 1030 21439
rect 1076 21393 1089 21439
rect 1001 21331 1089 21393
rect 1001 21285 1030 21331
rect 1076 21285 1089 21331
rect 1001 21223 1089 21285
rect 1001 21177 1030 21223
rect 1076 21177 1089 21223
rect 1001 21115 1089 21177
rect 1001 21069 1030 21115
rect 1076 21069 1089 21115
rect 1001 21007 1089 21069
rect 1001 20961 1030 21007
rect 1076 20961 1089 21007
rect 1001 20900 1089 20961
rect 1001 20854 1030 20900
rect 1076 20854 1089 20900
rect 1001 20793 1089 20854
rect 1001 20747 1030 20793
rect 1076 20747 1089 20793
rect 1001 20686 1089 20747
rect 1001 20640 1030 20686
rect 1076 20640 1089 20686
rect 1001 20579 1089 20640
rect 1001 20533 1030 20579
rect 1076 20533 1089 20579
rect 1001 20472 1089 20533
rect 1001 20426 1030 20472
rect 1076 20426 1089 20472
rect 1001 20365 1089 20426
rect 1001 20319 1030 20365
rect 1076 20319 1089 20365
rect 1001 20306 1089 20319
rect 1413 21655 1501 21668
rect 1413 21609 1426 21655
rect 1472 21609 1501 21655
rect 1413 21547 1501 21609
rect 1413 21501 1426 21547
rect 1472 21501 1501 21547
rect 1413 21439 1501 21501
rect 1413 21393 1426 21439
rect 1472 21393 1501 21439
rect 1413 21331 1501 21393
rect 1413 21285 1426 21331
rect 1472 21285 1501 21331
rect 1413 21223 1501 21285
rect 1413 21177 1426 21223
rect 1472 21177 1501 21223
rect 1413 21115 1501 21177
rect 1413 21069 1426 21115
rect 1472 21069 1501 21115
rect 1413 21007 1501 21069
rect 1413 20961 1426 21007
rect 1472 20961 1501 21007
rect 1413 20900 1501 20961
rect 1413 20854 1426 20900
rect 1472 20854 1501 20900
rect 1413 20793 1501 20854
rect 1413 20747 1426 20793
rect 1472 20747 1501 20793
rect 1413 20686 1501 20747
rect 1413 20640 1426 20686
rect 1472 20640 1501 20686
rect 1413 20579 1501 20640
rect 1413 20533 1426 20579
rect 1472 20533 1501 20579
rect 1413 20472 1501 20533
rect 1413 20426 1426 20472
rect 1472 20426 1501 20472
rect 1413 20365 1501 20426
rect 1413 20319 1426 20365
rect 1472 20319 1501 20365
rect 1413 20306 1501 20319
rect 1621 21655 1709 21668
rect 1621 21609 1650 21655
rect 1696 21609 1709 21655
rect 1621 21547 1709 21609
rect 1621 21501 1650 21547
rect 1696 21501 1709 21547
rect 1621 21439 1709 21501
rect 1621 21393 1650 21439
rect 1696 21393 1709 21439
rect 1621 21331 1709 21393
rect 1621 21285 1650 21331
rect 1696 21285 1709 21331
rect 1621 21223 1709 21285
rect 1621 21177 1650 21223
rect 1696 21177 1709 21223
rect 1621 21115 1709 21177
rect 1621 21069 1650 21115
rect 1696 21069 1709 21115
rect 1621 21007 1709 21069
rect 1621 20961 1650 21007
rect 1696 20961 1709 21007
rect 1621 20900 1709 20961
rect 1621 20854 1650 20900
rect 1696 20854 1709 20900
rect 1621 20793 1709 20854
rect 1621 20747 1650 20793
rect 1696 20747 1709 20793
rect 1621 20686 1709 20747
rect 1621 20640 1650 20686
rect 1696 20640 1709 20686
rect 1621 20579 1709 20640
rect 1621 20533 1650 20579
rect 1696 20533 1709 20579
rect 1621 20472 1709 20533
rect 1621 20426 1650 20472
rect 1696 20426 1709 20472
rect 1621 20365 1709 20426
rect 1621 20319 1650 20365
rect 1696 20319 1709 20365
rect 1621 20306 1709 20319
rect 2032 21655 2120 21668
rect 2032 21609 2045 21655
rect 2091 21609 2120 21655
rect 2032 21547 2120 21609
rect 2032 21501 2045 21547
rect 2091 21501 2120 21547
rect 2032 21439 2120 21501
rect 2032 21393 2045 21439
rect 2091 21393 2120 21439
rect 2032 21331 2120 21393
rect 2032 21285 2045 21331
rect 2091 21285 2120 21331
rect 2032 21223 2120 21285
rect 2032 21177 2045 21223
rect 2091 21177 2120 21223
rect 2032 21115 2120 21177
rect 2032 21069 2045 21115
rect 2091 21069 2120 21115
rect 2032 21007 2120 21069
rect 2032 20961 2045 21007
rect 2091 20961 2120 21007
rect 2032 20900 2120 20961
rect 2032 20854 2045 20900
rect 2091 20854 2120 20900
rect 2032 20793 2120 20854
rect 2032 20747 2045 20793
rect 2091 20747 2120 20793
rect 2032 20686 2120 20747
rect 2032 20640 2045 20686
rect 2091 20640 2120 20686
rect 2032 20579 2120 20640
rect 2032 20533 2045 20579
rect 2091 20533 2120 20579
rect 2032 20472 2120 20533
rect 2032 20426 2045 20472
rect 2091 20426 2120 20472
rect 2032 20365 2120 20426
rect 2032 20319 2045 20365
rect 2091 20319 2120 20365
rect 2032 20306 2120 20319
rect 2240 21655 2328 21668
rect 2240 21609 2269 21655
rect 2315 21609 2328 21655
rect 2240 21547 2328 21609
rect 2240 21501 2269 21547
rect 2315 21501 2328 21547
rect 2240 21439 2328 21501
rect 2240 21393 2269 21439
rect 2315 21393 2328 21439
rect 2240 21331 2328 21393
rect 2240 21285 2269 21331
rect 2315 21285 2328 21331
rect 2240 21223 2328 21285
rect 2240 21177 2269 21223
rect 2315 21177 2328 21223
rect 2240 21115 2328 21177
rect 2240 21069 2269 21115
rect 2315 21069 2328 21115
rect 2240 21007 2328 21069
rect 2240 20961 2269 21007
rect 2315 20961 2328 21007
rect 2240 20900 2328 20961
rect 2240 20854 2269 20900
rect 2315 20854 2328 20900
rect 2240 20793 2328 20854
rect 2240 20747 2269 20793
rect 2315 20747 2328 20793
rect 2240 20686 2328 20747
rect 2240 20640 2269 20686
rect 2315 20640 2328 20686
rect 2240 20579 2328 20640
rect 2240 20533 2269 20579
rect 2315 20533 2328 20579
rect 2240 20472 2328 20533
rect 2240 20426 2269 20472
rect 2315 20426 2328 20472
rect 2240 20365 2328 20426
rect 2240 20319 2269 20365
rect 2315 20319 2328 20365
rect 2240 20306 2328 20319
rect 2652 21655 2740 21668
rect 2652 21609 2665 21655
rect 2711 21609 2740 21655
rect 2652 21547 2740 21609
rect 2652 21501 2665 21547
rect 2711 21501 2740 21547
rect 2652 21439 2740 21501
rect 2652 21393 2665 21439
rect 2711 21393 2740 21439
rect 2652 21331 2740 21393
rect 2652 21285 2665 21331
rect 2711 21285 2740 21331
rect 2652 21223 2740 21285
rect 2652 21177 2665 21223
rect 2711 21177 2740 21223
rect 2652 21115 2740 21177
rect 2652 21069 2665 21115
rect 2711 21069 2740 21115
rect 2652 21007 2740 21069
rect 2652 20961 2665 21007
rect 2711 20961 2740 21007
rect 2652 20900 2740 20961
rect 2652 20854 2665 20900
rect 2711 20854 2740 20900
rect 2652 20793 2740 20854
rect 2652 20747 2665 20793
rect 2711 20747 2740 20793
rect 2652 20686 2740 20747
rect 2652 20640 2665 20686
rect 2711 20640 2740 20686
rect 2652 20579 2740 20640
rect 2652 20533 2665 20579
rect 2711 20533 2740 20579
rect 2652 20472 2740 20533
rect 2652 20426 2665 20472
rect 2711 20426 2740 20472
rect 2652 20365 2740 20426
rect 2652 20319 2665 20365
rect 2711 20319 2740 20365
rect 2652 20306 2740 20319
rect 2860 21655 2948 21668
rect 2860 21609 2889 21655
rect 2935 21609 2948 21655
rect 2860 21547 2948 21609
rect 2860 21501 2889 21547
rect 2935 21501 2948 21547
rect 2860 21439 2948 21501
rect 2860 21393 2889 21439
rect 2935 21393 2948 21439
rect 2860 21331 2948 21393
rect 2860 21285 2889 21331
rect 2935 21285 2948 21331
rect 2860 21223 2948 21285
rect 2860 21177 2889 21223
rect 2935 21177 2948 21223
rect 2860 21115 2948 21177
rect 2860 21069 2889 21115
rect 2935 21069 2948 21115
rect 2860 21007 2948 21069
rect 2860 20961 2889 21007
rect 2935 20961 2948 21007
rect 2860 20900 2948 20961
rect 2860 20854 2889 20900
rect 2935 20854 2948 20900
rect 2860 20793 2948 20854
rect 2860 20747 2889 20793
rect 2935 20747 2948 20793
rect 2860 20686 2948 20747
rect 2860 20640 2889 20686
rect 2935 20640 2948 20686
rect 2860 20579 2948 20640
rect 2860 20533 2889 20579
rect 2935 20533 2948 20579
rect 2860 20472 2948 20533
rect 2860 20426 2889 20472
rect 2935 20426 2948 20472
rect 2860 20365 2948 20426
rect 2860 20319 2889 20365
rect 2935 20319 2948 20365
rect 2860 20306 2948 20319
rect 3270 21655 3358 21668
rect 3270 21609 3283 21655
rect 3329 21609 3358 21655
rect 3270 21547 3358 21609
rect 3270 21501 3283 21547
rect 3329 21501 3358 21547
rect 3270 21439 3358 21501
rect 3270 21393 3283 21439
rect 3329 21393 3358 21439
rect 3270 21331 3358 21393
rect 3270 21285 3283 21331
rect 3329 21285 3358 21331
rect 3270 21223 3358 21285
rect 3270 21177 3283 21223
rect 3329 21177 3358 21223
rect 3270 21115 3358 21177
rect 3270 21069 3283 21115
rect 3329 21069 3358 21115
rect 3270 21007 3358 21069
rect 3270 20961 3283 21007
rect 3329 20961 3358 21007
rect 3270 20900 3358 20961
rect 3270 20854 3283 20900
rect 3329 20854 3358 20900
rect 3270 20793 3358 20854
rect 3270 20747 3283 20793
rect 3329 20747 3358 20793
rect 3270 20686 3358 20747
rect 3270 20640 3283 20686
rect 3329 20640 3358 20686
rect 3270 20579 3358 20640
rect 3270 20533 3283 20579
rect 3329 20533 3358 20579
rect 3270 20472 3358 20533
rect 3270 20426 3283 20472
rect 3329 20426 3358 20472
rect 3270 20365 3358 20426
rect 3270 20319 3283 20365
rect 3329 20319 3358 20365
rect 3270 20306 3358 20319
rect 3478 21655 3566 21668
rect 3478 21609 3507 21655
rect 3553 21609 3566 21655
rect 3478 21547 3566 21609
rect 3478 21501 3507 21547
rect 3553 21501 3566 21547
rect 3478 21439 3566 21501
rect 3478 21393 3507 21439
rect 3553 21393 3566 21439
rect 3478 21331 3566 21393
rect 3478 21285 3507 21331
rect 3553 21285 3566 21331
rect 3478 21223 3566 21285
rect 3478 21177 3507 21223
rect 3553 21177 3566 21223
rect 3478 21115 3566 21177
rect 3478 21069 3507 21115
rect 3553 21069 3566 21115
rect 3478 21007 3566 21069
rect 3478 20961 3507 21007
rect 3553 20961 3566 21007
rect 3478 20900 3566 20961
rect 3478 20854 3507 20900
rect 3553 20854 3566 20900
rect 3478 20793 3566 20854
rect 3478 20747 3507 20793
rect 3553 20747 3566 20793
rect 3478 20686 3566 20747
rect 3478 20640 3507 20686
rect 3553 20640 3566 20686
rect 3478 20579 3566 20640
rect 3478 20533 3507 20579
rect 3553 20533 3566 20579
rect 3478 20472 3566 20533
rect 3478 20426 3507 20472
rect 3553 20426 3566 20472
rect 3478 20365 3566 20426
rect 3478 20319 3507 20365
rect 3553 20319 3566 20365
rect 3478 20306 3566 20319
rect 3890 21655 3978 21668
rect 3890 21609 3903 21655
rect 3949 21609 3978 21655
rect 3890 21547 3978 21609
rect 3890 21501 3903 21547
rect 3949 21501 3978 21547
rect 3890 21439 3978 21501
rect 3890 21393 3903 21439
rect 3949 21393 3978 21439
rect 3890 21331 3978 21393
rect 3890 21285 3903 21331
rect 3949 21285 3978 21331
rect 3890 21223 3978 21285
rect 3890 21177 3903 21223
rect 3949 21177 3978 21223
rect 3890 21115 3978 21177
rect 3890 21069 3903 21115
rect 3949 21069 3978 21115
rect 3890 21007 3978 21069
rect 3890 20961 3903 21007
rect 3949 20961 3978 21007
rect 3890 20900 3978 20961
rect 3890 20854 3903 20900
rect 3949 20854 3978 20900
rect 3890 20793 3978 20854
rect 3890 20747 3903 20793
rect 3949 20747 3978 20793
rect 3890 20686 3978 20747
rect 3890 20640 3903 20686
rect 3949 20640 3978 20686
rect 3890 20579 3978 20640
rect 3890 20533 3903 20579
rect 3949 20533 3978 20579
rect 3890 20472 3978 20533
rect 3890 20426 3903 20472
rect 3949 20426 3978 20472
rect 3890 20365 3978 20426
rect 3890 20319 3903 20365
rect 3949 20319 3978 20365
rect 3890 20306 3978 20319
rect 4098 21655 4186 21668
rect 4098 21609 4127 21655
rect 4173 21609 4186 21655
rect 4098 21547 4186 21609
rect 4098 21501 4127 21547
rect 4173 21501 4186 21547
rect 4098 21439 4186 21501
rect 4098 21393 4127 21439
rect 4173 21393 4186 21439
rect 4098 21331 4186 21393
rect 4098 21285 4127 21331
rect 4173 21285 4186 21331
rect 4098 21223 4186 21285
rect 4098 21177 4127 21223
rect 4173 21177 4186 21223
rect 4098 21115 4186 21177
rect 4098 21069 4127 21115
rect 4173 21069 4186 21115
rect 4098 21007 4186 21069
rect 4098 20961 4127 21007
rect 4173 20961 4186 21007
rect 4098 20900 4186 20961
rect 4098 20854 4127 20900
rect 4173 20854 4186 20900
rect 4098 20793 4186 20854
rect 4098 20747 4127 20793
rect 4173 20747 4186 20793
rect 4098 20686 4186 20747
rect 4098 20640 4127 20686
rect 4173 20640 4186 20686
rect 4098 20579 4186 20640
rect 4098 20533 4127 20579
rect 4173 20533 4186 20579
rect 4098 20472 4186 20533
rect 4098 20426 4127 20472
rect 4173 20426 4186 20472
rect 4098 20365 4186 20426
rect 4098 20319 4127 20365
rect 4173 20319 4186 20365
rect 4098 20306 4186 20319
rect 4509 21655 4597 21668
rect 4509 21609 4522 21655
rect 4568 21609 4597 21655
rect 4509 21547 4597 21609
rect 4509 21501 4522 21547
rect 4568 21501 4597 21547
rect 4509 21439 4597 21501
rect 4509 21393 4522 21439
rect 4568 21393 4597 21439
rect 4509 21331 4597 21393
rect 4509 21285 4522 21331
rect 4568 21285 4597 21331
rect 4509 21223 4597 21285
rect 4509 21177 4522 21223
rect 4568 21177 4597 21223
rect 4509 21115 4597 21177
rect 4509 21069 4522 21115
rect 4568 21069 4597 21115
rect 4509 21007 4597 21069
rect 4509 20961 4522 21007
rect 4568 20961 4597 21007
rect 4509 20900 4597 20961
rect 4509 20854 4522 20900
rect 4568 20854 4597 20900
rect 4509 20793 4597 20854
rect 4509 20747 4522 20793
rect 4568 20747 4597 20793
rect 4509 20686 4597 20747
rect 4509 20640 4522 20686
rect 4568 20640 4597 20686
rect 4509 20579 4597 20640
rect 4509 20533 4522 20579
rect 4568 20533 4597 20579
rect 4509 20472 4597 20533
rect 4509 20426 4522 20472
rect 4568 20426 4597 20472
rect 4509 20365 4597 20426
rect 4509 20319 4522 20365
rect 4568 20319 4597 20365
rect 4509 20306 4597 20319
rect 4717 21655 4805 21668
rect 4717 21609 4746 21655
rect 4792 21609 4805 21655
rect 4717 21547 4805 21609
rect 4717 21501 4746 21547
rect 4792 21501 4805 21547
rect 4717 21439 4805 21501
rect 4717 21393 4746 21439
rect 4792 21393 4805 21439
rect 4717 21331 4805 21393
rect 4717 21285 4746 21331
rect 4792 21285 4805 21331
rect 4717 21223 4805 21285
rect 4717 21177 4746 21223
rect 4792 21177 4805 21223
rect 4717 21115 4805 21177
rect 4717 21069 4746 21115
rect 4792 21069 4805 21115
rect 4717 21007 4805 21069
rect 4717 20961 4746 21007
rect 4792 20961 4805 21007
rect 4717 20900 4805 20961
rect 4717 20854 4746 20900
rect 4792 20854 4805 20900
rect 4717 20793 4805 20854
rect 4717 20747 4746 20793
rect 4792 20747 4805 20793
rect 4717 20686 4805 20747
rect 4717 20640 4746 20686
rect 4792 20640 4805 20686
rect 4717 20579 4805 20640
rect 4717 20533 4746 20579
rect 4792 20533 4805 20579
rect 4717 20472 4805 20533
rect 4717 20426 4746 20472
rect 4792 20426 4805 20472
rect 4717 20365 4805 20426
rect 4717 20319 4746 20365
rect 4792 20319 4805 20365
rect 4717 20306 4805 20319
rect 5129 21655 5217 21668
rect 5129 21609 5142 21655
rect 5188 21609 5217 21655
rect 5129 21547 5217 21609
rect 5129 21501 5142 21547
rect 5188 21501 5217 21547
rect 5129 21439 5217 21501
rect 5129 21393 5142 21439
rect 5188 21393 5217 21439
rect 5129 21331 5217 21393
rect 5129 21285 5142 21331
rect 5188 21285 5217 21331
rect 5129 21223 5217 21285
rect 5129 21177 5142 21223
rect 5188 21177 5217 21223
rect 5129 21115 5217 21177
rect 5129 21069 5142 21115
rect 5188 21069 5217 21115
rect 5129 21007 5217 21069
rect 5129 20961 5142 21007
rect 5188 20961 5217 21007
rect 5129 20900 5217 20961
rect 5129 20854 5142 20900
rect 5188 20854 5217 20900
rect 5129 20793 5217 20854
rect 5129 20747 5142 20793
rect 5188 20747 5217 20793
rect 5129 20686 5217 20747
rect 5129 20640 5142 20686
rect 5188 20640 5217 20686
rect 5129 20579 5217 20640
rect 5129 20533 5142 20579
rect 5188 20533 5217 20579
rect 5129 20472 5217 20533
rect 5129 20426 5142 20472
rect 5188 20426 5217 20472
rect 5129 20365 5217 20426
rect 5129 20319 5142 20365
rect 5188 20319 5217 20365
rect 5129 20306 5217 20319
rect 5337 21655 5425 21668
rect 5337 21609 5366 21655
rect 5412 21609 5425 21655
rect 5337 21547 5425 21609
rect 5337 21501 5366 21547
rect 5412 21501 5425 21547
rect 5337 21439 5425 21501
rect 5337 21393 5366 21439
rect 5412 21393 5425 21439
rect 5337 21331 5425 21393
rect 5337 21285 5366 21331
rect 5412 21285 5425 21331
rect 5337 21223 5425 21285
rect 5337 21177 5366 21223
rect 5412 21177 5425 21223
rect 5337 21115 5425 21177
rect 5337 21069 5366 21115
rect 5412 21069 5425 21115
rect 5337 21007 5425 21069
rect 5337 20961 5366 21007
rect 5412 20961 5425 21007
rect 5337 20900 5425 20961
rect 5337 20854 5366 20900
rect 5412 20854 5425 20900
rect 5337 20793 5425 20854
rect 5337 20747 5366 20793
rect 5412 20747 5425 20793
rect 5337 20686 5425 20747
rect 5337 20640 5366 20686
rect 5412 20640 5425 20686
rect 5337 20579 5425 20640
rect 5337 20533 5366 20579
rect 5412 20533 5425 20579
rect 5337 20472 5425 20533
rect 5337 20426 5366 20472
rect 5412 20426 5425 20472
rect 5337 20365 5425 20426
rect 5337 20319 5366 20365
rect 5412 20319 5425 20365
rect 5337 20306 5425 20319
rect 767 17216 855 17250
rect 767 17170 780 17216
rect 826 17170 855 17216
rect 767 17136 855 17170
rect 975 17216 1079 17250
rect 975 17170 1004 17216
rect 1050 17170 1079 17216
rect 975 17136 1079 17170
rect 1199 17216 1303 17250
rect 1199 17170 1228 17216
rect 1274 17170 1303 17216
rect 1199 17136 1303 17170
rect 1423 17216 1527 17250
rect 1423 17170 1452 17216
rect 1498 17170 1527 17216
rect 1423 17136 1527 17170
rect 1647 17216 1735 17250
rect 1647 17170 1676 17216
rect 1722 17170 1735 17216
rect 1647 17136 1735 17170
rect 2006 17216 2094 17250
rect 2006 17170 2019 17216
rect 2065 17170 2094 17216
rect 2006 17136 2094 17170
rect 2214 17216 2318 17250
rect 2214 17170 2243 17216
rect 2289 17170 2318 17216
rect 2214 17136 2318 17170
rect 2438 17216 2542 17250
rect 2438 17170 2467 17216
rect 2513 17170 2542 17216
rect 2438 17136 2542 17170
rect 2662 17216 2766 17250
rect 2662 17170 2691 17216
rect 2737 17170 2766 17216
rect 2662 17136 2766 17170
rect 2886 17216 2974 17250
rect 2886 17170 2915 17216
rect 2961 17170 2974 17216
rect 2886 17136 2974 17170
rect 3244 17216 3332 17250
rect 3244 17170 3257 17216
rect 3303 17170 3332 17216
rect 3244 17136 3332 17170
rect 3452 17216 3556 17250
rect 3452 17170 3481 17216
rect 3527 17170 3556 17216
rect 3452 17136 3556 17170
rect 3676 17216 3780 17250
rect 3676 17170 3705 17216
rect 3751 17170 3780 17216
rect 3676 17136 3780 17170
rect 3900 17216 4004 17250
rect 3900 17170 3929 17216
rect 3975 17170 4004 17216
rect 3900 17136 4004 17170
rect 4124 17216 4212 17250
rect 4124 17170 4153 17216
rect 4199 17170 4212 17216
rect 4124 17136 4212 17170
rect 4483 17216 4571 17250
rect 4483 17170 4496 17216
rect 4542 17170 4571 17216
rect 4483 17136 4571 17170
rect 4691 17216 4795 17250
rect 4691 17170 4720 17216
rect 4766 17170 4795 17216
rect 4691 17136 4795 17170
rect 4915 17216 5019 17250
rect 4915 17170 4944 17216
rect 4990 17170 5019 17216
rect 4915 17136 5019 17170
rect 5139 17216 5243 17250
rect 5139 17170 5168 17216
rect 5214 17170 5243 17216
rect 5139 17136 5243 17170
rect 5363 17216 5451 17250
rect 5363 17170 5392 17216
rect 5438 17170 5451 17216
rect 5363 17136 5451 17170
rect 904 15584 1043 15697
rect 904 15538 948 15584
rect 994 15538 1043 15584
rect 904 15469 1043 15538
rect 1163 15584 1301 15697
rect 1163 15538 1211 15584
rect 1257 15538 1301 15584
rect 1163 15469 1301 15538
rect 287 12600 375 12613
rect 287 9904 300 12600
rect 346 9904 375 12600
rect 287 9891 375 9904
rect 495 12600 583 12613
rect 495 9904 524 12600
rect 570 9904 583 12600
rect 735 12599 823 12612
rect 735 12553 748 12599
rect 794 12553 823 12599
rect 735 12495 823 12553
rect 735 12449 748 12495
rect 794 12449 823 12495
rect 735 12391 823 12449
rect 735 12345 748 12391
rect 794 12345 823 12391
rect 735 12287 823 12345
rect 735 12241 748 12287
rect 794 12241 823 12287
rect 735 12183 823 12241
rect 735 12137 748 12183
rect 794 12137 823 12183
rect 735 12079 823 12137
rect 735 12033 748 12079
rect 794 12033 823 12079
rect 735 11975 823 12033
rect 735 11929 748 11975
rect 794 11929 823 11975
rect 735 11871 823 11929
rect 735 11825 748 11871
rect 794 11825 823 11871
rect 735 11767 823 11825
rect 735 11721 748 11767
rect 794 11721 823 11767
rect 735 11663 823 11721
rect 735 11617 748 11663
rect 794 11617 823 11663
rect 735 11558 823 11617
rect 735 11512 748 11558
rect 794 11512 823 11558
rect 735 11453 823 11512
rect 735 11407 748 11453
rect 794 11407 823 11453
rect 735 11348 823 11407
rect 735 11302 748 11348
rect 794 11302 823 11348
rect 735 11243 823 11302
rect 735 11197 748 11243
rect 794 11197 823 11243
rect 735 11138 823 11197
rect 735 11092 748 11138
rect 794 11092 823 11138
rect 735 11033 823 11092
rect 735 10987 748 11033
rect 794 10987 823 11033
rect 735 10928 823 10987
rect 735 10882 748 10928
rect 794 10882 823 10928
rect 735 10823 823 10882
rect 735 10777 748 10823
rect 794 10777 823 10823
rect 735 10718 823 10777
rect 735 10672 748 10718
rect 794 10672 823 10718
rect 735 10613 823 10672
rect 735 10567 748 10613
rect 794 10567 823 10613
rect 735 10508 823 10567
rect 735 10462 748 10508
rect 794 10462 823 10508
rect 735 10403 823 10462
rect 735 10357 748 10403
rect 794 10357 823 10403
rect 735 10344 823 10357
rect 943 12599 1031 12612
rect 943 12553 972 12599
rect 1018 12553 1031 12599
rect 943 12495 1031 12553
rect 943 12449 972 12495
rect 1018 12449 1031 12495
rect 943 12391 1031 12449
rect 943 12345 972 12391
rect 1018 12345 1031 12391
rect 943 12287 1031 12345
rect 943 12241 972 12287
rect 1018 12241 1031 12287
rect 943 12183 1031 12241
rect 943 12137 972 12183
rect 1018 12137 1031 12183
rect 943 12079 1031 12137
rect 943 12033 972 12079
rect 1018 12033 1031 12079
rect 943 11975 1031 12033
rect 943 11929 972 11975
rect 1018 11929 1031 11975
rect 943 11871 1031 11929
rect 943 11825 972 11871
rect 1018 11825 1031 11871
rect 943 11767 1031 11825
rect 943 11721 972 11767
rect 1018 11721 1031 11767
rect 943 11663 1031 11721
rect 943 11617 972 11663
rect 1018 11617 1031 11663
rect 943 11558 1031 11617
rect 943 11512 972 11558
rect 1018 11512 1031 11558
rect 943 11453 1031 11512
rect 943 11407 972 11453
rect 1018 11407 1031 11453
rect 943 11348 1031 11407
rect 943 11302 972 11348
rect 1018 11302 1031 11348
rect 943 11243 1031 11302
rect 943 11197 972 11243
rect 1018 11197 1031 11243
rect 943 11138 1031 11197
rect 943 11092 972 11138
rect 1018 11092 1031 11138
rect 943 11033 1031 11092
rect 943 10987 972 11033
rect 1018 10987 1031 11033
rect 943 10928 1031 10987
rect 943 10882 972 10928
rect 1018 10882 1031 10928
rect 943 10823 1031 10882
rect 943 10777 972 10823
rect 1018 10777 1031 10823
rect 943 10718 1031 10777
rect 943 10672 972 10718
rect 1018 10672 1031 10718
rect 943 10613 1031 10672
rect 943 10567 972 10613
rect 1018 10567 1031 10613
rect 943 10508 1031 10567
rect 943 10462 972 10508
rect 1018 10462 1031 10508
rect 943 10403 1031 10462
rect 943 10357 972 10403
rect 1018 10357 1031 10403
rect 943 10344 1031 10357
rect 1183 12599 1271 12612
rect 1183 12553 1196 12599
rect 1242 12553 1271 12599
rect 1183 12495 1271 12553
rect 1183 12449 1196 12495
rect 1242 12449 1271 12495
rect 1183 12391 1271 12449
rect 1183 12345 1196 12391
rect 1242 12345 1271 12391
rect 1183 12287 1271 12345
rect 1183 12241 1196 12287
rect 1242 12241 1271 12287
rect 1183 12183 1271 12241
rect 1183 12137 1196 12183
rect 1242 12137 1271 12183
rect 1183 12079 1271 12137
rect 1183 12033 1196 12079
rect 1242 12033 1271 12079
rect 1183 11975 1271 12033
rect 1183 11929 1196 11975
rect 1242 11929 1271 11975
rect 1183 11871 1271 11929
rect 1183 11825 1196 11871
rect 1242 11825 1271 11871
rect 1183 11767 1271 11825
rect 1183 11721 1196 11767
rect 1242 11721 1271 11767
rect 1183 11663 1271 11721
rect 1183 11617 1196 11663
rect 1242 11617 1271 11663
rect 1183 11558 1271 11617
rect 1183 11512 1196 11558
rect 1242 11512 1271 11558
rect 1183 11453 1271 11512
rect 1183 11407 1196 11453
rect 1242 11407 1271 11453
rect 1183 11348 1271 11407
rect 1183 11302 1196 11348
rect 1242 11302 1271 11348
rect 1183 11243 1271 11302
rect 1183 11197 1196 11243
rect 1242 11197 1271 11243
rect 1183 11138 1271 11197
rect 1183 11092 1196 11138
rect 1242 11092 1271 11138
rect 1183 11033 1271 11092
rect 1183 10987 1196 11033
rect 1242 10987 1271 11033
rect 1183 10928 1271 10987
rect 1183 10882 1196 10928
rect 1242 10882 1271 10928
rect 1183 10823 1271 10882
rect 1183 10777 1196 10823
rect 1242 10777 1271 10823
rect 1183 10718 1271 10777
rect 1183 10672 1196 10718
rect 1242 10672 1271 10718
rect 1183 10613 1271 10672
rect 1183 10567 1196 10613
rect 1242 10567 1271 10613
rect 1183 10508 1271 10567
rect 1183 10462 1196 10508
rect 1242 10462 1271 10508
rect 1183 10403 1271 10462
rect 1183 10357 1196 10403
rect 1242 10357 1271 10403
rect 1183 10344 1271 10357
rect 1391 12599 1479 12612
rect 1391 12553 1420 12599
rect 1466 12553 1479 12599
rect 1391 12495 1479 12553
rect 1391 12449 1420 12495
rect 1466 12449 1479 12495
rect 1391 12391 1479 12449
rect 1391 12345 1420 12391
rect 1466 12345 1479 12391
rect 1391 12287 1479 12345
rect 1391 12241 1420 12287
rect 1466 12241 1479 12287
rect 1391 12183 1479 12241
rect 1391 12137 1420 12183
rect 1466 12137 1479 12183
rect 1391 12079 1479 12137
rect 1391 12033 1420 12079
rect 1466 12033 1479 12079
rect 1391 11975 1479 12033
rect 1391 11929 1420 11975
rect 1466 11929 1479 11975
rect 1391 11871 1479 11929
rect 1391 11825 1420 11871
rect 1466 11825 1479 11871
rect 1391 11767 1479 11825
rect 1391 11721 1420 11767
rect 1466 11721 1479 11767
rect 1391 11663 1479 11721
rect 1391 11617 1420 11663
rect 1466 11617 1479 11663
rect 1391 11558 1479 11617
rect 1391 11512 1420 11558
rect 1466 11512 1479 11558
rect 1391 11453 1479 11512
rect 1391 11407 1420 11453
rect 1466 11407 1479 11453
rect 1391 11348 1479 11407
rect 1391 11302 1420 11348
rect 1466 11302 1479 11348
rect 1391 11243 1479 11302
rect 1391 11197 1420 11243
rect 1466 11197 1479 11243
rect 1391 11138 1479 11197
rect 1391 11092 1420 11138
rect 1466 11092 1479 11138
rect 1391 11033 1479 11092
rect 1391 10987 1420 11033
rect 1466 10987 1479 11033
rect 1391 10928 1479 10987
rect 1391 10882 1420 10928
rect 1466 10882 1479 10928
rect 1391 10823 1479 10882
rect 1391 10777 1420 10823
rect 1466 10777 1479 10823
rect 1391 10718 1479 10777
rect 1391 10672 1420 10718
rect 1466 10672 1479 10718
rect 1391 10613 1479 10672
rect 1391 10567 1420 10613
rect 1466 10567 1479 10613
rect 1391 10508 1479 10567
rect 1391 10462 1420 10508
rect 1466 10462 1479 10508
rect 1391 10403 1479 10462
rect 1391 10357 1420 10403
rect 1466 10357 1479 10403
rect 1391 10344 1479 10357
rect 1631 12599 1719 12612
rect 1631 12553 1644 12599
rect 1690 12553 1719 12599
rect 1631 12495 1719 12553
rect 1631 12449 1644 12495
rect 1690 12449 1719 12495
rect 1631 12391 1719 12449
rect 1631 12345 1644 12391
rect 1690 12345 1719 12391
rect 1631 12287 1719 12345
rect 1631 12241 1644 12287
rect 1690 12241 1719 12287
rect 1631 12183 1719 12241
rect 1631 12137 1644 12183
rect 1690 12137 1719 12183
rect 1631 12079 1719 12137
rect 1631 12033 1644 12079
rect 1690 12033 1719 12079
rect 1631 11975 1719 12033
rect 1631 11929 1644 11975
rect 1690 11929 1719 11975
rect 1631 11871 1719 11929
rect 1631 11825 1644 11871
rect 1690 11825 1719 11871
rect 1631 11767 1719 11825
rect 1631 11721 1644 11767
rect 1690 11721 1719 11767
rect 1631 11663 1719 11721
rect 1631 11617 1644 11663
rect 1690 11617 1719 11663
rect 1631 11558 1719 11617
rect 1631 11512 1644 11558
rect 1690 11512 1719 11558
rect 1631 11453 1719 11512
rect 1631 11407 1644 11453
rect 1690 11407 1719 11453
rect 1631 11348 1719 11407
rect 1631 11302 1644 11348
rect 1690 11302 1719 11348
rect 1631 11243 1719 11302
rect 1631 11197 1644 11243
rect 1690 11197 1719 11243
rect 1631 11138 1719 11197
rect 1631 11092 1644 11138
rect 1690 11092 1719 11138
rect 1631 11033 1719 11092
rect 1631 10987 1644 11033
rect 1690 10987 1719 11033
rect 1631 10928 1719 10987
rect 1631 10882 1644 10928
rect 1690 10882 1719 10928
rect 1631 10823 1719 10882
rect 1631 10777 1644 10823
rect 1690 10777 1719 10823
rect 1631 10718 1719 10777
rect 1631 10672 1644 10718
rect 1690 10672 1719 10718
rect 1631 10613 1719 10672
rect 1631 10567 1644 10613
rect 1690 10567 1719 10613
rect 1631 10508 1719 10567
rect 1631 10462 1644 10508
rect 1690 10462 1719 10508
rect 1631 10403 1719 10462
rect 1631 10357 1644 10403
rect 1690 10357 1719 10403
rect 1631 10344 1719 10357
rect 1839 12599 1927 12612
rect 1839 12553 1868 12599
rect 1914 12553 1927 12599
rect 1839 12495 1927 12553
rect 1839 12449 1868 12495
rect 1914 12449 1927 12495
rect 1839 12391 1927 12449
rect 1839 12345 1868 12391
rect 1914 12345 1927 12391
rect 1839 12287 1927 12345
rect 1839 12241 1868 12287
rect 1914 12241 1927 12287
rect 1839 12183 1927 12241
rect 1839 12137 1868 12183
rect 1914 12137 1927 12183
rect 1839 12079 1927 12137
rect 1839 12033 1868 12079
rect 1914 12033 1927 12079
rect 1839 11975 1927 12033
rect 1839 11929 1868 11975
rect 1914 11929 1927 11975
rect 1839 11871 1927 11929
rect 1839 11825 1868 11871
rect 1914 11825 1927 11871
rect 1839 11767 1927 11825
rect 1839 11721 1868 11767
rect 1914 11721 1927 11767
rect 1839 11663 1927 11721
rect 1839 11617 1868 11663
rect 1914 11617 1927 11663
rect 1839 11558 1927 11617
rect 1839 11512 1868 11558
rect 1914 11512 1927 11558
rect 1839 11453 1927 11512
rect 1839 11407 1868 11453
rect 1914 11407 1927 11453
rect 1839 11348 1927 11407
rect 1839 11302 1868 11348
rect 1914 11302 1927 11348
rect 1839 11243 1927 11302
rect 1839 11197 1868 11243
rect 1914 11197 1927 11243
rect 1839 11138 1927 11197
rect 1839 11092 1868 11138
rect 1914 11092 1927 11138
rect 1839 11033 1927 11092
rect 1839 10987 1868 11033
rect 1914 10987 1927 11033
rect 1839 10928 1927 10987
rect 1839 10882 1868 10928
rect 1914 10882 1927 10928
rect 1839 10823 1927 10882
rect 1839 10777 1868 10823
rect 1914 10777 1927 10823
rect 1839 10718 1927 10777
rect 1839 10672 1868 10718
rect 1914 10672 1927 10718
rect 1839 10613 1927 10672
rect 1839 10567 1868 10613
rect 1914 10567 1927 10613
rect 1839 10508 1927 10567
rect 1839 10462 1868 10508
rect 1914 10462 1927 10508
rect 1839 10403 1927 10462
rect 1839 10357 1868 10403
rect 1914 10357 1927 10403
rect 1839 10344 1927 10357
rect 2468 9977 2556 9990
rect 2468 9931 2481 9977
rect 2527 9931 2556 9977
rect 495 9891 583 9904
rect 1616 9891 1704 9904
rect 1616 9845 1629 9891
rect 1675 9845 1704 9891
rect 898 9791 986 9804
rect 898 9745 911 9791
rect 957 9745 986 9791
rect 898 9671 986 9745
rect 898 9625 911 9671
rect 957 9625 986 9671
rect 898 9612 986 9625
rect 1106 9791 1194 9804
rect 1106 9745 1135 9791
rect 1181 9745 1194 9791
rect 1106 9671 1194 9745
rect 1616 9771 1704 9845
rect 1616 9725 1629 9771
rect 1675 9725 1704 9771
rect 1616 9712 1704 9725
rect 1824 9891 1912 9904
rect 1824 9845 1853 9891
rect 1899 9845 1912 9891
rect 1824 9771 1912 9845
rect 1824 9725 1853 9771
rect 1899 9725 1912 9771
rect 1824 9712 1912 9725
rect 2468 9849 2556 9931
rect 2468 9803 2481 9849
rect 2527 9803 2556 9849
rect 2468 9722 2556 9803
rect 1106 9625 1135 9671
rect 1181 9625 1194 9671
rect 1106 9612 1194 9625
rect 2468 9676 2481 9722
rect 2527 9676 2556 9722
rect 2468 9595 2556 9676
rect 2468 9549 2481 9595
rect 2527 9549 2556 9595
rect 2468 9536 2556 9549
rect 2676 9977 2764 9990
rect 2676 9931 2705 9977
rect 2751 9931 2764 9977
rect 2676 9849 2764 9931
rect 2676 9803 2705 9849
rect 2751 9803 2764 9849
rect 2676 9722 2764 9803
rect 2676 9676 2705 9722
rect 2751 9676 2764 9722
rect 2676 9595 2764 9676
rect 2676 9549 2705 9595
rect 2751 9549 2764 9595
rect 2676 9536 2764 9549
rect 788 8150 876 8163
rect 788 8104 801 8150
rect 847 8104 876 8150
rect 788 8030 876 8104
rect 788 7984 801 8030
rect 847 7984 876 8030
rect 788 7971 876 7984
rect 996 8150 1100 8163
rect 996 8104 1025 8150
rect 1071 8104 1100 8150
rect 996 8030 1100 8104
rect 996 7984 1025 8030
rect 1071 7984 1100 8030
rect 996 7971 1100 7984
rect 1220 8150 1308 8163
rect 1220 8104 1249 8150
rect 1295 8104 1308 8150
rect 1220 8030 1308 8104
rect 1220 7984 1249 8030
rect 1295 7984 1308 8030
rect 1220 7971 1308 7984
rect 1616 8129 1704 8142
rect 1616 8083 1629 8129
rect 1675 8083 1704 8129
rect 1616 8009 1704 8083
rect 1616 7963 1629 8009
rect 1675 7963 1704 8009
rect 1616 7950 1704 7963
rect 1824 8129 1928 8142
rect 1824 8083 1853 8129
rect 1899 8083 1928 8129
rect 1824 8009 1928 8083
rect 1824 7963 1853 8009
rect 1899 7963 1928 8009
rect 1824 7950 1928 7963
rect 2048 8129 2136 8142
rect 2048 8083 2077 8129
rect 2123 8083 2136 8129
rect 2048 8009 2136 8083
rect 2048 7963 2077 8009
rect 2123 7963 2136 8009
rect 2048 7950 2136 7963
<< mvpdiff >>
rect 601 28581 769 28626
rect 601 28535 692 28581
rect 738 28535 769 28581
rect 601 28399 769 28535
rect 601 28353 692 28399
rect 738 28353 769 28399
rect 601 28218 769 28353
rect 601 28172 692 28218
rect 738 28172 769 28218
rect 601 28036 769 28172
rect 601 27990 692 28036
rect 738 27990 769 28036
rect 601 27944 769 27990
rect 889 28581 993 28626
rect 889 28535 918 28581
rect 964 28535 993 28581
rect 889 28399 993 28535
rect 889 28353 918 28399
rect 964 28353 993 28399
rect 889 28218 993 28353
rect 889 28172 918 28218
rect 964 28172 993 28218
rect 889 28036 993 28172
rect 889 27990 918 28036
rect 964 27990 993 28036
rect 889 27944 993 27990
rect 1113 28581 1389 28626
rect 1113 28535 1228 28581
rect 1274 28535 1389 28581
rect 1113 28399 1389 28535
rect 1113 28353 1228 28399
rect 1274 28353 1389 28399
rect 1113 28218 1389 28353
rect 1113 28172 1228 28218
rect 1274 28172 1389 28218
rect 1113 28036 1389 28172
rect 1113 27990 1228 28036
rect 1274 27990 1389 28036
rect 1113 27944 1389 27990
rect 1509 28581 1613 28626
rect 1509 28535 1538 28581
rect 1584 28535 1613 28581
rect 1509 28399 1613 28535
rect 1509 28353 1538 28399
rect 1584 28353 1613 28399
rect 1509 28218 1613 28353
rect 1509 28172 1538 28218
rect 1584 28172 1613 28218
rect 1509 28036 1613 28172
rect 1509 27990 1538 28036
rect 1584 27990 1613 28036
rect 1509 27944 1613 27990
rect 1733 28581 2008 28626
rect 1733 28535 1764 28581
rect 1810 28535 1931 28581
rect 1977 28535 2008 28581
rect 1733 28399 2008 28535
rect 1733 28353 1764 28399
rect 1810 28353 1931 28399
rect 1977 28353 2008 28399
rect 1733 28218 2008 28353
rect 1733 28172 1764 28218
rect 1810 28172 1931 28218
rect 1977 28172 2008 28218
rect 1733 28036 2008 28172
rect 1733 27990 1764 28036
rect 1810 27990 1931 28036
rect 1977 27990 2008 28036
rect 1733 27944 2008 27990
rect 2128 28581 2232 28626
rect 2128 28535 2157 28581
rect 2203 28535 2232 28581
rect 2128 28399 2232 28535
rect 2128 28353 2157 28399
rect 2203 28353 2232 28399
rect 2128 28218 2232 28353
rect 2128 28172 2157 28218
rect 2203 28172 2232 28218
rect 2128 28036 2232 28172
rect 2128 27990 2157 28036
rect 2203 27990 2232 28036
rect 2128 27944 2232 27990
rect 2352 28581 2628 28626
rect 2352 28535 2467 28581
rect 2513 28535 2628 28581
rect 2352 28399 2628 28535
rect 2352 28353 2467 28399
rect 2513 28353 2628 28399
rect 2352 28218 2628 28353
rect 2352 28172 2467 28218
rect 2513 28172 2628 28218
rect 2352 28036 2628 28172
rect 2352 27990 2467 28036
rect 2513 27990 2628 28036
rect 2352 27944 2628 27990
rect 2748 28581 2852 28626
rect 2748 28535 2777 28581
rect 2823 28535 2852 28581
rect 2748 28399 2852 28535
rect 2748 28353 2777 28399
rect 2823 28353 2852 28399
rect 2748 28218 2852 28353
rect 2748 28172 2777 28218
rect 2823 28172 2852 28218
rect 2748 28036 2852 28172
rect 2748 27990 2777 28036
rect 2823 27990 2852 28036
rect 2748 27944 2852 27990
rect 2972 28581 3246 28626
rect 2972 28535 3003 28581
rect 3049 28535 3169 28581
rect 3215 28535 3246 28581
rect 2972 28399 3246 28535
rect 2972 28353 3003 28399
rect 3049 28353 3169 28399
rect 3215 28353 3246 28399
rect 2972 28218 3246 28353
rect 2972 28172 3003 28218
rect 3049 28172 3169 28218
rect 3215 28172 3246 28218
rect 2972 28036 3246 28172
rect 2972 27990 3003 28036
rect 3049 27990 3169 28036
rect 3215 27990 3246 28036
rect 2972 27944 3246 27990
rect 3366 28581 3470 28626
rect 3366 28535 3395 28581
rect 3441 28535 3470 28581
rect 3366 28399 3470 28535
rect 3366 28353 3395 28399
rect 3441 28353 3470 28399
rect 3366 28218 3470 28353
rect 3366 28172 3395 28218
rect 3441 28172 3470 28218
rect 3366 28036 3470 28172
rect 3366 27990 3395 28036
rect 3441 27990 3470 28036
rect 3366 27944 3470 27990
rect 3590 28581 3866 28626
rect 3590 28535 3705 28581
rect 3751 28535 3866 28581
rect 3590 28399 3866 28535
rect 3590 28353 3705 28399
rect 3751 28353 3866 28399
rect 3590 28218 3866 28353
rect 3590 28172 3705 28218
rect 3751 28172 3866 28218
rect 3590 28036 3866 28172
rect 3590 27990 3705 28036
rect 3751 27990 3866 28036
rect 3590 27944 3866 27990
rect 3986 28581 4090 28626
rect 3986 28535 4015 28581
rect 4061 28535 4090 28581
rect 3986 28399 4090 28535
rect 3986 28353 4015 28399
rect 4061 28353 4090 28399
rect 3986 28218 4090 28353
rect 3986 28172 4015 28218
rect 4061 28172 4090 28218
rect 3986 28036 4090 28172
rect 3986 27990 4015 28036
rect 4061 27990 4090 28036
rect 3986 27944 4090 27990
rect 4210 28581 4485 28626
rect 4210 28535 4241 28581
rect 4287 28535 4408 28581
rect 4454 28535 4485 28581
rect 4210 28399 4485 28535
rect 4210 28353 4241 28399
rect 4287 28353 4408 28399
rect 4454 28353 4485 28399
rect 4210 28218 4485 28353
rect 4210 28172 4241 28218
rect 4287 28172 4408 28218
rect 4454 28172 4485 28218
rect 4210 28036 4485 28172
rect 4210 27990 4241 28036
rect 4287 27990 4408 28036
rect 4454 27990 4485 28036
rect 4210 27944 4485 27990
rect 4605 28581 4709 28626
rect 4605 28535 4634 28581
rect 4680 28535 4709 28581
rect 4605 28399 4709 28535
rect 4605 28353 4634 28399
rect 4680 28353 4709 28399
rect 4605 28218 4709 28353
rect 4605 28172 4634 28218
rect 4680 28172 4709 28218
rect 4605 28036 4709 28172
rect 4605 27990 4634 28036
rect 4680 27990 4709 28036
rect 4605 27944 4709 27990
rect 4829 28581 5069 28626
rect 4829 28535 4944 28581
rect 4990 28535 5069 28581
rect 4829 28399 5069 28535
rect 4829 28353 4944 28399
rect 4990 28353 5069 28399
rect 4829 28218 5069 28353
rect 4829 28172 4944 28218
rect 4990 28172 5069 28218
rect 4829 28036 5069 28172
rect 4829 27990 4944 28036
rect 4990 27990 5069 28036
rect 4829 27944 5069 27990
rect 5189 28581 5294 28626
rect 5189 28535 5219 28581
rect 5265 28535 5294 28581
rect 5189 28399 5294 28535
rect 5189 28353 5219 28399
rect 5265 28353 5294 28399
rect 5189 28218 5294 28353
rect 5189 28172 5219 28218
rect 5265 28172 5294 28218
rect 5189 28036 5294 28172
rect 5189 27990 5219 28036
rect 5265 27990 5294 28036
rect 5189 27944 5294 27990
rect 5414 28581 5618 28626
rect 5414 28535 5480 28581
rect 5526 28535 5618 28581
rect 5414 28399 5618 28535
rect 5414 28353 5480 28399
rect 5526 28353 5618 28399
rect 5414 28218 5618 28353
rect 5414 28172 5480 28218
rect 5526 28172 5618 28218
rect 5414 28036 5618 28172
rect 5414 27990 5480 28036
rect 5526 27990 5618 28036
rect 5414 27944 5618 27990
rect 601 27805 769 27851
rect 601 27759 692 27805
rect 738 27759 769 27805
rect 601 27624 769 27759
rect 601 27578 692 27624
rect 738 27578 769 27624
rect 601 27443 769 27578
rect 601 27397 692 27443
rect 738 27397 769 27443
rect 601 27261 769 27397
rect 601 27215 692 27261
rect 738 27215 769 27261
rect 601 27169 769 27215
rect 889 27805 993 27851
rect 889 27759 918 27805
rect 964 27759 993 27805
rect 889 27624 993 27759
rect 889 27578 918 27624
rect 964 27578 993 27624
rect 889 27443 993 27578
rect 889 27397 918 27443
rect 964 27397 993 27443
rect 889 27261 993 27397
rect 889 27215 918 27261
rect 964 27215 993 27261
rect 889 27169 993 27215
rect 1113 27805 1389 27851
rect 1113 27759 1228 27805
rect 1274 27759 1389 27805
rect 1113 27624 1389 27759
rect 1113 27578 1228 27624
rect 1274 27578 1389 27624
rect 1113 27443 1389 27578
rect 1113 27397 1228 27443
rect 1274 27397 1389 27443
rect 1113 27261 1389 27397
rect 1113 27215 1228 27261
rect 1274 27215 1389 27261
rect 1113 27169 1389 27215
rect 1509 27805 1613 27851
rect 1509 27759 1538 27805
rect 1584 27759 1613 27805
rect 1509 27624 1613 27759
rect 1509 27578 1538 27624
rect 1584 27578 1613 27624
rect 1509 27443 1613 27578
rect 1509 27397 1538 27443
rect 1584 27397 1613 27443
rect 1509 27261 1613 27397
rect 1509 27215 1538 27261
rect 1584 27215 1613 27261
rect 1509 27169 1613 27215
rect 1733 27805 2008 27851
rect 1733 27759 1764 27805
rect 1810 27759 1931 27805
rect 1977 27759 2008 27805
rect 1733 27624 2008 27759
rect 1733 27578 1764 27624
rect 1810 27578 1931 27624
rect 1977 27578 2008 27624
rect 1733 27443 2008 27578
rect 1733 27397 1764 27443
rect 1810 27397 1931 27443
rect 1977 27397 2008 27443
rect 1733 27261 2008 27397
rect 1733 27215 1764 27261
rect 1810 27215 1931 27261
rect 1977 27215 2008 27261
rect 1733 27169 2008 27215
rect 2128 27805 2232 27851
rect 2128 27759 2157 27805
rect 2203 27759 2232 27805
rect 2128 27624 2232 27759
rect 2128 27578 2157 27624
rect 2203 27578 2232 27624
rect 2128 27443 2232 27578
rect 2128 27397 2157 27443
rect 2203 27397 2232 27443
rect 2128 27261 2232 27397
rect 2128 27215 2157 27261
rect 2203 27215 2232 27261
rect 2128 27169 2232 27215
rect 2352 27805 2628 27851
rect 2352 27759 2467 27805
rect 2513 27759 2628 27805
rect 2352 27624 2628 27759
rect 2352 27578 2467 27624
rect 2513 27578 2628 27624
rect 2352 27443 2628 27578
rect 2352 27397 2467 27443
rect 2513 27397 2628 27443
rect 2352 27261 2628 27397
rect 2352 27215 2467 27261
rect 2513 27215 2628 27261
rect 2352 27169 2628 27215
rect 2748 27805 2852 27851
rect 2748 27759 2777 27805
rect 2823 27759 2852 27805
rect 2748 27624 2852 27759
rect 2748 27578 2777 27624
rect 2823 27578 2852 27624
rect 2748 27443 2852 27578
rect 2748 27397 2777 27443
rect 2823 27397 2852 27443
rect 2748 27261 2852 27397
rect 2748 27215 2777 27261
rect 2823 27215 2852 27261
rect 2748 27169 2852 27215
rect 2972 27805 3246 27851
rect 2972 27759 3003 27805
rect 3049 27759 3169 27805
rect 3215 27759 3246 27805
rect 2972 27624 3246 27759
rect 2972 27578 3003 27624
rect 3049 27578 3169 27624
rect 3215 27578 3246 27624
rect 2972 27443 3246 27578
rect 2972 27397 3003 27443
rect 3049 27397 3169 27443
rect 3215 27397 3246 27443
rect 2972 27261 3246 27397
rect 2972 27215 3003 27261
rect 3049 27215 3169 27261
rect 3215 27215 3246 27261
rect 2972 27169 3246 27215
rect 3366 27805 3470 27851
rect 3366 27759 3395 27805
rect 3441 27759 3470 27805
rect 3366 27624 3470 27759
rect 3366 27578 3395 27624
rect 3441 27578 3470 27624
rect 3366 27443 3470 27578
rect 3366 27397 3395 27443
rect 3441 27397 3470 27443
rect 3366 27261 3470 27397
rect 3366 27215 3395 27261
rect 3441 27215 3470 27261
rect 3366 27169 3470 27215
rect 3590 27805 3866 27851
rect 3590 27759 3705 27805
rect 3751 27759 3866 27805
rect 3590 27624 3866 27759
rect 3590 27578 3705 27624
rect 3751 27578 3866 27624
rect 3590 27443 3866 27578
rect 3590 27397 3705 27443
rect 3751 27397 3866 27443
rect 3590 27261 3866 27397
rect 3590 27215 3705 27261
rect 3751 27215 3866 27261
rect 3590 27169 3866 27215
rect 3986 27805 4090 27851
rect 3986 27759 4015 27805
rect 4061 27759 4090 27805
rect 3986 27624 4090 27759
rect 3986 27578 4015 27624
rect 4061 27578 4090 27624
rect 3986 27443 4090 27578
rect 3986 27397 4015 27443
rect 4061 27397 4090 27443
rect 3986 27261 4090 27397
rect 3986 27215 4015 27261
rect 4061 27215 4090 27261
rect 3986 27169 4090 27215
rect 4210 27805 4485 27851
rect 4210 27759 4241 27805
rect 4287 27759 4408 27805
rect 4454 27759 4485 27805
rect 4210 27624 4485 27759
rect 4210 27578 4241 27624
rect 4287 27578 4408 27624
rect 4454 27578 4485 27624
rect 4210 27443 4485 27578
rect 4210 27397 4241 27443
rect 4287 27397 4408 27443
rect 4454 27397 4485 27443
rect 4210 27261 4485 27397
rect 4210 27215 4241 27261
rect 4287 27215 4408 27261
rect 4454 27215 4485 27261
rect 4210 27169 4485 27215
rect 4605 27805 4709 27851
rect 4605 27759 4634 27805
rect 4680 27759 4709 27805
rect 4605 27624 4709 27759
rect 4605 27578 4634 27624
rect 4680 27578 4709 27624
rect 4605 27443 4709 27578
rect 4605 27397 4634 27443
rect 4680 27397 4709 27443
rect 4605 27261 4709 27397
rect 4605 27215 4634 27261
rect 4680 27215 4709 27261
rect 4605 27169 4709 27215
rect 4829 27805 5069 27851
rect 4829 27759 4944 27805
rect 4990 27759 5069 27805
rect 4829 27624 5069 27759
rect 4829 27578 4944 27624
rect 4990 27578 5069 27624
rect 4829 27443 5069 27578
rect 4829 27397 4944 27443
rect 4990 27397 5069 27443
rect 4829 27261 5069 27397
rect 4829 27215 4944 27261
rect 4990 27215 5069 27261
rect 4829 27169 5069 27215
rect 5189 27805 5294 27851
rect 5189 27759 5219 27805
rect 5265 27759 5294 27805
rect 5189 27624 5294 27759
rect 5189 27578 5219 27624
rect 5265 27578 5294 27624
rect 5189 27443 5294 27578
rect 5189 27397 5219 27443
rect 5265 27397 5294 27443
rect 5189 27261 5294 27397
rect 5189 27215 5219 27261
rect 5265 27215 5294 27261
rect 5189 27169 5294 27215
rect 5414 27805 5618 27851
rect 5414 27759 5480 27805
rect 5526 27759 5618 27805
rect 5414 27624 5618 27759
rect 5414 27578 5480 27624
rect 5526 27578 5618 27624
rect 5414 27443 5618 27578
rect 5414 27397 5480 27443
rect 5526 27397 5618 27443
rect 5414 27261 5618 27397
rect 5414 27215 5480 27261
rect 5526 27215 5618 27261
rect 5414 27169 5618 27215
rect 795 26937 883 26950
rect 795 26891 808 26937
rect 854 26891 883 26937
rect 795 26829 883 26891
rect 795 26783 808 26829
rect 854 26783 883 26829
rect 795 26721 883 26783
rect 795 26675 808 26721
rect 854 26675 883 26721
rect 795 26613 883 26675
rect 795 26567 808 26613
rect 854 26567 883 26613
rect 795 26505 883 26567
rect 795 26459 808 26505
rect 854 26459 883 26505
rect 795 26397 883 26459
rect 795 26351 808 26397
rect 854 26351 883 26397
rect 795 26289 883 26351
rect 795 26243 808 26289
rect 854 26243 883 26289
rect 795 26182 883 26243
rect 795 26136 808 26182
rect 854 26136 883 26182
rect 795 26075 883 26136
rect 795 26029 808 26075
rect 854 26029 883 26075
rect 795 25968 883 26029
rect 795 25922 808 25968
rect 854 25922 883 25968
rect 795 25861 883 25922
rect 795 25815 808 25861
rect 854 25815 883 25861
rect 795 25754 883 25815
rect 795 25708 808 25754
rect 854 25708 883 25754
rect 795 25647 883 25708
rect 795 25601 808 25647
rect 854 25601 883 25647
rect 795 25588 883 25601
rect 1003 26937 1091 26950
rect 1003 26891 1032 26937
rect 1078 26891 1091 26937
rect 1003 26829 1091 26891
rect 1003 26783 1032 26829
rect 1078 26783 1091 26829
rect 1003 26721 1091 26783
rect 1003 26675 1032 26721
rect 1078 26675 1091 26721
rect 1003 26613 1091 26675
rect 1003 26567 1032 26613
rect 1078 26567 1091 26613
rect 1003 26505 1091 26567
rect 1003 26459 1032 26505
rect 1078 26459 1091 26505
rect 1003 26397 1091 26459
rect 1003 26351 1032 26397
rect 1078 26351 1091 26397
rect 1003 26289 1091 26351
rect 1003 26243 1032 26289
rect 1078 26243 1091 26289
rect 1003 26182 1091 26243
rect 1003 26136 1032 26182
rect 1078 26136 1091 26182
rect 1003 26075 1091 26136
rect 1003 26029 1032 26075
rect 1078 26029 1091 26075
rect 1003 25968 1091 26029
rect 1003 25922 1032 25968
rect 1078 25922 1091 25968
rect 1003 25861 1091 25922
rect 1003 25815 1032 25861
rect 1078 25815 1091 25861
rect 1003 25754 1091 25815
rect 1003 25708 1032 25754
rect 1078 25708 1091 25754
rect 1003 25647 1091 25708
rect 1003 25601 1032 25647
rect 1078 25601 1091 25647
rect 1003 25588 1091 25601
rect 1411 26937 1499 26950
rect 1411 26891 1424 26937
rect 1470 26891 1499 26937
rect 1411 26829 1499 26891
rect 1411 26783 1424 26829
rect 1470 26783 1499 26829
rect 1411 26721 1499 26783
rect 1411 26675 1424 26721
rect 1470 26675 1499 26721
rect 1411 26613 1499 26675
rect 1411 26567 1424 26613
rect 1470 26567 1499 26613
rect 1411 26505 1499 26567
rect 1411 26459 1424 26505
rect 1470 26459 1499 26505
rect 1411 26397 1499 26459
rect 1411 26351 1424 26397
rect 1470 26351 1499 26397
rect 1411 26289 1499 26351
rect 1411 26243 1424 26289
rect 1470 26243 1499 26289
rect 1411 26182 1499 26243
rect 1411 26136 1424 26182
rect 1470 26136 1499 26182
rect 1411 26075 1499 26136
rect 1411 26029 1424 26075
rect 1470 26029 1499 26075
rect 1411 25968 1499 26029
rect 1411 25922 1424 25968
rect 1470 25922 1499 25968
rect 1411 25861 1499 25922
rect 1411 25815 1424 25861
rect 1470 25815 1499 25861
rect 1411 25754 1499 25815
rect 1411 25708 1424 25754
rect 1470 25708 1499 25754
rect 1411 25647 1499 25708
rect 1411 25601 1424 25647
rect 1470 25601 1499 25647
rect 1411 25588 1499 25601
rect 1619 26937 1707 26950
rect 1619 26891 1648 26937
rect 1694 26891 1707 26937
rect 1619 26829 1707 26891
rect 1619 26783 1648 26829
rect 1694 26783 1707 26829
rect 1619 26721 1707 26783
rect 1619 26675 1648 26721
rect 1694 26675 1707 26721
rect 1619 26613 1707 26675
rect 1619 26567 1648 26613
rect 1694 26567 1707 26613
rect 1619 26505 1707 26567
rect 1619 26459 1648 26505
rect 1694 26459 1707 26505
rect 1619 26397 1707 26459
rect 1619 26351 1648 26397
rect 1694 26351 1707 26397
rect 1619 26289 1707 26351
rect 1619 26243 1648 26289
rect 1694 26243 1707 26289
rect 1619 26182 1707 26243
rect 1619 26136 1648 26182
rect 1694 26136 1707 26182
rect 1619 26075 1707 26136
rect 1619 26029 1648 26075
rect 1694 26029 1707 26075
rect 1619 25968 1707 26029
rect 1619 25922 1648 25968
rect 1694 25922 1707 25968
rect 1619 25861 1707 25922
rect 1619 25815 1648 25861
rect 1694 25815 1707 25861
rect 1619 25754 1707 25815
rect 1619 25708 1648 25754
rect 1694 25708 1707 25754
rect 1619 25647 1707 25708
rect 1619 25601 1648 25647
rect 1694 25601 1707 25647
rect 1619 25588 1707 25601
rect 2034 26937 2122 26950
rect 2034 26891 2047 26937
rect 2093 26891 2122 26937
rect 2034 26829 2122 26891
rect 2034 26783 2047 26829
rect 2093 26783 2122 26829
rect 2034 26721 2122 26783
rect 2034 26675 2047 26721
rect 2093 26675 2122 26721
rect 2034 26613 2122 26675
rect 2034 26567 2047 26613
rect 2093 26567 2122 26613
rect 2034 26505 2122 26567
rect 2034 26459 2047 26505
rect 2093 26459 2122 26505
rect 2034 26397 2122 26459
rect 2034 26351 2047 26397
rect 2093 26351 2122 26397
rect 2034 26289 2122 26351
rect 2034 26243 2047 26289
rect 2093 26243 2122 26289
rect 2034 26182 2122 26243
rect 2034 26136 2047 26182
rect 2093 26136 2122 26182
rect 2034 26075 2122 26136
rect 2034 26029 2047 26075
rect 2093 26029 2122 26075
rect 2034 25968 2122 26029
rect 2034 25922 2047 25968
rect 2093 25922 2122 25968
rect 2034 25861 2122 25922
rect 2034 25815 2047 25861
rect 2093 25815 2122 25861
rect 2034 25754 2122 25815
rect 2034 25708 2047 25754
rect 2093 25708 2122 25754
rect 2034 25647 2122 25708
rect 2034 25601 2047 25647
rect 2093 25601 2122 25647
rect 2034 25588 2122 25601
rect 2242 26937 2330 26950
rect 2242 26891 2271 26937
rect 2317 26891 2330 26937
rect 2242 26829 2330 26891
rect 2242 26783 2271 26829
rect 2317 26783 2330 26829
rect 2242 26721 2330 26783
rect 2242 26675 2271 26721
rect 2317 26675 2330 26721
rect 2242 26613 2330 26675
rect 2242 26567 2271 26613
rect 2317 26567 2330 26613
rect 2242 26505 2330 26567
rect 2242 26459 2271 26505
rect 2317 26459 2330 26505
rect 2242 26397 2330 26459
rect 2242 26351 2271 26397
rect 2317 26351 2330 26397
rect 2242 26289 2330 26351
rect 2242 26243 2271 26289
rect 2317 26243 2330 26289
rect 2242 26182 2330 26243
rect 2242 26136 2271 26182
rect 2317 26136 2330 26182
rect 2242 26075 2330 26136
rect 2242 26029 2271 26075
rect 2317 26029 2330 26075
rect 2242 25968 2330 26029
rect 2242 25922 2271 25968
rect 2317 25922 2330 25968
rect 2242 25861 2330 25922
rect 2242 25815 2271 25861
rect 2317 25815 2330 25861
rect 2242 25754 2330 25815
rect 2242 25708 2271 25754
rect 2317 25708 2330 25754
rect 2242 25647 2330 25708
rect 2242 25601 2271 25647
rect 2317 25601 2330 25647
rect 2242 25588 2330 25601
rect 2650 26937 2738 26950
rect 2650 26891 2663 26937
rect 2709 26891 2738 26937
rect 2650 26829 2738 26891
rect 2650 26783 2663 26829
rect 2709 26783 2738 26829
rect 2650 26721 2738 26783
rect 2650 26675 2663 26721
rect 2709 26675 2738 26721
rect 2650 26613 2738 26675
rect 2650 26567 2663 26613
rect 2709 26567 2738 26613
rect 2650 26505 2738 26567
rect 2650 26459 2663 26505
rect 2709 26459 2738 26505
rect 2650 26397 2738 26459
rect 2650 26351 2663 26397
rect 2709 26351 2738 26397
rect 2650 26289 2738 26351
rect 2650 26243 2663 26289
rect 2709 26243 2738 26289
rect 2650 26182 2738 26243
rect 2650 26136 2663 26182
rect 2709 26136 2738 26182
rect 2650 26075 2738 26136
rect 2650 26029 2663 26075
rect 2709 26029 2738 26075
rect 2650 25968 2738 26029
rect 2650 25922 2663 25968
rect 2709 25922 2738 25968
rect 2650 25861 2738 25922
rect 2650 25815 2663 25861
rect 2709 25815 2738 25861
rect 2650 25754 2738 25815
rect 2650 25708 2663 25754
rect 2709 25708 2738 25754
rect 2650 25647 2738 25708
rect 2650 25601 2663 25647
rect 2709 25601 2738 25647
rect 2650 25588 2738 25601
rect 2858 26937 2946 26950
rect 2858 26891 2887 26937
rect 2933 26891 2946 26937
rect 2858 26829 2946 26891
rect 2858 26783 2887 26829
rect 2933 26783 2946 26829
rect 2858 26721 2946 26783
rect 2858 26675 2887 26721
rect 2933 26675 2946 26721
rect 2858 26613 2946 26675
rect 2858 26567 2887 26613
rect 2933 26567 2946 26613
rect 2858 26505 2946 26567
rect 2858 26459 2887 26505
rect 2933 26459 2946 26505
rect 2858 26397 2946 26459
rect 2858 26351 2887 26397
rect 2933 26351 2946 26397
rect 2858 26289 2946 26351
rect 2858 26243 2887 26289
rect 2933 26243 2946 26289
rect 2858 26182 2946 26243
rect 2858 26136 2887 26182
rect 2933 26136 2946 26182
rect 2858 26075 2946 26136
rect 2858 26029 2887 26075
rect 2933 26029 2946 26075
rect 2858 25968 2946 26029
rect 2858 25922 2887 25968
rect 2933 25922 2946 25968
rect 2858 25861 2946 25922
rect 2858 25815 2887 25861
rect 2933 25815 2946 25861
rect 2858 25754 2946 25815
rect 2858 25708 2887 25754
rect 2933 25708 2946 25754
rect 2858 25647 2946 25708
rect 2858 25601 2887 25647
rect 2933 25601 2946 25647
rect 2858 25588 2946 25601
rect 3272 26937 3360 26950
rect 3272 26891 3285 26937
rect 3331 26891 3360 26937
rect 3272 26829 3360 26891
rect 3272 26783 3285 26829
rect 3331 26783 3360 26829
rect 3272 26721 3360 26783
rect 3272 26675 3285 26721
rect 3331 26675 3360 26721
rect 3272 26613 3360 26675
rect 3272 26567 3285 26613
rect 3331 26567 3360 26613
rect 3272 26505 3360 26567
rect 3272 26459 3285 26505
rect 3331 26459 3360 26505
rect 3272 26397 3360 26459
rect 3272 26351 3285 26397
rect 3331 26351 3360 26397
rect 3272 26289 3360 26351
rect 3272 26243 3285 26289
rect 3331 26243 3360 26289
rect 3272 26182 3360 26243
rect 3272 26136 3285 26182
rect 3331 26136 3360 26182
rect 3272 26075 3360 26136
rect 3272 26029 3285 26075
rect 3331 26029 3360 26075
rect 3272 25968 3360 26029
rect 3272 25922 3285 25968
rect 3331 25922 3360 25968
rect 3272 25861 3360 25922
rect 3272 25815 3285 25861
rect 3331 25815 3360 25861
rect 3272 25754 3360 25815
rect 3272 25708 3285 25754
rect 3331 25708 3360 25754
rect 3272 25647 3360 25708
rect 3272 25601 3285 25647
rect 3331 25601 3360 25647
rect 3272 25588 3360 25601
rect 3480 26937 3568 26950
rect 3480 26891 3509 26937
rect 3555 26891 3568 26937
rect 3480 26829 3568 26891
rect 3480 26783 3509 26829
rect 3555 26783 3568 26829
rect 3480 26721 3568 26783
rect 3480 26675 3509 26721
rect 3555 26675 3568 26721
rect 3480 26613 3568 26675
rect 3480 26567 3509 26613
rect 3555 26567 3568 26613
rect 3480 26505 3568 26567
rect 3480 26459 3509 26505
rect 3555 26459 3568 26505
rect 3480 26397 3568 26459
rect 3480 26351 3509 26397
rect 3555 26351 3568 26397
rect 3480 26289 3568 26351
rect 3480 26243 3509 26289
rect 3555 26243 3568 26289
rect 3480 26182 3568 26243
rect 3480 26136 3509 26182
rect 3555 26136 3568 26182
rect 3480 26075 3568 26136
rect 3480 26029 3509 26075
rect 3555 26029 3568 26075
rect 3480 25968 3568 26029
rect 3480 25922 3509 25968
rect 3555 25922 3568 25968
rect 3480 25861 3568 25922
rect 3480 25815 3509 25861
rect 3555 25815 3568 25861
rect 3480 25754 3568 25815
rect 3480 25708 3509 25754
rect 3555 25708 3568 25754
rect 3480 25647 3568 25708
rect 3480 25601 3509 25647
rect 3555 25601 3568 25647
rect 3480 25588 3568 25601
rect 3888 26937 3976 26950
rect 3888 26891 3901 26937
rect 3947 26891 3976 26937
rect 3888 26829 3976 26891
rect 3888 26783 3901 26829
rect 3947 26783 3976 26829
rect 3888 26721 3976 26783
rect 3888 26675 3901 26721
rect 3947 26675 3976 26721
rect 3888 26613 3976 26675
rect 3888 26567 3901 26613
rect 3947 26567 3976 26613
rect 3888 26505 3976 26567
rect 3888 26459 3901 26505
rect 3947 26459 3976 26505
rect 3888 26397 3976 26459
rect 3888 26351 3901 26397
rect 3947 26351 3976 26397
rect 3888 26289 3976 26351
rect 3888 26243 3901 26289
rect 3947 26243 3976 26289
rect 3888 26182 3976 26243
rect 3888 26136 3901 26182
rect 3947 26136 3976 26182
rect 3888 26075 3976 26136
rect 3888 26029 3901 26075
rect 3947 26029 3976 26075
rect 3888 25968 3976 26029
rect 3888 25922 3901 25968
rect 3947 25922 3976 25968
rect 3888 25861 3976 25922
rect 3888 25815 3901 25861
rect 3947 25815 3976 25861
rect 3888 25754 3976 25815
rect 3888 25708 3901 25754
rect 3947 25708 3976 25754
rect 3888 25647 3976 25708
rect 3888 25601 3901 25647
rect 3947 25601 3976 25647
rect 3888 25588 3976 25601
rect 4096 26937 4184 26950
rect 4096 26891 4125 26937
rect 4171 26891 4184 26937
rect 4096 26829 4184 26891
rect 4096 26783 4125 26829
rect 4171 26783 4184 26829
rect 4096 26721 4184 26783
rect 4096 26675 4125 26721
rect 4171 26675 4184 26721
rect 4096 26613 4184 26675
rect 4096 26567 4125 26613
rect 4171 26567 4184 26613
rect 4096 26505 4184 26567
rect 4096 26459 4125 26505
rect 4171 26459 4184 26505
rect 4096 26397 4184 26459
rect 4096 26351 4125 26397
rect 4171 26351 4184 26397
rect 4096 26289 4184 26351
rect 4096 26243 4125 26289
rect 4171 26243 4184 26289
rect 4096 26182 4184 26243
rect 4096 26136 4125 26182
rect 4171 26136 4184 26182
rect 4096 26075 4184 26136
rect 4096 26029 4125 26075
rect 4171 26029 4184 26075
rect 4096 25968 4184 26029
rect 4096 25922 4125 25968
rect 4171 25922 4184 25968
rect 4096 25861 4184 25922
rect 4096 25815 4125 25861
rect 4171 25815 4184 25861
rect 4096 25754 4184 25815
rect 4096 25708 4125 25754
rect 4171 25708 4184 25754
rect 4096 25647 4184 25708
rect 4096 25601 4125 25647
rect 4171 25601 4184 25647
rect 4096 25588 4184 25601
rect 4511 26937 4599 26950
rect 4511 26891 4524 26937
rect 4570 26891 4599 26937
rect 4511 26829 4599 26891
rect 4511 26783 4524 26829
rect 4570 26783 4599 26829
rect 4511 26721 4599 26783
rect 4511 26675 4524 26721
rect 4570 26675 4599 26721
rect 4511 26613 4599 26675
rect 4511 26567 4524 26613
rect 4570 26567 4599 26613
rect 4511 26505 4599 26567
rect 4511 26459 4524 26505
rect 4570 26459 4599 26505
rect 4511 26397 4599 26459
rect 4511 26351 4524 26397
rect 4570 26351 4599 26397
rect 4511 26289 4599 26351
rect 4511 26243 4524 26289
rect 4570 26243 4599 26289
rect 4511 26182 4599 26243
rect 4511 26136 4524 26182
rect 4570 26136 4599 26182
rect 4511 26075 4599 26136
rect 4511 26029 4524 26075
rect 4570 26029 4599 26075
rect 4511 25968 4599 26029
rect 4511 25922 4524 25968
rect 4570 25922 4599 25968
rect 4511 25861 4599 25922
rect 4511 25815 4524 25861
rect 4570 25815 4599 25861
rect 4511 25754 4599 25815
rect 4511 25708 4524 25754
rect 4570 25708 4599 25754
rect 4511 25647 4599 25708
rect 4511 25601 4524 25647
rect 4570 25601 4599 25647
rect 4511 25588 4599 25601
rect 4719 26937 4807 26950
rect 4719 26891 4748 26937
rect 4794 26891 4807 26937
rect 4719 26829 4807 26891
rect 4719 26783 4748 26829
rect 4794 26783 4807 26829
rect 4719 26721 4807 26783
rect 4719 26675 4748 26721
rect 4794 26675 4807 26721
rect 4719 26613 4807 26675
rect 4719 26567 4748 26613
rect 4794 26567 4807 26613
rect 4719 26505 4807 26567
rect 4719 26459 4748 26505
rect 4794 26459 4807 26505
rect 4719 26397 4807 26459
rect 4719 26351 4748 26397
rect 4794 26351 4807 26397
rect 4719 26289 4807 26351
rect 4719 26243 4748 26289
rect 4794 26243 4807 26289
rect 4719 26182 4807 26243
rect 4719 26136 4748 26182
rect 4794 26136 4807 26182
rect 4719 26075 4807 26136
rect 4719 26029 4748 26075
rect 4794 26029 4807 26075
rect 4719 25968 4807 26029
rect 4719 25922 4748 25968
rect 4794 25922 4807 25968
rect 4719 25861 4807 25922
rect 4719 25815 4748 25861
rect 4794 25815 4807 25861
rect 4719 25754 4807 25815
rect 4719 25708 4748 25754
rect 4794 25708 4807 25754
rect 4719 25647 4807 25708
rect 4719 25601 4748 25647
rect 4794 25601 4807 25647
rect 4719 25588 4807 25601
rect 5127 26937 5215 26950
rect 5127 26891 5140 26937
rect 5186 26891 5215 26937
rect 5127 26829 5215 26891
rect 5127 26783 5140 26829
rect 5186 26783 5215 26829
rect 5127 26721 5215 26783
rect 5127 26675 5140 26721
rect 5186 26675 5215 26721
rect 5127 26613 5215 26675
rect 5127 26567 5140 26613
rect 5186 26567 5215 26613
rect 5127 26505 5215 26567
rect 5127 26459 5140 26505
rect 5186 26459 5215 26505
rect 5127 26397 5215 26459
rect 5127 26351 5140 26397
rect 5186 26351 5215 26397
rect 5127 26289 5215 26351
rect 5127 26243 5140 26289
rect 5186 26243 5215 26289
rect 5127 26182 5215 26243
rect 5127 26136 5140 26182
rect 5186 26136 5215 26182
rect 5127 26075 5215 26136
rect 5127 26029 5140 26075
rect 5186 26029 5215 26075
rect 5127 25968 5215 26029
rect 5127 25922 5140 25968
rect 5186 25922 5215 25968
rect 5127 25861 5215 25922
rect 5127 25815 5140 25861
rect 5186 25815 5215 25861
rect 5127 25754 5215 25815
rect 5127 25708 5140 25754
rect 5186 25708 5215 25754
rect 5127 25647 5215 25708
rect 5127 25601 5140 25647
rect 5186 25601 5215 25647
rect 5127 25588 5215 25601
rect 5335 26937 5423 26950
rect 5335 26891 5364 26937
rect 5410 26891 5423 26937
rect 5335 26829 5423 26891
rect 5335 26783 5364 26829
rect 5410 26783 5423 26829
rect 5335 26721 5423 26783
rect 5335 26675 5364 26721
rect 5410 26675 5423 26721
rect 5335 26613 5423 26675
rect 5335 26567 5364 26613
rect 5410 26567 5423 26613
rect 5335 26505 5423 26567
rect 5335 26459 5364 26505
rect 5410 26459 5423 26505
rect 5335 26397 5423 26459
rect 5335 26351 5364 26397
rect 5410 26351 5423 26397
rect 5335 26289 5423 26351
rect 5335 26243 5364 26289
rect 5410 26243 5423 26289
rect 5335 26182 5423 26243
rect 5335 26136 5364 26182
rect 5410 26136 5423 26182
rect 5335 26075 5423 26136
rect 5335 26029 5364 26075
rect 5410 26029 5423 26075
rect 5335 25968 5423 26029
rect 5335 25922 5364 25968
rect 5410 25922 5423 25968
rect 5335 25861 5423 25922
rect 5335 25815 5364 25861
rect 5410 25815 5423 25861
rect 5335 25754 5423 25815
rect 5335 25708 5364 25754
rect 5410 25708 5423 25754
rect 5335 25647 5423 25708
rect 5335 25601 5364 25647
rect 5410 25601 5423 25647
rect 5335 25588 5423 25601
rect 793 25350 881 25363
rect 793 25304 806 25350
rect 852 25304 881 25350
rect 793 25242 881 25304
rect 793 25196 806 25242
rect 852 25196 881 25242
rect 793 25134 881 25196
rect 793 25088 806 25134
rect 852 25088 881 25134
rect 793 25026 881 25088
rect 793 24980 806 25026
rect 852 24980 881 25026
rect 793 24918 881 24980
rect 793 24872 806 24918
rect 852 24872 881 24918
rect 793 24810 881 24872
rect 793 24764 806 24810
rect 852 24764 881 24810
rect 793 24702 881 24764
rect 793 24656 806 24702
rect 852 24656 881 24702
rect 793 24595 881 24656
rect 793 24549 806 24595
rect 852 24549 881 24595
rect 793 24488 881 24549
rect 793 24442 806 24488
rect 852 24442 881 24488
rect 793 24381 881 24442
rect 793 24335 806 24381
rect 852 24335 881 24381
rect 793 24274 881 24335
rect 793 24228 806 24274
rect 852 24228 881 24274
rect 793 24167 881 24228
rect 793 24121 806 24167
rect 852 24121 881 24167
rect 793 24060 881 24121
rect 793 24014 806 24060
rect 852 24014 881 24060
rect 793 24001 881 24014
rect 1001 25350 1089 25363
rect 1001 25304 1030 25350
rect 1076 25304 1089 25350
rect 1001 25242 1089 25304
rect 1001 25196 1030 25242
rect 1076 25196 1089 25242
rect 1001 25134 1089 25196
rect 1001 25088 1030 25134
rect 1076 25088 1089 25134
rect 1001 25026 1089 25088
rect 1001 24980 1030 25026
rect 1076 24980 1089 25026
rect 1001 24918 1089 24980
rect 1001 24872 1030 24918
rect 1076 24872 1089 24918
rect 1001 24810 1089 24872
rect 1001 24764 1030 24810
rect 1076 24764 1089 24810
rect 1001 24702 1089 24764
rect 1001 24656 1030 24702
rect 1076 24656 1089 24702
rect 1413 25350 1501 25363
rect 1413 25304 1426 25350
rect 1472 25304 1501 25350
rect 1413 25242 1501 25304
rect 1413 25196 1426 25242
rect 1472 25196 1501 25242
rect 1413 25134 1501 25196
rect 1413 25088 1426 25134
rect 1472 25088 1501 25134
rect 1413 25026 1501 25088
rect 1413 24980 1426 25026
rect 1472 24980 1501 25026
rect 1413 24918 1501 24980
rect 1413 24872 1426 24918
rect 1472 24872 1501 24918
rect 1413 24810 1501 24872
rect 1413 24764 1426 24810
rect 1472 24764 1501 24810
rect 1413 24702 1501 24764
rect 1001 24595 1089 24656
rect 1001 24549 1030 24595
rect 1076 24549 1089 24595
rect 1001 24488 1089 24549
rect 1001 24442 1030 24488
rect 1076 24442 1089 24488
rect 1001 24381 1089 24442
rect 1413 24656 1426 24702
rect 1472 24656 1501 24702
rect 1413 24595 1501 24656
rect 1413 24549 1426 24595
rect 1472 24549 1501 24595
rect 1413 24488 1501 24549
rect 1413 24442 1426 24488
rect 1472 24442 1501 24488
rect 1001 24335 1030 24381
rect 1076 24335 1089 24381
rect 1001 24274 1089 24335
rect 1001 24228 1030 24274
rect 1076 24228 1089 24274
rect 1001 24167 1089 24228
rect 1001 24121 1030 24167
rect 1076 24121 1089 24167
rect 1001 24060 1089 24121
rect 1001 24014 1030 24060
rect 1076 24014 1089 24060
rect 1001 24001 1089 24014
rect 1413 24381 1501 24442
rect 1413 24335 1426 24381
rect 1472 24335 1501 24381
rect 1413 24274 1501 24335
rect 1413 24228 1426 24274
rect 1472 24228 1501 24274
rect 1413 24167 1501 24228
rect 1413 24121 1426 24167
rect 1472 24121 1501 24167
rect 1413 24060 1501 24121
rect 1413 24014 1426 24060
rect 1472 24014 1501 24060
rect 1413 24001 1501 24014
rect 1621 25350 1709 25363
rect 1621 25304 1650 25350
rect 1696 25304 1709 25350
rect 1621 25242 1709 25304
rect 1621 25196 1650 25242
rect 1696 25196 1709 25242
rect 1621 25134 1709 25196
rect 1621 25088 1650 25134
rect 1696 25088 1709 25134
rect 1621 25026 1709 25088
rect 1621 24980 1650 25026
rect 1696 24980 1709 25026
rect 1621 24918 1709 24980
rect 1621 24872 1650 24918
rect 1696 24872 1709 24918
rect 1621 24810 1709 24872
rect 1621 24764 1650 24810
rect 1696 24764 1709 24810
rect 1621 24702 1709 24764
rect 1621 24656 1650 24702
rect 1696 24656 1709 24702
rect 1621 24595 1709 24656
rect 1621 24549 1650 24595
rect 1696 24549 1709 24595
rect 1621 24488 1709 24549
rect 1621 24442 1650 24488
rect 1696 24442 1709 24488
rect 1621 24381 1709 24442
rect 1621 24335 1650 24381
rect 1696 24335 1709 24381
rect 1621 24274 1709 24335
rect 1621 24228 1650 24274
rect 1696 24228 1709 24274
rect 1621 24167 1709 24228
rect 1621 24121 1650 24167
rect 1696 24121 1709 24167
rect 1621 24060 1709 24121
rect 1621 24014 1650 24060
rect 1696 24014 1709 24060
rect 1621 24001 1709 24014
rect 2032 25350 2120 25363
rect 2032 25304 2045 25350
rect 2091 25304 2120 25350
rect 2032 25242 2120 25304
rect 2032 25196 2045 25242
rect 2091 25196 2120 25242
rect 2032 25134 2120 25196
rect 2032 25088 2045 25134
rect 2091 25088 2120 25134
rect 2032 25026 2120 25088
rect 2032 24980 2045 25026
rect 2091 24980 2120 25026
rect 2032 24918 2120 24980
rect 2032 24872 2045 24918
rect 2091 24872 2120 24918
rect 2032 24810 2120 24872
rect 2032 24764 2045 24810
rect 2091 24764 2120 24810
rect 2032 24702 2120 24764
rect 2032 24656 2045 24702
rect 2091 24656 2120 24702
rect 2032 24595 2120 24656
rect 2032 24549 2045 24595
rect 2091 24549 2120 24595
rect 2032 24488 2120 24549
rect 2032 24442 2045 24488
rect 2091 24442 2120 24488
rect 2032 24381 2120 24442
rect 2032 24335 2045 24381
rect 2091 24335 2120 24381
rect 2032 24274 2120 24335
rect 2032 24228 2045 24274
rect 2091 24228 2120 24274
rect 2032 24167 2120 24228
rect 2032 24121 2045 24167
rect 2091 24121 2120 24167
rect 2032 24060 2120 24121
rect 2032 24014 2045 24060
rect 2091 24014 2120 24060
rect 2032 24001 2120 24014
rect 2240 25350 2328 25363
rect 2240 25304 2269 25350
rect 2315 25304 2328 25350
rect 2240 25242 2328 25304
rect 2240 25196 2269 25242
rect 2315 25196 2328 25242
rect 2240 25134 2328 25196
rect 2240 25088 2269 25134
rect 2315 25088 2328 25134
rect 2240 25026 2328 25088
rect 2240 24980 2269 25026
rect 2315 24980 2328 25026
rect 2240 24918 2328 24980
rect 2240 24872 2269 24918
rect 2315 24872 2328 24918
rect 2240 24810 2328 24872
rect 2240 24764 2269 24810
rect 2315 24764 2328 24810
rect 2240 24702 2328 24764
rect 2240 24656 2269 24702
rect 2315 24656 2328 24702
rect 2652 25350 2740 25363
rect 2652 25304 2665 25350
rect 2711 25304 2740 25350
rect 2652 25242 2740 25304
rect 2652 25196 2665 25242
rect 2711 25196 2740 25242
rect 2652 25134 2740 25196
rect 2652 25088 2665 25134
rect 2711 25088 2740 25134
rect 2652 25026 2740 25088
rect 2652 24980 2665 25026
rect 2711 24980 2740 25026
rect 2652 24918 2740 24980
rect 2652 24872 2665 24918
rect 2711 24872 2740 24918
rect 2652 24810 2740 24872
rect 2652 24764 2665 24810
rect 2711 24764 2740 24810
rect 2652 24702 2740 24764
rect 2240 24595 2328 24656
rect 2240 24549 2269 24595
rect 2315 24549 2328 24595
rect 2240 24488 2328 24549
rect 2240 24442 2269 24488
rect 2315 24442 2328 24488
rect 2240 24381 2328 24442
rect 2652 24656 2665 24702
rect 2711 24656 2740 24702
rect 2652 24595 2740 24656
rect 2652 24549 2665 24595
rect 2711 24549 2740 24595
rect 2652 24488 2740 24549
rect 2652 24442 2665 24488
rect 2711 24442 2740 24488
rect 2240 24335 2269 24381
rect 2315 24335 2328 24381
rect 2240 24274 2328 24335
rect 2240 24228 2269 24274
rect 2315 24228 2328 24274
rect 2240 24167 2328 24228
rect 2240 24121 2269 24167
rect 2315 24121 2328 24167
rect 2240 24060 2328 24121
rect 2240 24014 2269 24060
rect 2315 24014 2328 24060
rect 2240 24001 2328 24014
rect 2652 24381 2740 24442
rect 2652 24335 2665 24381
rect 2711 24335 2740 24381
rect 2652 24274 2740 24335
rect 2652 24228 2665 24274
rect 2711 24228 2740 24274
rect 2652 24167 2740 24228
rect 2652 24121 2665 24167
rect 2711 24121 2740 24167
rect 2652 24060 2740 24121
rect 2652 24014 2665 24060
rect 2711 24014 2740 24060
rect 2652 24001 2740 24014
rect 2860 25350 2948 25363
rect 2860 25304 2889 25350
rect 2935 25304 2948 25350
rect 2860 25242 2948 25304
rect 2860 25196 2889 25242
rect 2935 25196 2948 25242
rect 2860 25134 2948 25196
rect 2860 25088 2889 25134
rect 2935 25088 2948 25134
rect 2860 25026 2948 25088
rect 2860 24980 2889 25026
rect 2935 24980 2948 25026
rect 2860 24918 2948 24980
rect 2860 24872 2889 24918
rect 2935 24872 2948 24918
rect 2860 24810 2948 24872
rect 2860 24764 2889 24810
rect 2935 24764 2948 24810
rect 2860 24702 2948 24764
rect 2860 24656 2889 24702
rect 2935 24656 2948 24702
rect 2860 24595 2948 24656
rect 2860 24549 2889 24595
rect 2935 24549 2948 24595
rect 2860 24488 2948 24549
rect 2860 24442 2889 24488
rect 2935 24442 2948 24488
rect 2860 24381 2948 24442
rect 2860 24335 2889 24381
rect 2935 24335 2948 24381
rect 2860 24274 2948 24335
rect 2860 24228 2889 24274
rect 2935 24228 2948 24274
rect 2860 24167 2948 24228
rect 2860 24121 2889 24167
rect 2935 24121 2948 24167
rect 2860 24060 2948 24121
rect 2860 24014 2889 24060
rect 2935 24014 2948 24060
rect 2860 24001 2948 24014
rect 3270 25350 3358 25363
rect 3270 25304 3283 25350
rect 3329 25304 3358 25350
rect 3270 25242 3358 25304
rect 3270 25196 3283 25242
rect 3329 25196 3358 25242
rect 3270 25134 3358 25196
rect 3270 25088 3283 25134
rect 3329 25088 3358 25134
rect 3270 25026 3358 25088
rect 3270 24980 3283 25026
rect 3329 24980 3358 25026
rect 3270 24918 3358 24980
rect 3270 24872 3283 24918
rect 3329 24872 3358 24918
rect 3270 24810 3358 24872
rect 3270 24764 3283 24810
rect 3329 24764 3358 24810
rect 3270 24702 3358 24764
rect 3270 24656 3283 24702
rect 3329 24656 3358 24702
rect 3270 24595 3358 24656
rect 3270 24549 3283 24595
rect 3329 24549 3358 24595
rect 3270 24488 3358 24549
rect 3270 24442 3283 24488
rect 3329 24442 3358 24488
rect 3270 24381 3358 24442
rect 3270 24335 3283 24381
rect 3329 24335 3358 24381
rect 3270 24274 3358 24335
rect 3270 24228 3283 24274
rect 3329 24228 3358 24274
rect 3270 24167 3358 24228
rect 3270 24121 3283 24167
rect 3329 24121 3358 24167
rect 3270 24060 3358 24121
rect 3270 24014 3283 24060
rect 3329 24014 3358 24060
rect 3270 24001 3358 24014
rect 3478 25350 3566 25363
rect 3478 25304 3507 25350
rect 3553 25304 3566 25350
rect 3478 25242 3566 25304
rect 3478 25196 3507 25242
rect 3553 25196 3566 25242
rect 3478 25134 3566 25196
rect 3478 25088 3507 25134
rect 3553 25088 3566 25134
rect 3478 25026 3566 25088
rect 3478 24980 3507 25026
rect 3553 24980 3566 25026
rect 3478 24918 3566 24980
rect 3478 24872 3507 24918
rect 3553 24872 3566 24918
rect 3478 24810 3566 24872
rect 3478 24764 3507 24810
rect 3553 24764 3566 24810
rect 3478 24702 3566 24764
rect 3478 24656 3507 24702
rect 3553 24656 3566 24702
rect 3890 25350 3978 25363
rect 3890 25304 3903 25350
rect 3949 25304 3978 25350
rect 3890 25242 3978 25304
rect 3890 25196 3903 25242
rect 3949 25196 3978 25242
rect 3890 25134 3978 25196
rect 3890 25088 3903 25134
rect 3949 25088 3978 25134
rect 3890 25026 3978 25088
rect 3890 24980 3903 25026
rect 3949 24980 3978 25026
rect 3890 24918 3978 24980
rect 3890 24872 3903 24918
rect 3949 24872 3978 24918
rect 3890 24810 3978 24872
rect 3890 24764 3903 24810
rect 3949 24764 3978 24810
rect 3890 24702 3978 24764
rect 3478 24595 3566 24656
rect 3478 24549 3507 24595
rect 3553 24549 3566 24595
rect 3478 24488 3566 24549
rect 3478 24442 3507 24488
rect 3553 24442 3566 24488
rect 3478 24381 3566 24442
rect 3890 24656 3903 24702
rect 3949 24656 3978 24702
rect 3890 24595 3978 24656
rect 3890 24549 3903 24595
rect 3949 24549 3978 24595
rect 3890 24488 3978 24549
rect 3890 24442 3903 24488
rect 3949 24442 3978 24488
rect 3478 24335 3507 24381
rect 3553 24335 3566 24381
rect 3478 24274 3566 24335
rect 3478 24228 3507 24274
rect 3553 24228 3566 24274
rect 3478 24167 3566 24228
rect 3478 24121 3507 24167
rect 3553 24121 3566 24167
rect 3478 24060 3566 24121
rect 3478 24014 3507 24060
rect 3553 24014 3566 24060
rect 3478 24001 3566 24014
rect 3890 24381 3978 24442
rect 3890 24335 3903 24381
rect 3949 24335 3978 24381
rect 3890 24274 3978 24335
rect 3890 24228 3903 24274
rect 3949 24228 3978 24274
rect 3890 24167 3978 24228
rect 3890 24121 3903 24167
rect 3949 24121 3978 24167
rect 3890 24060 3978 24121
rect 3890 24014 3903 24060
rect 3949 24014 3978 24060
rect 3890 24001 3978 24014
rect 4098 25350 4186 25363
rect 4098 25304 4127 25350
rect 4173 25304 4186 25350
rect 4098 25242 4186 25304
rect 4098 25196 4127 25242
rect 4173 25196 4186 25242
rect 4098 25134 4186 25196
rect 4098 25088 4127 25134
rect 4173 25088 4186 25134
rect 4098 25026 4186 25088
rect 4098 24980 4127 25026
rect 4173 24980 4186 25026
rect 4098 24918 4186 24980
rect 4098 24872 4127 24918
rect 4173 24872 4186 24918
rect 4098 24810 4186 24872
rect 4098 24764 4127 24810
rect 4173 24764 4186 24810
rect 4098 24702 4186 24764
rect 4098 24656 4127 24702
rect 4173 24656 4186 24702
rect 4098 24595 4186 24656
rect 4098 24549 4127 24595
rect 4173 24549 4186 24595
rect 4098 24488 4186 24549
rect 4098 24442 4127 24488
rect 4173 24442 4186 24488
rect 4098 24381 4186 24442
rect 4098 24335 4127 24381
rect 4173 24335 4186 24381
rect 4098 24274 4186 24335
rect 4098 24228 4127 24274
rect 4173 24228 4186 24274
rect 4098 24167 4186 24228
rect 4098 24121 4127 24167
rect 4173 24121 4186 24167
rect 4098 24060 4186 24121
rect 4098 24014 4127 24060
rect 4173 24014 4186 24060
rect 4098 24001 4186 24014
rect 4509 25350 4597 25363
rect 4509 25304 4522 25350
rect 4568 25304 4597 25350
rect 4509 25242 4597 25304
rect 4509 25196 4522 25242
rect 4568 25196 4597 25242
rect 4509 25134 4597 25196
rect 4509 25088 4522 25134
rect 4568 25088 4597 25134
rect 4509 25026 4597 25088
rect 4509 24980 4522 25026
rect 4568 24980 4597 25026
rect 4509 24918 4597 24980
rect 4509 24872 4522 24918
rect 4568 24872 4597 24918
rect 4509 24810 4597 24872
rect 4509 24764 4522 24810
rect 4568 24764 4597 24810
rect 4509 24702 4597 24764
rect 4509 24656 4522 24702
rect 4568 24656 4597 24702
rect 4509 24595 4597 24656
rect 4509 24549 4522 24595
rect 4568 24549 4597 24595
rect 4509 24488 4597 24549
rect 4509 24442 4522 24488
rect 4568 24442 4597 24488
rect 4509 24381 4597 24442
rect 4509 24335 4522 24381
rect 4568 24335 4597 24381
rect 4509 24274 4597 24335
rect 4509 24228 4522 24274
rect 4568 24228 4597 24274
rect 4509 24167 4597 24228
rect 4509 24121 4522 24167
rect 4568 24121 4597 24167
rect 4509 24060 4597 24121
rect 4509 24014 4522 24060
rect 4568 24014 4597 24060
rect 4509 24001 4597 24014
rect 4717 25350 4805 25363
rect 4717 25304 4746 25350
rect 4792 25304 4805 25350
rect 4717 25242 4805 25304
rect 4717 25196 4746 25242
rect 4792 25196 4805 25242
rect 4717 25134 4805 25196
rect 4717 25088 4746 25134
rect 4792 25088 4805 25134
rect 4717 25026 4805 25088
rect 4717 24980 4746 25026
rect 4792 24980 4805 25026
rect 4717 24918 4805 24980
rect 4717 24872 4746 24918
rect 4792 24872 4805 24918
rect 4717 24810 4805 24872
rect 4717 24764 4746 24810
rect 4792 24764 4805 24810
rect 4717 24702 4805 24764
rect 4717 24656 4746 24702
rect 4792 24656 4805 24702
rect 5129 25350 5217 25363
rect 5129 25304 5142 25350
rect 5188 25304 5217 25350
rect 5129 25242 5217 25304
rect 5129 25196 5142 25242
rect 5188 25196 5217 25242
rect 5129 25134 5217 25196
rect 5129 25088 5142 25134
rect 5188 25088 5217 25134
rect 5129 25026 5217 25088
rect 5129 24980 5142 25026
rect 5188 24980 5217 25026
rect 5129 24918 5217 24980
rect 5129 24872 5142 24918
rect 5188 24872 5217 24918
rect 5129 24810 5217 24872
rect 5129 24764 5142 24810
rect 5188 24764 5217 24810
rect 5129 24702 5217 24764
rect 4717 24595 4805 24656
rect 4717 24549 4746 24595
rect 4792 24549 4805 24595
rect 4717 24488 4805 24549
rect 4717 24442 4746 24488
rect 4792 24442 4805 24488
rect 4717 24381 4805 24442
rect 5129 24656 5142 24702
rect 5188 24656 5217 24702
rect 5129 24595 5217 24656
rect 5129 24549 5142 24595
rect 5188 24549 5217 24595
rect 5129 24488 5217 24549
rect 5129 24442 5142 24488
rect 5188 24442 5217 24488
rect 4717 24335 4746 24381
rect 4792 24335 4805 24381
rect 4717 24274 4805 24335
rect 4717 24228 4746 24274
rect 4792 24228 4805 24274
rect 4717 24167 4805 24228
rect 4717 24121 4746 24167
rect 4792 24121 4805 24167
rect 4717 24060 4805 24121
rect 4717 24014 4746 24060
rect 4792 24014 4805 24060
rect 4717 24001 4805 24014
rect 5129 24381 5217 24442
rect 5129 24335 5142 24381
rect 5188 24335 5217 24381
rect 5129 24274 5217 24335
rect 5129 24228 5142 24274
rect 5188 24228 5217 24274
rect 5129 24167 5217 24228
rect 5129 24121 5142 24167
rect 5188 24121 5217 24167
rect 5129 24060 5217 24121
rect 5129 24014 5142 24060
rect 5188 24014 5217 24060
rect 5129 24001 5217 24014
rect 5337 25350 5425 25363
rect 5337 25304 5366 25350
rect 5412 25304 5425 25350
rect 5337 25242 5425 25304
rect 5337 25196 5366 25242
rect 5412 25196 5425 25242
rect 5337 25134 5425 25196
rect 5337 25088 5366 25134
rect 5412 25088 5425 25134
rect 5337 25026 5425 25088
rect 5337 24980 5366 25026
rect 5412 24980 5425 25026
rect 5337 24918 5425 24980
rect 5337 24872 5366 24918
rect 5412 24872 5425 24918
rect 5337 24810 5425 24872
rect 5337 24764 5366 24810
rect 5412 24764 5425 24810
rect 5337 24702 5425 24764
rect 5337 24656 5366 24702
rect 5412 24656 5425 24702
rect 5337 24595 5425 24656
rect 5337 24549 5366 24595
rect 5412 24549 5425 24595
rect 5337 24488 5425 24549
rect 5337 24442 5366 24488
rect 5412 24442 5425 24488
rect 5337 24381 5425 24442
rect 5337 24335 5366 24381
rect 5412 24335 5425 24381
rect 5337 24274 5425 24335
rect 5337 24228 5366 24274
rect 5412 24228 5425 24274
rect 5337 24167 5425 24228
rect 5337 24121 5366 24167
rect 5412 24121 5425 24167
rect 5337 24060 5425 24121
rect 5337 24014 5366 24060
rect 5412 24014 5425 24060
rect 5337 24001 5425 24014
rect 793 19800 881 19813
rect 793 19754 806 19800
rect 852 19754 881 19800
rect 793 19692 881 19754
rect 793 19646 806 19692
rect 852 19646 881 19692
rect 793 19584 881 19646
rect 793 19538 806 19584
rect 852 19538 881 19584
rect 793 19476 881 19538
rect 793 19430 806 19476
rect 852 19430 881 19476
rect 793 19368 881 19430
rect 793 19322 806 19368
rect 852 19322 881 19368
rect 793 19260 881 19322
rect 793 19214 806 19260
rect 852 19214 881 19260
rect 793 19152 881 19214
rect 793 19106 806 19152
rect 852 19106 881 19152
rect 793 19045 881 19106
rect 793 18999 806 19045
rect 852 18999 881 19045
rect 793 18938 881 18999
rect 793 18892 806 18938
rect 852 18892 881 18938
rect 793 18831 881 18892
rect 793 18785 806 18831
rect 852 18785 881 18831
rect 793 18724 881 18785
rect 793 18678 806 18724
rect 852 18678 881 18724
rect 793 18617 881 18678
rect 793 18571 806 18617
rect 852 18571 881 18617
rect 793 18510 881 18571
rect 793 18464 806 18510
rect 852 18464 881 18510
rect 793 18451 881 18464
rect 1001 19800 1089 19813
rect 1001 19754 1030 19800
rect 1076 19754 1089 19800
rect 1001 19692 1089 19754
rect 1001 19646 1030 19692
rect 1076 19646 1089 19692
rect 1001 19584 1089 19646
rect 1001 19538 1030 19584
rect 1076 19538 1089 19584
rect 1001 19476 1089 19538
rect 1001 19430 1030 19476
rect 1076 19430 1089 19476
rect 1001 19368 1089 19430
rect 1001 19322 1030 19368
rect 1076 19322 1089 19368
rect 1001 19260 1089 19322
rect 1001 19214 1030 19260
rect 1076 19214 1089 19260
rect 1001 19152 1089 19214
rect 1001 19106 1030 19152
rect 1076 19106 1089 19152
rect 1001 19045 1089 19106
rect 1001 18999 1030 19045
rect 1076 18999 1089 19045
rect 1001 18938 1089 18999
rect 1001 18892 1030 18938
rect 1076 18892 1089 18938
rect 1001 18831 1089 18892
rect 1001 18785 1030 18831
rect 1076 18785 1089 18831
rect 1001 18724 1089 18785
rect 1001 18678 1030 18724
rect 1076 18678 1089 18724
rect 1001 18617 1089 18678
rect 1001 18571 1030 18617
rect 1076 18571 1089 18617
rect 1001 18510 1089 18571
rect 1001 18464 1030 18510
rect 1076 18464 1089 18510
rect 1001 18451 1089 18464
rect 1413 19800 1501 19813
rect 1413 19754 1426 19800
rect 1472 19754 1501 19800
rect 1413 19692 1501 19754
rect 1413 19646 1426 19692
rect 1472 19646 1501 19692
rect 1413 19584 1501 19646
rect 1413 19538 1426 19584
rect 1472 19538 1501 19584
rect 1413 19476 1501 19538
rect 1413 19430 1426 19476
rect 1472 19430 1501 19476
rect 1413 19368 1501 19430
rect 1413 19322 1426 19368
rect 1472 19322 1501 19368
rect 1413 19260 1501 19322
rect 1413 19214 1426 19260
rect 1472 19214 1501 19260
rect 1413 19152 1501 19214
rect 1413 19106 1426 19152
rect 1472 19106 1501 19152
rect 1413 19045 1501 19106
rect 1413 18999 1426 19045
rect 1472 18999 1501 19045
rect 1413 18938 1501 18999
rect 1413 18892 1426 18938
rect 1472 18892 1501 18938
rect 1413 18831 1501 18892
rect 1413 18785 1426 18831
rect 1472 18785 1501 18831
rect 1413 18724 1501 18785
rect 1413 18678 1426 18724
rect 1472 18678 1501 18724
rect 1413 18617 1501 18678
rect 1413 18571 1426 18617
rect 1472 18571 1501 18617
rect 1413 18510 1501 18571
rect 1413 18464 1426 18510
rect 1472 18464 1501 18510
rect 1413 18451 1501 18464
rect 1621 19800 1709 19813
rect 1621 19754 1650 19800
rect 1696 19754 1709 19800
rect 1621 19692 1709 19754
rect 1621 19646 1650 19692
rect 1696 19646 1709 19692
rect 1621 19584 1709 19646
rect 1621 19538 1650 19584
rect 1696 19538 1709 19584
rect 1621 19476 1709 19538
rect 1621 19430 1650 19476
rect 1696 19430 1709 19476
rect 1621 19368 1709 19430
rect 1621 19322 1650 19368
rect 1696 19322 1709 19368
rect 1621 19260 1709 19322
rect 1621 19214 1650 19260
rect 1696 19214 1709 19260
rect 1621 19152 1709 19214
rect 1621 19106 1650 19152
rect 1696 19106 1709 19152
rect 1621 19045 1709 19106
rect 1621 18999 1650 19045
rect 1696 18999 1709 19045
rect 1621 18938 1709 18999
rect 1621 18892 1650 18938
rect 1696 18892 1709 18938
rect 1621 18831 1709 18892
rect 1621 18785 1650 18831
rect 1696 18785 1709 18831
rect 1621 18724 1709 18785
rect 1621 18678 1650 18724
rect 1696 18678 1709 18724
rect 1621 18617 1709 18678
rect 1621 18571 1650 18617
rect 1696 18571 1709 18617
rect 1621 18510 1709 18571
rect 1621 18464 1650 18510
rect 1696 18464 1709 18510
rect 1621 18451 1709 18464
rect 2032 19800 2120 19813
rect 2032 19754 2045 19800
rect 2091 19754 2120 19800
rect 2032 19692 2120 19754
rect 2032 19646 2045 19692
rect 2091 19646 2120 19692
rect 2032 19584 2120 19646
rect 2032 19538 2045 19584
rect 2091 19538 2120 19584
rect 2032 19476 2120 19538
rect 2032 19430 2045 19476
rect 2091 19430 2120 19476
rect 2032 19368 2120 19430
rect 2032 19322 2045 19368
rect 2091 19322 2120 19368
rect 2032 19260 2120 19322
rect 2032 19214 2045 19260
rect 2091 19214 2120 19260
rect 2032 19152 2120 19214
rect 2032 19106 2045 19152
rect 2091 19106 2120 19152
rect 2032 19045 2120 19106
rect 2032 18999 2045 19045
rect 2091 18999 2120 19045
rect 2032 18938 2120 18999
rect 2032 18892 2045 18938
rect 2091 18892 2120 18938
rect 2032 18831 2120 18892
rect 2032 18785 2045 18831
rect 2091 18785 2120 18831
rect 2032 18724 2120 18785
rect 2032 18678 2045 18724
rect 2091 18678 2120 18724
rect 2032 18617 2120 18678
rect 2032 18571 2045 18617
rect 2091 18571 2120 18617
rect 2032 18510 2120 18571
rect 2032 18464 2045 18510
rect 2091 18464 2120 18510
rect 2032 18451 2120 18464
rect 2240 19800 2328 19813
rect 2240 19754 2269 19800
rect 2315 19754 2328 19800
rect 2240 19692 2328 19754
rect 2240 19646 2269 19692
rect 2315 19646 2328 19692
rect 2240 19584 2328 19646
rect 2240 19538 2269 19584
rect 2315 19538 2328 19584
rect 2240 19476 2328 19538
rect 2240 19430 2269 19476
rect 2315 19430 2328 19476
rect 2240 19368 2328 19430
rect 2240 19322 2269 19368
rect 2315 19322 2328 19368
rect 2240 19260 2328 19322
rect 2240 19214 2269 19260
rect 2315 19214 2328 19260
rect 2240 19152 2328 19214
rect 2240 19106 2269 19152
rect 2315 19106 2328 19152
rect 2240 19045 2328 19106
rect 2240 18999 2269 19045
rect 2315 18999 2328 19045
rect 2240 18938 2328 18999
rect 2240 18892 2269 18938
rect 2315 18892 2328 18938
rect 2240 18831 2328 18892
rect 2240 18785 2269 18831
rect 2315 18785 2328 18831
rect 2240 18724 2328 18785
rect 2240 18678 2269 18724
rect 2315 18678 2328 18724
rect 2240 18617 2328 18678
rect 2240 18571 2269 18617
rect 2315 18571 2328 18617
rect 2240 18510 2328 18571
rect 2240 18464 2269 18510
rect 2315 18464 2328 18510
rect 2240 18451 2328 18464
rect 2652 19800 2740 19813
rect 2652 19754 2665 19800
rect 2711 19754 2740 19800
rect 2652 19692 2740 19754
rect 2652 19646 2665 19692
rect 2711 19646 2740 19692
rect 2652 19584 2740 19646
rect 2652 19538 2665 19584
rect 2711 19538 2740 19584
rect 2652 19476 2740 19538
rect 2652 19430 2665 19476
rect 2711 19430 2740 19476
rect 2652 19368 2740 19430
rect 2652 19322 2665 19368
rect 2711 19322 2740 19368
rect 2652 19260 2740 19322
rect 2652 19214 2665 19260
rect 2711 19214 2740 19260
rect 2652 19152 2740 19214
rect 2652 19106 2665 19152
rect 2711 19106 2740 19152
rect 2652 19045 2740 19106
rect 2652 18999 2665 19045
rect 2711 18999 2740 19045
rect 2652 18938 2740 18999
rect 2652 18892 2665 18938
rect 2711 18892 2740 18938
rect 2652 18831 2740 18892
rect 2652 18785 2665 18831
rect 2711 18785 2740 18831
rect 2652 18724 2740 18785
rect 2652 18678 2665 18724
rect 2711 18678 2740 18724
rect 2652 18617 2740 18678
rect 2652 18571 2665 18617
rect 2711 18571 2740 18617
rect 2652 18510 2740 18571
rect 2652 18464 2665 18510
rect 2711 18464 2740 18510
rect 2652 18451 2740 18464
rect 2860 19800 2948 19813
rect 2860 19754 2889 19800
rect 2935 19754 2948 19800
rect 2860 19692 2948 19754
rect 2860 19646 2889 19692
rect 2935 19646 2948 19692
rect 2860 19584 2948 19646
rect 2860 19538 2889 19584
rect 2935 19538 2948 19584
rect 2860 19476 2948 19538
rect 2860 19430 2889 19476
rect 2935 19430 2948 19476
rect 2860 19368 2948 19430
rect 2860 19322 2889 19368
rect 2935 19322 2948 19368
rect 2860 19260 2948 19322
rect 2860 19214 2889 19260
rect 2935 19214 2948 19260
rect 2860 19152 2948 19214
rect 2860 19106 2889 19152
rect 2935 19106 2948 19152
rect 2860 19045 2948 19106
rect 2860 18999 2889 19045
rect 2935 18999 2948 19045
rect 2860 18938 2948 18999
rect 2860 18892 2889 18938
rect 2935 18892 2948 18938
rect 2860 18831 2948 18892
rect 2860 18785 2889 18831
rect 2935 18785 2948 18831
rect 2860 18724 2948 18785
rect 2860 18678 2889 18724
rect 2935 18678 2948 18724
rect 2860 18617 2948 18678
rect 2860 18571 2889 18617
rect 2935 18571 2948 18617
rect 2860 18510 2948 18571
rect 2860 18464 2889 18510
rect 2935 18464 2948 18510
rect 2860 18451 2948 18464
rect 3270 19800 3358 19813
rect 3270 19754 3283 19800
rect 3329 19754 3358 19800
rect 3270 19692 3358 19754
rect 3270 19646 3283 19692
rect 3329 19646 3358 19692
rect 3270 19584 3358 19646
rect 3270 19538 3283 19584
rect 3329 19538 3358 19584
rect 3270 19476 3358 19538
rect 3270 19430 3283 19476
rect 3329 19430 3358 19476
rect 3270 19368 3358 19430
rect 3270 19322 3283 19368
rect 3329 19322 3358 19368
rect 3270 19260 3358 19322
rect 3270 19214 3283 19260
rect 3329 19214 3358 19260
rect 3270 19152 3358 19214
rect 3270 19106 3283 19152
rect 3329 19106 3358 19152
rect 3270 19045 3358 19106
rect 3270 18999 3283 19045
rect 3329 18999 3358 19045
rect 3270 18938 3358 18999
rect 3270 18892 3283 18938
rect 3329 18892 3358 18938
rect 3270 18831 3358 18892
rect 3270 18785 3283 18831
rect 3329 18785 3358 18831
rect 3270 18724 3358 18785
rect 3270 18678 3283 18724
rect 3329 18678 3358 18724
rect 3270 18617 3358 18678
rect 3270 18571 3283 18617
rect 3329 18571 3358 18617
rect 3270 18510 3358 18571
rect 3270 18464 3283 18510
rect 3329 18464 3358 18510
rect 3270 18451 3358 18464
rect 3478 19800 3566 19813
rect 3478 19754 3507 19800
rect 3553 19754 3566 19800
rect 3478 19692 3566 19754
rect 3478 19646 3507 19692
rect 3553 19646 3566 19692
rect 3478 19584 3566 19646
rect 3478 19538 3507 19584
rect 3553 19538 3566 19584
rect 3478 19476 3566 19538
rect 3478 19430 3507 19476
rect 3553 19430 3566 19476
rect 3478 19368 3566 19430
rect 3478 19322 3507 19368
rect 3553 19322 3566 19368
rect 3478 19260 3566 19322
rect 3478 19214 3507 19260
rect 3553 19214 3566 19260
rect 3478 19152 3566 19214
rect 3478 19106 3507 19152
rect 3553 19106 3566 19152
rect 3478 19045 3566 19106
rect 3478 18999 3507 19045
rect 3553 18999 3566 19045
rect 3478 18938 3566 18999
rect 3478 18892 3507 18938
rect 3553 18892 3566 18938
rect 3478 18831 3566 18892
rect 3478 18785 3507 18831
rect 3553 18785 3566 18831
rect 3478 18724 3566 18785
rect 3478 18678 3507 18724
rect 3553 18678 3566 18724
rect 3478 18617 3566 18678
rect 3478 18571 3507 18617
rect 3553 18571 3566 18617
rect 3478 18510 3566 18571
rect 3478 18464 3507 18510
rect 3553 18464 3566 18510
rect 3478 18451 3566 18464
rect 3890 19800 3978 19813
rect 3890 19754 3903 19800
rect 3949 19754 3978 19800
rect 3890 19692 3978 19754
rect 3890 19646 3903 19692
rect 3949 19646 3978 19692
rect 3890 19584 3978 19646
rect 3890 19538 3903 19584
rect 3949 19538 3978 19584
rect 3890 19476 3978 19538
rect 3890 19430 3903 19476
rect 3949 19430 3978 19476
rect 3890 19368 3978 19430
rect 3890 19322 3903 19368
rect 3949 19322 3978 19368
rect 3890 19260 3978 19322
rect 3890 19214 3903 19260
rect 3949 19214 3978 19260
rect 3890 19152 3978 19214
rect 3890 19106 3903 19152
rect 3949 19106 3978 19152
rect 3890 19045 3978 19106
rect 3890 18999 3903 19045
rect 3949 18999 3978 19045
rect 3890 18938 3978 18999
rect 3890 18892 3903 18938
rect 3949 18892 3978 18938
rect 3890 18831 3978 18892
rect 3890 18785 3903 18831
rect 3949 18785 3978 18831
rect 3890 18724 3978 18785
rect 3890 18678 3903 18724
rect 3949 18678 3978 18724
rect 3890 18617 3978 18678
rect 3890 18571 3903 18617
rect 3949 18571 3978 18617
rect 3890 18510 3978 18571
rect 3890 18464 3903 18510
rect 3949 18464 3978 18510
rect 3890 18451 3978 18464
rect 4098 19800 4186 19813
rect 4098 19754 4127 19800
rect 4173 19754 4186 19800
rect 4098 19692 4186 19754
rect 4098 19646 4127 19692
rect 4173 19646 4186 19692
rect 4098 19584 4186 19646
rect 4098 19538 4127 19584
rect 4173 19538 4186 19584
rect 4098 19476 4186 19538
rect 4098 19430 4127 19476
rect 4173 19430 4186 19476
rect 4098 19368 4186 19430
rect 4098 19322 4127 19368
rect 4173 19322 4186 19368
rect 4098 19260 4186 19322
rect 4098 19214 4127 19260
rect 4173 19214 4186 19260
rect 4098 19152 4186 19214
rect 4098 19106 4127 19152
rect 4173 19106 4186 19152
rect 4098 19045 4186 19106
rect 4098 18999 4127 19045
rect 4173 18999 4186 19045
rect 4098 18938 4186 18999
rect 4098 18892 4127 18938
rect 4173 18892 4186 18938
rect 4098 18831 4186 18892
rect 4098 18785 4127 18831
rect 4173 18785 4186 18831
rect 4098 18724 4186 18785
rect 4098 18678 4127 18724
rect 4173 18678 4186 18724
rect 4098 18617 4186 18678
rect 4098 18571 4127 18617
rect 4173 18571 4186 18617
rect 4098 18510 4186 18571
rect 4098 18464 4127 18510
rect 4173 18464 4186 18510
rect 4098 18451 4186 18464
rect 4509 19800 4597 19813
rect 4509 19754 4522 19800
rect 4568 19754 4597 19800
rect 4509 19692 4597 19754
rect 4509 19646 4522 19692
rect 4568 19646 4597 19692
rect 4509 19584 4597 19646
rect 4509 19538 4522 19584
rect 4568 19538 4597 19584
rect 4509 19476 4597 19538
rect 4509 19430 4522 19476
rect 4568 19430 4597 19476
rect 4509 19368 4597 19430
rect 4509 19322 4522 19368
rect 4568 19322 4597 19368
rect 4509 19260 4597 19322
rect 4509 19214 4522 19260
rect 4568 19214 4597 19260
rect 4509 19152 4597 19214
rect 4509 19106 4522 19152
rect 4568 19106 4597 19152
rect 4509 19045 4597 19106
rect 4509 18999 4522 19045
rect 4568 18999 4597 19045
rect 4509 18938 4597 18999
rect 4509 18892 4522 18938
rect 4568 18892 4597 18938
rect 4509 18831 4597 18892
rect 4509 18785 4522 18831
rect 4568 18785 4597 18831
rect 4509 18724 4597 18785
rect 4509 18678 4522 18724
rect 4568 18678 4597 18724
rect 4509 18617 4597 18678
rect 4509 18571 4522 18617
rect 4568 18571 4597 18617
rect 4509 18510 4597 18571
rect 4509 18464 4522 18510
rect 4568 18464 4597 18510
rect 4509 18451 4597 18464
rect 4717 19800 4805 19813
rect 4717 19754 4746 19800
rect 4792 19754 4805 19800
rect 4717 19692 4805 19754
rect 4717 19646 4746 19692
rect 4792 19646 4805 19692
rect 4717 19584 4805 19646
rect 4717 19538 4746 19584
rect 4792 19538 4805 19584
rect 4717 19476 4805 19538
rect 4717 19430 4746 19476
rect 4792 19430 4805 19476
rect 4717 19368 4805 19430
rect 4717 19322 4746 19368
rect 4792 19322 4805 19368
rect 4717 19260 4805 19322
rect 4717 19214 4746 19260
rect 4792 19214 4805 19260
rect 4717 19152 4805 19214
rect 4717 19106 4746 19152
rect 4792 19106 4805 19152
rect 4717 19045 4805 19106
rect 4717 18999 4746 19045
rect 4792 18999 4805 19045
rect 4717 18938 4805 18999
rect 4717 18892 4746 18938
rect 4792 18892 4805 18938
rect 4717 18831 4805 18892
rect 4717 18785 4746 18831
rect 4792 18785 4805 18831
rect 4717 18724 4805 18785
rect 4717 18678 4746 18724
rect 4792 18678 4805 18724
rect 4717 18617 4805 18678
rect 4717 18571 4746 18617
rect 4792 18571 4805 18617
rect 4717 18510 4805 18571
rect 4717 18464 4746 18510
rect 4792 18464 4805 18510
rect 4717 18451 4805 18464
rect 5129 19800 5217 19813
rect 5129 19754 5142 19800
rect 5188 19754 5217 19800
rect 5129 19692 5217 19754
rect 5129 19646 5142 19692
rect 5188 19646 5217 19692
rect 5129 19584 5217 19646
rect 5129 19538 5142 19584
rect 5188 19538 5217 19584
rect 5129 19476 5217 19538
rect 5129 19430 5142 19476
rect 5188 19430 5217 19476
rect 5129 19368 5217 19430
rect 5129 19322 5142 19368
rect 5188 19322 5217 19368
rect 5129 19260 5217 19322
rect 5129 19214 5142 19260
rect 5188 19214 5217 19260
rect 5129 19152 5217 19214
rect 5129 19106 5142 19152
rect 5188 19106 5217 19152
rect 5129 19045 5217 19106
rect 5129 18999 5142 19045
rect 5188 18999 5217 19045
rect 5129 18938 5217 18999
rect 5129 18892 5142 18938
rect 5188 18892 5217 18938
rect 5129 18831 5217 18892
rect 5129 18785 5142 18831
rect 5188 18785 5217 18831
rect 5129 18724 5217 18785
rect 5129 18678 5142 18724
rect 5188 18678 5217 18724
rect 5129 18617 5217 18678
rect 5129 18571 5142 18617
rect 5188 18571 5217 18617
rect 5129 18510 5217 18571
rect 5129 18464 5142 18510
rect 5188 18464 5217 18510
rect 5129 18451 5217 18464
rect 5337 19800 5425 19813
rect 5337 19754 5366 19800
rect 5412 19754 5425 19800
rect 5337 19692 5425 19754
rect 5337 19646 5366 19692
rect 5412 19646 5425 19692
rect 5337 19584 5425 19646
rect 5337 19538 5366 19584
rect 5412 19538 5425 19584
rect 5337 19476 5425 19538
rect 5337 19430 5366 19476
rect 5412 19430 5425 19476
rect 5337 19368 5425 19430
rect 5337 19322 5366 19368
rect 5412 19322 5425 19368
rect 5337 19260 5425 19322
rect 5337 19214 5366 19260
rect 5412 19214 5425 19260
rect 5337 19152 5425 19214
rect 5337 19106 5366 19152
rect 5412 19106 5425 19152
rect 5337 19045 5425 19106
rect 5337 18999 5366 19045
rect 5412 18999 5425 19045
rect 5337 18938 5425 18999
rect 5337 18892 5366 18938
rect 5412 18892 5425 18938
rect 5337 18831 5425 18892
rect 5337 18785 5366 18831
rect 5412 18785 5425 18831
rect 5337 18724 5425 18785
rect 5337 18678 5366 18724
rect 5412 18678 5425 18724
rect 5337 18617 5425 18678
rect 5337 18571 5366 18617
rect 5412 18571 5425 18617
rect 5337 18510 5425 18571
rect 5337 18464 5366 18510
rect 5412 18464 5425 18510
rect 5337 18451 5425 18464
rect 631 17713 812 17838
rect 631 17667 725 17713
rect 771 17667 812 17713
rect 631 17541 812 17667
rect 932 17713 1064 17838
rect 932 17667 975 17713
rect 1021 17667 1064 17713
rect 932 17541 1064 17667
rect 1184 17713 1318 17838
rect 1184 17667 1228 17713
rect 1274 17667 1318 17713
rect 1184 17541 1318 17667
rect 1438 17713 1570 17838
rect 1438 17667 1481 17713
rect 1527 17667 1570 17713
rect 1438 17541 1570 17667
rect 1690 17713 2051 17838
rect 1690 17667 1731 17713
rect 1777 17667 1964 17713
rect 2010 17667 2051 17713
rect 1690 17541 2051 17667
rect 2171 17713 2303 17838
rect 2171 17667 2214 17713
rect 2260 17667 2303 17713
rect 2171 17541 2303 17667
rect 2423 17713 2557 17838
rect 2423 17667 2467 17713
rect 2513 17667 2557 17713
rect 2423 17541 2557 17667
rect 2677 17713 2809 17838
rect 2677 17667 2720 17713
rect 2766 17667 2809 17713
rect 2677 17541 2809 17667
rect 2929 17713 3289 17838
rect 2929 17667 2970 17713
rect 3016 17667 3202 17713
rect 3248 17667 3289 17713
rect 2929 17541 3289 17667
rect 3409 17713 3541 17838
rect 3409 17667 3452 17713
rect 3498 17667 3541 17713
rect 3409 17541 3541 17667
rect 3661 17713 3795 17838
rect 3661 17667 3705 17713
rect 3751 17667 3795 17713
rect 3661 17541 3795 17667
rect 3915 17713 4047 17838
rect 3915 17667 3958 17713
rect 4004 17667 4047 17713
rect 3915 17541 4047 17667
rect 4167 17713 4528 17838
rect 4167 17667 4208 17713
rect 4254 17667 4441 17713
rect 4487 17667 4528 17713
rect 4167 17541 4528 17667
rect 4648 17713 4780 17838
rect 4648 17667 4691 17713
rect 4737 17667 4780 17713
rect 4648 17541 4780 17667
rect 4900 17713 5034 17838
rect 4900 17667 4944 17713
rect 4990 17667 5034 17713
rect 4900 17541 5034 17667
rect 5154 17713 5285 17838
rect 5154 17667 5197 17713
rect 5243 17667 5285 17713
rect 5154 17541 5285 17667
rect 5405 17713 5587 17838
rect 5405 17667 5447 17713
rect 5493 17667 5587 17713
rect 5405 17541 5587 17667
rect 287 15758 375 15771
rect 287 13062 300 15758
rect 346 13062 375 15758
rect 287 13049 375 13062
rect 495 15758 583 15771
rect 495 13062 524 15758
rect 570 13062 583 15758
rect 1631 15304 1719 15317
rect 1631 15258 1644 15304
rect 1690 15258 1719 15304
rect 1631 15200 1719 15258
rect 810 15065 928 15190
rect 810 15019 853 15065
rect 899 15019 928 15065
rect 810 14893 928 15019
rect 1048 15065 1201 15190
rect 1048 15019 1117 15065
rect 1163 15019 1201 15065
rect 1048 14893 1201 15019
rect 1321 15065 1439 15190
rect 1321 15019 1350 15065
rect 1396 15019 1439 15065
rect 1321 14893 1439 15019
rect 1631 15154 1644 15200
rect 1690 15154 1719 15200
rect 1631 15096 1719 15154
rect 1631 15050 1644 15096
rect 1690 15050 1719 15096
rect 1631 14992 1719 15050
rect 1631 14946 1644 14992
rect 1690 14946 1719 14992
rect 1631 14888 1719 14946
rect 1631 14842 1644 14888
rect 1690 14842 1719 14888
rect 1631 14784 1719 14842
rect 1631 14738 1644 14784
rect 1690 14738 1719 14784
rect 1631 14680 1719 14738
rect 1631 14634 1644 14680
rect 1690 14634 1719 14680
rect 1631 14576 1719 14634
rect 1631 14530 1644 14576
rect 1690 14530 1719 14576
rect 1631 14472 1719 14530
rect 1631 14426 1644 14472
rect 1690 14426 1719 14472
rect 495 13049 583 13062
rect 735 14398 823 14411
rect 735 14352 748 14398
rect 794 14352 823 14398
rect 735 14291 823 14352
rect 735 14245 748 14291
rect 794 14245 823 14291
rect 735 14184 823 14245
rect 735 14138 748 14184
rect 794 14138 823 14184
rect 735 14077 823 14138
rect 735 14031 748 14077
rect 794 14031 823 14077
rect 735 13970 823 14031
rect 735 13924 748 13970
rect 794 13924 823 13970
rect 735 13863 823 13924
rect 735 13817 748 13863
rect 794 13817 823 13863
rect 735 13756 823 13817
rect 735 13710 748 13756
rect 794 13710 823 13756
rect 735 13648 823 13710
rect 735 13602 748 13648
rect 794 13602 823 13648
rect 735 13540 823 13602
rect 735 13494 748 13540
rect 794 13494 823 13540
rect 735 13432 823 13494
rect 735 13386 748 13432
rect 794 13386 823 13432
rect 735 13324 823 13386
rect 735 13278 748 13324
rect 794 13278 823 13324
rect 735 13216 823 13278
rect 735 13170 748 13216
rect 794 13170 823 13216
rect 735 13108 823 13170
rect 735 13062 748 13108
rect 794 13062 823 13108
rect 735 13049 823 13062
rect 943 14398 1031 14411
rect 943 14352 972 14398
rect 1018 14352 1031 14398
rect 943 14291 1031 14352
rect 943 14245 972 14291
rect 1018 14245 1031 14291
rect 943 14184 1031 14245
rect 943 14138 972 14184
rect 1018 14138 1031 14184
rect 943 14077 1031 14138
rect 943 14031 972 14077
rect 1018 14031 1031 14077
rect 943 13970 1031 14031
rect 943 13924 972 13970
rect 1018 13924 1031 13970
rect 943 13863 1031 13924
rect 943 13817 972 13863
rect 1018 13817 1031 13863
rect 943 13756 1031 13817
rect 943 13710 972 13756
rect 1018 13710 1031 13756
rect 943 13648 1031 13710
rect 943 13602 972 13648
rect 1018 13602 1031 13648
rect 943 13540 1031 13602
rect 943 13494 972 13540
rect 1018 13494 1031 13540
rect 943 13432 1031 13494
rect 943 13386 972 13432
rect 1018 13386 1031 13432
rect 943 13324 1031 13386
rect 943 13278 972 13324
rect 1018 13278 1031 13324
rect 943 13216 1031 13278
rect 943 13170 972 13216
rect 1018 13170 1031 13216
rect 943 13108 1031 13170
rect 943 13062 972 13108
rect 1018 13062 1031 13108
rect 943 13049 1031 13062
rect 1183 14398 1271 14411
rect 1183 14352 1196 14398
rect 1242 14352 1271 14398
rect 1183 14291 1271 14352
rect 1183 14245 1196 14291
rect 1242 14245 1271 14291
rect 1183 14184 1271 14245
rect 1183 14138 1196 14184
rect 1242 14138 1271 14184
rect 1183 14077 1271 14138
rect 1183 14031 1196 14077
rect 1242 14031 1271 14077
rect 1183 13970 1271 14031
rect 1183 13924 1196 13970
rect 1242 13924 1271 13970
rect 1183 13863 1271 13924
rect 1183 13817 1196 13863
rect 1242 13817 1271 13863
rect 1183 13756 1271 13817
rect 1183 13710 1196 13756
rect 1242 13710 1271 13756
rect 1183 13648 1271 13710
rect 1183 13602 1196 13648
rect 1242 13602 1271 13648
rect 1183 13540 1271 13602
rect 1183 13494 1196 13540
rect 1242 13494 1271 13540
rect 1183 13432 1271 13494
rect 1183 13386 1196 13432
rect 1242 13386 1271 13432
rect 1183 13324 1271 13386
rect 1183 13278 1196 13324
rect 1242 13278 1271 13324
rect 1183 13216 1271 13278
rect 1183 13170 1196 13216
rect 1242 13170 1271 13216
rect 1183 13108 1271 13170
rect 1183 13062 1196 13108
rect 1242 13062 1271 13108
rect 1183 13049 1271 13062
rect 1391 14398 1479 14411
rect 1391 14352 1420 14398
rect 1466 14352 1479 14398
rect 1391 14291 1479 14352
rect 1391 14245 1420 14291
rect 1466 14245 1479 14291
rect 1391 14184 1479 14245
rect 1391 14138 1420 14184
rect 1466 14138 1479 14184
rect 1391 14077 1479 14138
rect 1391 14031 1420 14077
rect 1466 14031 1479 14077
rect 1391 13970 1479 14031
rect 1391 13924 1420 13970
rect 1466 13924 1479 13970
rect 1391 13863 1479 13924
rect 1391 13817 1420 13863
rect 1466 13817 1479 13863
rect 1391 13756 1479 13817
rect 1391 13710 1420 13756
rect 1466 13710 1479 13756
rect 1391 13648 1479 13710
rect 1391 13602 1420 13648
rect 1466 13602 1479 13648
rect 1391 13540 1479 13602
rect 1391 13494 1420 13540
rect 1466 13494 1479 13540
rect 1391 13432 1479 13494
rect 1391 13386 1420 13432
rect 1466 13386 1479 13432
rect 1391 13324 1479 13386
rect 1391 13278 1420 13324
rect 1466 13278 1479 13324
rect 1391 13216 1479 13278
rect 1391 13170 1420 13216
rect 1466 13170 1479 13216
rect 1391 13108 1479 13170
rect 1391 13062 1420 13108
rect 1466 13062 1479 13108
rect 1391 13049 1479 13062
rect 1631 14368 1719 14426
rect 1631 14322 1644 14368
rect 1690 14322 1719 14368
rect 1631 14263 1719 14322
rect 1631 14217 1644 14263
rect 1690 14217 1719 14263
rect 1631 14158 1719 14217
rect 1631 14112 1644 14158
rect 1690 14112 1719 14158
rect 1631 14053 1719 14112
rect 1631 14007 1644 14053
rect 1690 14007 1719 14053
rect 1631 13948 1719 14007
rect 1631 13902 1644 13948
rect 1690 13902 1719 13948
rect 1631 13843 1719 13902
rect 1631 13797 1644 13843
rect 1690 13797 1719 13843
rect 1631 13738 1719 13797
rect 1631 13692 1644 13738
rect 1690 13692 1719 13738
rect 1631 13633 1719 13692
rect 1631 13587 1644 13633
rect 1690 13587 1719 13633
rect 1631 13528 1719 13587
rect 1631 13482 1644 13528
rect 1690 13482 1719 13528
rect 1631 13423 1719 13482
rect 1631 13377 1644 13423
rect 1690 13377 1719 13423
rect 1631 13318 1719 13377
rect 1631 13272 1644 13318
rect 1690 13272 1719 13318
rect 1631 13213 1719 13272
rect 1631 13167 1644 13213
rect 1690 13167 1719 13213
rect 1631 13108 1719 13167
rect 1631 13062 1644 13108
rect 1690 13062 1719 13108
rect 1631 13049 1719 13062
rect 1839 15304 1927 15317
rect 1839 15258 1868 15304
rect 1914 15258 1927 15304
rect 1839 15200 1927 15258
rect 1839 15154 1868 15200
rect 1914 15154 1927 15200
rect 1839 15096 1927 15154
rect 1839 15050 1868 15096
rect 1914 15050 1927 15096
rect 1839 14992 1927 15050
rect 1839 14946 1868 14992
rect 1914 14946 1927 14992
rect 1839 14888 1927 14946
rect 1839 14842 1868 14888
rect 1914 14842 1927 14888
rect 1839 14784 1927 14842
rect 1839 14738 1868 14784
rect 1914 14738 1927 14784
rect 1839 14680 1927 14738
rect 1839 14634 1868 14680
rect 1914 14634 1927 14680
rect 1839 14576 1927 14634
rect 1839 14530 1868 14576
rect 1914 14530 1927 14576
rect 1839 14472 1927 14530
rect 1839 14426 1868 14472
rect 1914 14426 1927 14472
rect 1839 14368 1927 14426
rect 1839 14322 1868 14368
rect 1914 14322 1927 14368
rect 1839 14263 1927 14322
rect 1839 14217 1868 14263
rect 1914 14217 1927 14263
rect 1839 14158 1927 14217
rect 1839 14112 1868 14158
rect 1914 14112 1927 14158
rect 1839 14053 1927 14112
rect 1839 14007 1868 14053
rect 1914 14007 1927 14053
rect 1839 13948 1927 14007
rect 1839 13902 1868 13948
rect 1914 13902 1927 13948
rect 1839 13843 1927 13902
rect 1839 13797 1868 13843
rect 1914 13797 1927 13843
rect 1839 13738 1927 13797
rect 1839 13692 1868 13738
rect 1914 13692 1927 13738
rect 1839 13633 1927 13692
rect 1839 13587 1868 13633
rect 1914 13587 1927 13633
rect 1839 13528 1927 13587
rect 1839 13482 1868 13528
rect 1914 13482 1927 13528
rect 1839 13423 1927 13482
rect 1839 13377 1868 13423
rect 1914 13377 1927 13423
rect 1839 13318 1927 13377
rect 1839 13272 1868 13318
rect 1914 13272 1927 13318
rect 1839 13213 1927 13272
rect 1839 13167 1868 13213
rect 1914 13167 1927 13213
rect 1839 13108 1927 13167
rect 1839 13062 1868 13108
rect 1914 13062 1927 13108
rect 1839 13049 1927 13062
rect 1616 9420 1704 9433
rect 1616 9374 1629 9420
rect 1675 9374 1704 9420
rect 1616 9264 1704 9374
rect 788 9227 876 9240
rect 788 9181 801 9227
rect 847 9181 876 9227
rect 788 9071 876 9181
rect 788 9025 801 9071
rect 847 9025 876 9071
rect 788 9012 876 9025
rect 996 9227 1100 9240
rect 996 9181 1025 9227
rect 1071 9181 1100 9227
rect 996 9071 1100 9181
rect 996 9025 1025 9071
rect 1071 9025 1100 9071
rect 996 9012 1100 9025
rect 1220 9227 1308 9240
rect 1220 9181 1249 9227
rect 1295 9181 1308 9227
rect 1616 9218 1629 9264
rect 1675 9218 1704 9264
rect 1616 9205 1704 9218
rect 1824 9420 1928 9433
rect 1824 9374 1853 9420
rect 1899 9374 1928 9420
rect 1824 9264 1928 9374
rect 1824 9218 1853 9264
rect 1899 9218 1928 9264
rect 1824 9205 1928 9218
rect 2048 9420 2136 9433
rect 2048 9374 2077 9420
rect 2123 9374 2136 9420
rect 2048 9264 2136 9374
rect 2048 9218 2077 9264
rect 2123 9218 2136 9264
rect 2048 9205 2136 9218
rect 2468 9245 2556 9258
rect 1220 9071 1308 9181
rect 2468 9199 2481 9245
rect 2527 9199 2556 9245
rect 2468 9138 2556 9199
rect 1220 9025 1249 9071
rect 1295 9025 1308 9071
rect 2468 9092 2481 9138
rect 2527 9092 2556 9138
rect 1220 9012 1308 9025
rect 2468 9031 2556 9092
rect 2468 8985 2481 9031
rect 2527 8985 2556 9031
rect 2468 8924 2556 8985
rect 2468 8878 2481 8924
rect 2527 8878 2556 8924
rect 2468 8817 2556 8878
rect 2468 8771 2481 8817
rect 2527 8771 2556 8817
rect 1616 8705 1704 8718
rect 1616 8659 1629 8705
rect 1675 8659 1704 8705
rect 788 8623 876 8636
rect 788 8577 801 8623
rect 847 8577 876 8623
rect 788 8503 876 8577
rect 788 8457 801 8503
rect 847 8457 876 8503
rect 788 8444 876 8457
rect 996 8623 1100 8636
rect 996 8577 1025 8623
rect 1071 8577 1100 8623
rect 996 8503 1100 8577
rect 996 8457 1025 8503
rect 1071 8457 1100 8503
rect 996 8444 1100 8457
rect 1220 8623 1308 8636
rect 1220 8577 1249 8623
rect 1295 8577 1308 8623
rect 1220 8503 1308 8577
rect 1616 8585 1704 8659
rect 1616 8539 1629 8585
rect 1675 8539 1704 8585
rect 1616 8526 1704 8539
rect 1824 8705 1928 8718
rect 1824 8659 1853 8705
rect 1899 8659 1928 8705
rect 1824 8585 1928 8659
rect 1824 8539 1853 8585
rect 1899 8539 1928 8585
rect 1824 8526 1928 8539
rect 2048 8705 2136 8718
rect 2048 8659 2077 8705
rect 2123 8659 2136 8705
rect 2048 8585 2136 8659
rect 2048 8539 2077 8585
rect 2123 8539 2136 8585
rect 2048 8526 2136 8539
rect 2468 8710 2556 8771
rect 2468 8664 2481 8710
rect 2527 8664 2556 8710
rect 2468 8603 2556 8664
rect 2468 8557 2481 8603
rect 2527 8557 2556 8603
rect 1220 8457 1249 8503
rect 1295 8457 1308 8503
rect 1220 8444 1308 8457
rect 2468 8495 2556 8557
rect 2468 8449 2481 8495
rect 2527 8449 2556 8495
rect 2468 8387 2556 8449
rect 2468 8341 2481 8387
rect 2527 8341 2556 8387
rect 2468 8279 2556 8341
rect 2468 8233 2481 8279
rect 2527 8233 2556 8279
rect 2468 8171 2556 8233
rect 2468 8125 2481 8171
rect 2527 8125 2556 8171
rect 2468 8063 2556 8125
rect 2468 8017 2481 8063
rect 2527 8017 2556 8063
rect 2468 7955 2556 8017
rect 2468 7909 2481 7955
rect 2527 7909 2556 7955
rect 2468 7896 2556 7909
rect 2676 9245 2764 9258
rect 2676 9199 2705 9245
rect 2751 9199 2764 9245
rect 2676 9138 2764 9199
rect 2676 9092 2705 9138
rect 2751 9092 2764 9138
rect 2676 9031 2764 9092
rect 2676 8985 2705 9031
rect 2751 8985 2764 9031
rect 2676 8924 2764 8985
rect 2676 8878 2705 8924
rect 2751 8878 2764 8924
rect 2676 8817 2764 8878
rect 2676 8771 2705 8817
rect 2751 8771 2764 8817
rect 2676 8710 2764 8771
rect 2676 8664 2705 8710
rect 2751 8664 2764 8710
rect 2676 8603 2764 8664
rect 2676 8557 2705 8603
rect 2751 8557 2764 8603
rect 2676 8495 2764 8557
rect 2676 8449 2705 8495
rect 2751 8449 2764 8495
rect 2676 8387 2764 8449
rect 2676 8341 2705 8387
rect 2751 8341 2764 8387
rect 2676 8279 2764 8341
rect 2676 8233 2705 8279
rect 2751 8233 2764 8279
rect 2676 8171 2764 8233
rect 2676 8125 2705 8171
rect 2751 8125 2764 8171
rect 2676 8063 2764 8125
rect 2676 8017 2705 8063
rect 2751 8017 2764 8063
rect 2676 7955 2764 8017
rect 2676 7909 2705 7955
rect 2751 7909 2764 7955
rect 2676 7896 2764 7909
<< mvndiffc >>
rect 806 23613 852 23659
rect 806 23505 852 23551
rect 806 23397 852 23443
rect 806 23289 852 23335
rect 806 23181 852 23227
rect 806 23073 852 23119
rect 806 22965 852 23011
rect 806 22858 852 22904
rect 806 22751 852 22797
rect 806 22644 852 22690
rect 806 22537 852 22583
rect 806 22430 852 22476
rect 806 22323 852 22369
rect 1030 23613 1076 23659
rect 1030 23505 1076 23551
rect 1030 23397 1076 23443
rect 1030 23289 1076 23335
rect 1030 23181 1076 23227
rect 1030 23073 1076 23119
rect 1030 22965 1076 23011
rect 1030 22858 1076 22904
rect 1030 22751 1076 22797
rect 1030 22644 1076 22690
rect 1030 22537 1076 22583
rect 1030 22430 1076 22476
rect 1030 22323 1076 22369
rect 1426 23613 1472 23659
rect 1426 23505 1472 23551
rect 1426 23397 1472 23443
rect 1426 23289 1472 23335
rect 1426 23181 1472 23227
rect 1426 23073 1472 23119
rect 1426 22965 1472 23011
rect 1426 22858 1472 22904
rect 1426 22751 1472 22797
rect 1426 22644 1472 22690
rect 1426 22537 1472 22583
rect 1426 22430 1472 22476
rect 1426 22323 1472 22369
rect 1650 23613 1696 23659
rect 1650 23505 1696 23551
rect 1650 23397 1696 23443
rect 1650 23289 1696 23335
rect 1650 23181 1696 23227
rect 1650 23073 1696 23119
rect 1650 22965 1696 23011
rect 1650 22858 1696 22904
rect 1650 22751 1696 22797
rect 1650 22644 1696 22690
rect 1650 22537 1696 22583
rect 1650 22430 1696 22476
rect 1650 22323 1696 22369
rect 2045 23613 2091 23659
rect 2045 23505 2091 23551
rect 2045 23397 2091 23443
rect 2045 23289 2091 23335
rect 2045 23181 2091 23227
rect 2045 23073 2091 23119
rect 2045 22965 2091 23011
rect 2045 22858 2091 22904
rect 2045 22751 2091 22797
rect 2045 22644 2091 22690
rect 2045 22537 2091 22583
rect 2045 22430 2091 22476
rect 2045 22323 2091 22369
rect 2269 23613 2315 23659
rect 2269 23505 2315 23551
rect 2269 23397 2315 23443
rect 2269 23289 2315 23335
rect 2269 23181 2315 23227
rect 2269 23073 2315 23119
rect 2269 22965 2315 23011
rect 2269 22858 2315 22904
rect 2269 22751 2315 22797
rect 2269 22644 2315 22690
rect 2269 22537 2315 22583
rect 2269 22430 2315 22476
rect 2269 22323 2315 22369
rect 2665 23613 2711 23659
rect 2665 23505 2711 23551
rect 2665 23397 2711 23443
rect 2665 23289 2711 23335
rect 2665 23181 2711 23227
rect 2665 23073 2711 23119
rect 2665 22965 2711 23011
rect 2665 22858 2711 22904
rect 2665 22751 2711 22797
rect 2665 22644 2711 22690
rect 2665 22537 2711 22583
rect 2665 22430 2711 22476
rect 2665 22323 2711 22369
rect 2889 23613 2935 23659
rect 2889 23505 2935 23551
rect 2889 23397 2935 23443
rect 2889 23289 2935 23335
rect 2889 23181 2935 23227
rect 2889 23073 2935 23119
rect 2889 22965 2935 23011
rect 2889 22858 2935 22904
rect 2889 22751 2935 22797
rect 2889 22644 2935 22690
rect 2889 22537 2935 22583
rect 2889 22430 2935 22476
rect 2889 22323 2935 22369
rect 3283 23613 3329 23659
rect 3283 23505 3329 23551
rect 3283 23397 3329 23443
rect 3283 23289 3329 23335
rect 3283 23181 3329 23227
rect 3283 23073 3329 23119
rect 3283 22965 3329 23011
rect 3283 22858 3329 22904
rect 3283 22751 3329 22797
rect 3283 22644 3329 22690
rect 3283 22537 3329 22583
rect 3283 22430 3329 22476
rect 3283 22323 3329 22369
rect 3507 23613 3553 23659
rect 3507 23505 3553 23551
rect 3507 23397 3553 23443
rect 3507 23289 3553 23335
rect 3507 23181 3553 23227
rect 3507 23073 3553 23119
rect 3507 22965 3553 23011
rect 3507 22858 3553 22904
rect 3507 22751 3553 22797
rect 3507 22644 3553 22690
rect 3507 22537 3553 22583
rect 3507 22430 3553 22476
rect 3507 22323 3553 22369
rect 3903 23613 3949 23659
rect 3903 23505 3949 23551
rect 3903 23397 3949 23443
rect 3903 23289 3949 23335
rect 3903 23181 3949 23227
rect 3903 23073 3949 23119
rect 3903 22965 3949 23011
rect 3903 22858 3949 22904
rect 3903 22751 3949 22797
rect 3903 22644 3949 22690
rect 3903 22537 3949 22583
rect 3903 22430 3949 22476
rect 3903 22323 3949 22369
rect 4127 23613 4173 23659
rect 4127 23505 4173 23551
rect 4127 23397 4173 23443
rect 4127 23289 4173 23335
rect 4127 23181 4173 23227
rect 4127 23073 4173 23119
rect 4127 22965 4173 23011
rect 4127 22858 4173 22904
rect 4127 22751 4173 22797
rect 4127 22644 4173 22690
rect 4127 22537 4173 22583
rect 4127 22430 4173 22476
rect 4127 22323 4173 22369
rect 4522 23613 4568 23659
rect 4522 23505 4568 23551
rect 4522 23397 4568 23443
rect 4522 23289 4568 23335
rect 4522 23181 4568 23227
rect 4522 23073 4568 23119
rect 4522 22965 4568 23011
rect 4522 22858 4568 22904
rect 4522 22751 4568 22797
rect 4522 22644 4568 22690
rect 4522 22537 4568 22583
rect 4522 22430 4568 22476
rect 4522 22323 4568 22369
rect 4746 23613 4792 23659
rect 4746 23505 4792 23551
rect 4746 23397 4792 23443
rect 4746 23289 4792 23335
rect 4746 23181 4792 23227
rect 4746 23073 4792 23119
rect 4746 22965 4792 23011
rect 4746 22858 4792 22904
rect 4746 22751 4792 22797
rect 4746 22644 4792 22690
rect 4746 22537 4792 22583
rect 4746 22430 4792 22476
rect 4746 22323 4792 22369
rect 5142 23613 5188 23659
rect 5142 23505 5188 23551
rect 5142 23397 5188 23443
rect 5142 23289 5188 23335
rect 5142 23181 5188 23227
rect 5142 23073 5188 23119
rect 5142 22965 5188 23011
rect 5142 22858 5188 22904
rect 5142 22751 5188 22797
rect 5142 22644 5188 22690
rect 5142 22537 5188 22583
rect 5142 22430 5188 22476
rect 5142 22323 5188 22369
rect 5366 23613 5412 23659
rect 5366 23505 5412 23551
rect 5366 23397 5412 23443
rect 5366 23289 5412 23335
rect 5366 23181 5412 23227
rect 5366 23073 5412 23119
rect 5366 22965 5412 23011
rect 5366 22858 5412 22904
rect 5366 22751 5412 22797
rect 5366 22644 5412 22690
rect 5366 22537 5412 22583
rect 5366 22430 5412 22476
rect 5366 22323 5412 22369
rect 806 21609 852 21655
rect 806 21501 852 21547
rect 806 21393 852 21439
rect 806 21285 852 21331
rect 806 21177 852 21223
rect 806 21069 852 21115
rect 806 20961 852 21007
rect 806 20854 852 20900
rect 806 20747 852 20793
rect 806 20640 852 20686
rect 806 20533 852 20579
rect 806 20426 852 20472
rect 806 20319 852 20365
rect 1030 21609 1076 21655
rect 1030 21501 1076 21547
rect 1030 21393 1076 21439
rect 1030 21285 1076 21331
rect 1030 21177 1076 21223
rect 1030 21069 1076 21115
rect 1030 20961 1076 21007
rect 1030 20854 1076 20900
rect 1030 20747 1076 20793
rect 1030 20640 1076 20686
rect 1030 20533 1076 20579
rect 1030 20426 1076 20472
rect 1030 20319 1076 20365
rect 1426 21609 1472 21655
rect 1426 21501 1472 21547
rect 1426 21393 1472 21439
rect 1426 21285 1472 21331
rect 1426 21177 1472 21223
rect 1426 21069 1472 21115
rect 1426 20961 1472 21007
rect 1426 20854 1472 20900
rect 1426 20747 1472 20793
rect 1426 20640 1472 20686
rect 1426 20533 1472 20579
rect 1426 20426 1472 20472
rect 1426 20319 1472 20365
rect 1650 21609 1696 21655
rect 1650 21501 1696 21547
rect 1650 21393 1696 21439
rect 1650 21285 1696 21331
rect 1650 21177 1696 21223
rect 1650 21069 1696 21115
rect 1650 20961 1696 21007
rect 1650 20854 1696 20900
rect 1650 20747 1696 20793
rect 1650 20640 1696 20686
rect 1650 20533 1696 20579
rect 1650 20426 1696 20472
rect 1650 20319 1696 20365
rect 2045 21609 2091 21655
rect 2045 21501 2091 21547
rect 2045 21393 2091 21439
rect 2045 21285 2091 21331
rect 2045 21177 2091 21223
rect 2045 21069 2091 21115
rect 2045 20961 2091 21007
rect 2045 20854 2091 20900
rect 2045 20747 2091 20793
rect 2045 20640 2091 20686
rect 2045 20533 2091 20579
rect 2045 20426 2091 20472
rect 2045 20319 2091 20365
rect 2269 21609 2315 21655
rect 2269 21501 2315 21547
rect 2269 21393 2315 21439
rect 2269 21285 2315 21331
rect 2269 21177 2315 21223
rect 2269 21069 2315 21115
rect 2269 20961 2315 21007
rect 2269 20854 2315 20900
rect 2269 20747 2315 20793
rect 2269 20640 2315 20686
rect 2269 20533 2315 20579
rect 2269 20426 2315 20472
rect 2269 20319 2315 20365
rect 2665 21609 2711 21655
rect 2665 21501 2711 21547
rect 2665 21393 2711 21439
rect 2665 21285 2711 21331
rect 2665 21177 2711 21223
rect 2665 21069 2711 21115
rect 2665 20961 2711 21007
rect 2665 20854 2711 20900
rect 2665 20747 2711 20793
rect 2665 20640 2711 20686
rect 2665 20533 2711 20579
rect 2665 20426 2711 20472
rect 2665 20319 2711 20365
rect 2889 21609 2935 21655
rect 2889 21501 2935 21547
rect 2889 21393 2935 21439
rect 2889 21285 2935 21331
rect 2889 21177 2935 21223
rect 2889 21069 2935 21115
rect 2889 20961 2935 21007
rect 2889 20854 2935 20900
rect 2889 20747 2935 20793
rect 2889 20640 2935 20686
rect 2889 20533 2935 20579
rect 2889 20426 2935 20472
rect 2889 20319 2935 20365
rect 3283 21609 3329 21655
rect 3283 21501 3329 21547
rect 3283 21393 3329 21439
rect 3283 21285 3329 21331
rect 3283 21177 3329 21223
rect 3283 21069 3329 21115
rect 3283 20961 3329 21007
rect 3283 20854 3329 20900
rect 3283 20747 3329 20793
rect 3283 20640 3329 20686
rect 3283 20533 3329 20579
rect 3283 20426 3329 20472
rect 3283 20319 3329 20365
rect 3507 21609 3553 21655
rect 3507 21501 3553 21547
rect 3507 21393 3553 21439
rect 3507 21285 3553 21331
rect 3507 21177 3553 21223
rect 3507 21069 3553 21115
rect 3507 20961 3553 21007
rect 3507 20854 3553 20900
rect 3507 20747 3553 20793
rect 3507 20640 3553 20686
rect 3507 20533 3553 20579
rect 3507 20426 3553 20472
rect 3507 20319 3553 20365
rect 3903 21609 3949 21655
rect 3903 21501 3949 21547
rect 3903 21393 3949 21439
rect 3903 21285 3949 21331
rect 3903 21177 3949 21223
rect 3903 21069 3949 21115
rect 3903 20961 3949 21007
rect 3903 20854 3949 20900
rect 3903 20747 3949 20793
rect 3903 20640 3949 20686
rect 3903 20533 3949 20579
rect 3903 20426 3949 20472
rect 3903 20319 3949 20365
rect 4127 21609 4173 21655
rect 4127 21501 4173 21547
rect 4127 21393 4173 21439
rect 4127 21285 4173 21331
rect 4127 21177 4173 21223
rect 4127 21069 4173 21115
rect 4127 20961 4173 21007
rect 4127 20854 4173 20900
rect 4127 20747 4173 20793
rect 4127 20640 4173 20686
rect 4127 20533 4173 20579
rect 4127 20426 4173 20472
rect 4127 20319 4173 20365
rect 4522 21609 4568 21655
rect 4522 21501 4568 21547
rect 4522 21393 4568 21439
rect 4522 21285 4568 21331
rect 4522 21177 4568 21223
rect 4522 21069 4568 21115
rect 4522 20961 4568 21007
rect 4522 20854 4568 20900
rect 4522 20747 4568 20793
rect 4522 20640 4568 20686
rect 4522 20533 4568 20579
rect 4522 20426 4568 20472
rect 4522 20319 4568 20365
rect 4746 21609 4792 21655
rect 4746 21501 4792 21547
rect 4746 21393 4792 21439
rect 4746 21285 4792 21331
rect 4746 21177 4792 21223
rect 4746 21069 4792 21115
rect 4746 20961 4792 21007
rect 4746 20854 4792 20900
rect 4746 20747 4792 20793
rect 4746 20640 4792 20686
rect 4746 20533 4792 20579
rect 4746 20426 4792 20472
rect 4746 20319 4792 20365
rect 5142 21609 5188 21655
rect 5142 21501 5188 21547
rect 5142 21393 5188 21439
rect 5142 21285 5188 21331
rect 5142 21177 5188 21223
rect 5142 21069 5188 21115
rect 5142 20961 5188 21007
rect 5142 20854 5188 20900
rect 5142 20747 5188 20793
rect 5142 20640 5188 20686
rect 5142 20533 5188 20579
rect 5142 20426 5188 20472
rect 5142 20319 5188 20365
rect 5366 21609 5412 21655
rect 5366 21501 5412 21547
rect 5366 21393 5412 21439
rect 5366 21285 5412 21331
rect 5366 21177 5412 21223
rect 5366 21069 5412 21115
rect 5366 20961 5412 21007
rect 5366 20854 5412 20900
rect 5366 20747 5412 20793
rect 5366 20640 5412 20686
rect 5366 20533 5412 20579
rect 5366 20426 5412 20472
rect 5366 20319 5412 20365
rect 780 17170 826 17216
rect 1004 17170 1050 17216
rect 1228 17170 1274 17216
rect 1452 17170 1498 17216
rect 1676 17170 1722 17216
rect 2019 17170 2065 17216
rect 2243 17170 2289 17216
rect 2467 17170 2513 17216
rect 2691 17170 2737 17216
rect 2915 17170 2961 17216
rect 3257 17170 3303 17216
rect 3481 17170 3527 17216
rect 3705 17170 3751 17216
rect 3929 17170 3975 17216
rect 4153 17170 4199 17216
rect 4496 17170 4542 17216
rect 4720 17170 4766 17216
rect 4944 17170 4990 17216
rect 5168 17170 5214 17216
rect 5392 17170 5438 17216
rect 948 15538 994 15584
rect 1211 15538 1257 15584
rect 300 9904 346 12600
rect 524 9904 570 12600
rect 748 12553 794 12599
rect 748 12449 794 12495
rect 748 12345 794 12391
rect 748 12241 794 12287
rect 748 12137 794 12183
rect 748 12033 794 12079
rect 748 11929 794 11975
rect 748 11825 794 11871
rect 748 11721 794 11767
rect 748 11617 794 11663
rect 748 11512 794 11558
rect 748 11407 794 11453
rect 748 11302 794 11348
rect 748 11197 794 11243
rect 748 11092 794 11138
rect 748 10987 794 11033
rect 748 10882 794 10928
rect 748 10777 794 10823
rect 748 10672 794 10718
rect 748 10567 794 10613
rect 748 10462 794 10508
rect 748 10357 794 10403
rect 972 12553 1018 12599
rect 972 12449 1018 12495
rect 972 12345 1018 12391
rect 972 12241 1018 12287
rect 972 12137 1018 12183
rect 972 12033 1018 12079
rect 972 11929 1018 11975
rect 972 11825 1018 11871
rect 972 11721 1018 11767
rect 972 11617 1018 11663
rect 972 11512 1018 11558
rect 972 11407 1018 11453
rect 972 11302 1018 11348
rect 972 11197 1018 11243
rect 972 11092 1018 11138
rect 972 10987 1018 11033
rect 972 10882 1018 10928
rect 972 10777 1018 10823
rect 972 10672 1018 10718
rect 972 10567 1018 10613
rect 972 10462 1018 10508
rect 972 10357 1018 10403
rect 1196 12553 1242 12599
rect 1196 12449 1242 12495
rect 1196 12345 1242 12391
rect 1196 12241 1242 12287
rect 1196 12137 1242 12183
rect 1196 12033 1242 12079
rect 1196 11929 1242 11975
rect 1196 11825 1242 11871
rect 1196 11721 1242 11767
rect 1196 11617 1242 11663
rect 1196 11512 1242 11558
rect 1196 11407 1242 11453
rect 1196 11302 1242 11348
rect 1196 11197 1242 11243
rect 1196 11092 1242 11138
rect 1196 10987 1242 11033
rect 1196 10882 1242 10928
rect 1196 10777 1242 10823
rect 1196 10672 1242 10718
rect 1196 10567 1242 10613
rect 1196 10462 1242 10508
rect 1196 10357 1242 10403
rect 1420 12553 1466 12599
rect 1420 12449 1466 12495
rect 1420 12345 1466 12391
rect 1420 12241 1466 12287
rect 1420 12137 1466 12183
rect 1420 12033 1466 12079
rect 1420 11929 1466 11975
rect 1420 11825 1466 11871
rect 1420 11721 1466 11767
rect 1420 11617 1466 11663
rect 1420 11512 1466 11558
rect 1420 11407 1466 11453
rect 1420 11302 1466 11348
rect 1420 11197 1466 11243
rect 1420 11092 1466 11138
rect 1420 10987 1466 11033
rect 1420 10882 1466 10928
rect 1420 10777 1466 10823
rect 1420 10672 1466 10718
rect 1420 10567 1466 10613
rect 1420 10462 1466 10508
rect 1420 10357 1466 10403
rect 1644 12553 1690 12599
rect 1644 12449 1690 12495
rect 1644 12345 1690 12391
rect 1644 12241 1690 12287
rect 1644 12137 1690 12183
rect 1644 12033 1690 12079
rect 1644 11929 1690 11975
rect 1644 11825 1690 11871
rect 1644 11721 1690 11767
rect 1644 11617 1690 11663
rect 1644 11512 1690 11558
rect 1644 11407 1690 11453
rect 1644 11302 1690 11348
rect 1644 11197 1690 11243
rect 1644 11092 1690 11138
rect 1644 10987 1690 11033
rect 1644 10882 1690 10928
rect 1644 10777 1690 10823
rect 1644 10672 1690 10718
rect 1644 10567 1690 10613
rect 1644 10462 1690 10508
rect 1644 10357 1690 10403
rect 1868 12553 1914 12599
rect 1868 12449 1914 12495
rect 1868 12345 1914 12391
rect 1868 12241 1914 12287
rect 1868 12137 1914 12183
rect 1868 12033 1914 12079
rect 1868 11929 1914 11975
rect 1868 11825 1914 11871
rect 1868 11721 1914 11767
rect 1868 11617 1914 11663
rect 1868 11512 1914 11558
rect 1868 11407 1914 11453
rect 1868 11302 1914 11348
rect 1868 11197 1914 11243
rect 1868 11092 1914 11138
rect 1868 10987 1914 11033
rect 1868 10882 1914 10928
rect 1868 10777 1914 10823
rect 1868 10672 1914 10718
rect 1868 10567 1914 10613
rect 1868 10462 1914 10508
rect 1868 10357 1914 10403
rect 2481 9931 2527 9977
rect 1629 9845 1675 9891
rect 911 9745 957 9791
rect 911 9625 957 9671
rect 1135 9745 1181 9791
rect 1629 9725 1675 9771
rect 1853 9845 1899 9891
rect 1853 9725 1899 9771
rect 2481 9803 2527 9849
rect 1135 9625 1181 9671
rect 2481 9676 2527 9722
rect 2481 9549 2527 9595
rect 2705 9931 2751 9977
rect 2705 9803 2751 9849
rect 2705 9676 2751 9722
rect 2705 9549 2751 9595
rect 801 8104 847 8150
rect 801 7984 847 8030
rect 1025 8104 1071 8150
rect 1025 7984 1071 8030
rect 1249 8104 1295 8150
rect 1249 7984 1295 8030
rect 1629 8083 1675 8129
rect 1629 7963 1675 8009
rect 1853 8083 1899 8129
rect 1853 7963 1899 8009
rect 2077 8083 2123 8129
rect 2077 7963 2123 8009
<< mvpdiffc >>
rect 692 28535 738 28581
rect 692 28353 738 28399
rect 692 28172 738 28218
rect 692 27990 738 28036
rect 918 28535 964 28581
rect 918 28353 964 28399
rect 918 28172 964 28218
rect 918 27990 964 28036
rect 1228 28535 1274 28581
rect 1228 28353 1274 28399
rect 1228 28172 1274 28218
rect 1228 27990 1274 28036
rect 1538 28535 1584 28581
rect 1538 28353 1584 28399
rect 1538 28172 1584 28218
rect 1538 27990 1584 28036
rect 1764 28535 1810 28581
rect 1931 28535 1977 28581
rect 1764 28353 1810 28399
rect 1931 28353 1977 28399
rect 1764 28172 1810 28218
rect 1931 28172 1977 28218
rect 1764 27990 1810 28036
rect 1931 27990 1977 28036
rect 2157 28535 2203 28581
rect 2157 28353 2203 28399
rect 2157 28172 2203 28218
rect 2157 27990 2203 28036
rect 2467 28535 2513 28581
rect 2467 28353 2513 28399
rect 2467 28172 2513 28218
rect 2467 27990 2513 28036
rect 2777 28535 2823 28581
rect 2777 28353 2823 28399
rect 2777 28172 2823 28218
rect 2777 27990 2823 28036
rect 3003 28535 3049 28581
rect 3169 28535 3215 28581
rect 3003 28353 3049 28399
rect 3169 28353 3215 28399
rect 3003 28172 3049 28218
rect 3169 28172 3215 28218
rect 3003 27990 3049 28036
rect 3169 27990 3215 28036
rect 3395 28535 3441 28581
rect 3395 28353 3441 28399
rect 3395 28172 3441 28218
rect 3395 27990 3441 28036
rect 3705 28535 3751 28581
rect 3705 28353 3751 28399
rect 3705 28172 3751 28218
rect 3705 27990 3751 28036
rect 4015 28535 4061 28581
rect 4015 28353 4061 28399
rect 4015 28172 4061 28218
rect 4015 27990 4061 28036
rect 4241 28535 4287 28581
rect 4408 28535 4454 28581
rect 4241 28353 4287 28399
rect 4408 28353 4454 28399
rect 4241 28172 4287 28218
rect 4408 28172 4454 28218
rect 4241 27990 4287 28036
rect 4408 27990 4454 28036
rect 4634 28535 4680 28581
rect 4634 28353 4680 28399
rect 4634 28172 4680 28218
rect 4634 27990 4680 28036
rect 4944 28535 4990 28581
rect 4944 28353 4990 28399
rect 4944 28172 4990 28218
rect 4944 27990 4990 28036
rect 5219 28535 5265 28581
rect 5219 28353 5265 28399
rect 5219 28172 5265 28218
rect 5219 27990 5265 28036
rect 5480 28535 5526 28581
rect 5480 28353 5526 28399
rect 5480 28172 5526 28218
rect 5480 27990 5526 28036
rect 692 27759 738 27805
rect 692 27578 738 27624
rect 692 27397 738 27443
rect 692 27215 738 27261
rect 918 27759 964 27805
rect 918 27578 964 27624
rect 918 27397 964 27443
rect 918 27215 964 27261
rect 1228 27759 1274 27805
rect 1228 27578 1274 27624
rect 1228 27397 1274 27443
rect 1228 27215 1274 27261
rect 1538 27759 1584 27805
rect 1538 27578 1584 27624
rect 1538 27397 1584 27443
rect 1538 27215 1584 27261
rect 1764 27759 1810 27805
rect 1931 27759 1977 27805
rect 1764 27578 1810 27624
rect 1931 27578 1977 27624
rect 1764 27397 1810 27443
rect 1931 27397 1977 27443
rect 1764 27215 1810 27261
rect 1931 27215 1977 27261
rect 2157 27759 2203 27805
rect 2157 27578 2203 27624
rect 2157 27397 2203 27443
rect 2157 27215 2203 27261
rect 2467 27759 2513 27805
rect 2467 27578 2513 27624
rect 2467 27397 2513 27443
rect 2467 27215 2513 27261
rect 2777 27759 2823 27805
rect 2777 27578 2823 27624
rect 2777 27397 2823 27443
rect 2777 27215 2823 27261
rect 3003 27759 3049 27805
rect 3169 27759 3215 27805
rect 3003 27578 3049 27624
rect 3169 27578 3215 27624
rect 3003 27397 3049 27443
rect 3169 27397 3215 27443
rect 3003 27215 3049 27261
rect 3169 27215 3215 27261
rect 3395 27759 3441 27805
rect 3395 27578 3441 27624
rect 3395 27397 3441 27443
rect 3395 27215 3441 27261
rect 3705 27759 3751 27805
rect 3705 27578 3751 27624
rect 3705 27397 3751 27443
rect 3705 27215 3751 27261
rect 4015 27759 4061 27805
rect 4015 27578 4061 27624
rect 4015 27397 4061 27443
rect 4015 27215 4061 27261
rect 4241 27759 4287 27805
rect 4408 27759 4454 27805
rect 4241 27578 4287 27624
rect 4408 27578 4454 27624
rect 4241 27397 4287 27443
rect 4408 27397 4454 27443
rect 4241 27215 4287 27261
rect 4408 27215 4454 27261
rect 4634 27759 4680 27805
rect 4634 27578 4680 27624
rect 4634 27397 4680 27443
rect 4634 27215 4680 27261
rect 4944 27759 4990 27805
rect 4944 27578 4990 27624
rect 4944 27397 4990 27443
rect 4944 27215 4990 27261
rect 5219 27759 5265 27805
rect 5219 27578 5265 27624
rect 5219 27397 5265 27443
rect 5219 27215 5265 27261
rect 5480 27759 5526 27805
rect 5480 27578 5526 27624
rect 5480 27397 5526 27443
rect 5480 27215 5526 27261
rect 808 26891 854 26937
rect 808 26783 854 26829
rect 808 26675 854 26721
rect 808 26567 854 26613
rect 808 26459 854 26505
rect 808 26351 854 26397
rect 808 26243 854 26289
rect 808 26136 854 26182
rect 808 26029 854 26075
rect 808 25922 854 25968
rect 808 25815 854 25861
rect 808 25708 854 25754
rect 808 25601 854 25647
rect 1032 26891 1078 26937
rect 1032 26783 1078 26829
rect 1032 26675 1078 26721
rect 1032 26567 1078 26613
rect 1032 26459 1078 26505
rect 1032 26351 1078 26397
rect 1032 26243 1078 26289
rect 1032 26136 1078 26182
rect 1032 26029 1078 26075
rect 1032 25922 1078 25968
rect 1032 25815 1078 25861
rect 1032 25708 1078 25754
rect 1032 25601 1078 25647
rect 1424 26891 1470 26937
rect 1424 26783 1470 26829
rect 1424 26675 1470 26721
rect 1424 26567 1470 26613
rect 1424 26459 1470 26505
rect 1424 26351 1470 26397
rect 1424 26243 1470 26289
rect 1424 26136 1470 26182
rect 1424 26029 1470 26075
rect 1424 25922 1470 25968
rect 1424 25815 1470 25861
rect 1424 25708 1470 25754
rect 1424 25601 1470 25647
rect 1648 26891 1694 26937
rect 1648 26783 1694 26829
rect 1648 26675 1694 26721
rect 1648 26567 1694 26613
rect 1648 26459 1694 26505
rect 1648 26351 1694 26397
rect 1648 26243 1694 26289
rect 1648 26136 1694 26182
rect 1648 26029 1694 26075
rect 1648 25922 1694 25968
rect 1648 25815 1694 25861
rect 1648 25708 1694 25754
rect 1648 25601 1694 25647
rect 2047 26891 2093 26937
rect 2047 26783 2093 26829
rect 2047 26675 2093 26721
rect 2047 26567 2093 26613
rect 2047 26459 2093 26505
rect 2047 26351 2093 26397
rect 2047 26243 2093 26289
rect 2047 26136 2093 26182
rect 2047 26029 2093 26075
rect 2047 25922 2093 25968
rect 2047 25815 2093 25861
rect 2047 25708 2093 25754
rect 2047 25601 2093 25647
rect 2271 26891 2317 26937
rect 2271 26783 2317 26829
rect 2271 26675 2317 26721
rect 2271 26567 2317 26613
rect 2271 26459 2317 26505
rect 2271 26351 2317 26397
rect 2271 26243 2317 26289
rect 2271 26136 2317 26182
rect 2271 26029 2317 26075
rect 2271 25922 2317 25968
rect 2271 25815 2317 25861
rect 2271 25708 2317 25754
rect 2271 25601 2317 25647
rect 2663 26891 2709 26937
rect 2663 26783 2709 26829
rect 2663 26675 2709 26721
rect 2663 26567 2709 26613
rect 2663 26459 2709 26505
rect 2663 26351 2709 26397
rect 2663 26243 2709 26289
rect 2663 26136 2709 26182
rect 2663 26029 2709 26075
rect 2663 25922 2709 25968
rect 2663 25815 2709 25861
rect 2663 25708 2709 25754
rect 2663 25601 2709 25647
rect 2887 26891 2933 26937
rect 2887 26783 2933 26829
rect 2887 26675 2933 26721
rect 2887 26567 2933 26613
rect 2887 26459 2933 26505
rect 2887 26351 2933 26397
rect 2887 26243 2933 26289
rect 2887 26136 2933 26182
rect 2887 26029 2933 26075
rect 2887 25922 2933 25968
rect 2887 25815 2933 25861
rect 2887 25708 2933 25754
rect 2887 25601 2933 25647
rect 3285 26891 3331 26937
rect 3285 26783 3331 26829
rect 3285 26675 3331 26721
rect 3285 26567 3331 26613
rect 3285 26459 3331 26505
rect 3285 26351 3331 26397
rect 3285 26243 3331 26289
rect 3285 26136 3331 26182
rect 3285 26029 3331 26075
rect 3285 25922 3331 25968
rect 3285 25815 3331 25861
rect 3285 25708 3331 25754
rect 3285 25601 3331 25647
rect 3509 26891 3555 26937
rect 3509 26783 3555 26829
rect 3509 26675 3555 26721
rect 3509 26567 3555 26613
rect 3509 26459 3555 26505
rect 3509 26351 3555 26397
rect 3509 26243 3555 26289
rect 3509 26136 3555 26182
rect 3509 26029 3555 26075
rect 3509 25922 3555 25968
rect 3509 25815 3555 25861
rect 3509 25708 3555 25754
rect 3509 25601 3555 25647
rect 3901 26891 3947 26937
rect 3901 26783 3947 26829
rect 3901 26675 3947 26721
rect 3901 26567 3947 26613
rect 3901 26459 3947 26505
rect 3901 26351 3947 26397
rect 3901 26243 3947 26289
rect 3901 26136 3947 26182
rect 3901 26029 3947 26075
rect 3901 25922 3947 25968
rect 3901 25815 3947 25861
rect 3901 25708 3947 25754
rect 3901 25601 3947 25647
rect 4125 26891 4171 26937
rect 4125 26783 4171 26829
rect 4125 26675 4171 26721
rect 4125 26567 4171 26613
rect 4125 26459 4171 26505
rect 4125 26351 4171 26397
rect 4125 26243 4171 26289
rect 4125 26136 4171 26182
rect 4125 26029 4171 26075
rect 4125 25922 4171 25968
rect 4125 25815 4171 25861
rect 4125 25708 4171 25754
rect 4125 25601 4171 25647
rect 4524 26891 4570 26937
rect 4524 26783 4570 26829
rect 4524 26675 4570 26721
rect 4524 26567 4570 26613
rect 4524 26459 4570 26505
rect 4524 26351 4570 26397
rect 4524 26243 4570 26289
rect 4524 26136 4570 26182
rect 4524 26029 4570 26075
rect 4524 25922 4570 25968
rect 4524 25815 4570 25861
rect 4524 25708 4570 25754
rect 4524 25601 4570 25647
rect 4748 26891 4794 26937
rect 4748 26783 4794 26829
rect 4748 26675 4794 26721
rect 4748 26567 4794 26613
rect 4748 26459 4794 26505
rect 4748 26351 4794 26397
rect 4748 26243 4794 26289
rect 4748 26136 4794 26182
rect 4748 26029 4794 26075
rect 4748 25922 4794 25968
rect 4748 25815 4794 25861
rect 4748 25708 4794 25754
rect 4748 25601 4794 25647
rect 5140 26891 5186 26937
rect 5140 26783 5186 26829
rect 5140 26675 5186 26721
rect 5140 26567 5186 26613
rect 5140 26459 5186 26505
rect 5140 26351 5186 26397
rect 5140 26243 5186 26289
rect 5140 26136 5186 26182
rect 5140 26029 5186 26075
rect 5140 25922 5186 25968
rect 5140 25815 5186 25861
rect 5140 25708 5186 25754
rect 5140 25601 5186 25647
rect 5364 26891 5410 26937
rect 5364 26783 5410 26829
rect 5364 26675 5410 26721
rect 5364 26567 5410 26613
rect 5364 26459 5410 26505
rect 5364 26351 5410 26397
rect 5364 26243 5410 26289
rect 5364 26136 5410 26182
rect 5364 26029 5410 26075
rect 5364 25922 5410 25968
rect 5364 25815 5410 25861
rect 5364 25708 5410 25754
rect 5364 25601 5410 25647
rect 806 25304 852 25350
rect 806 25196 852 25242
rect 806 25088 852 25134
rect 806 24980 852 25026
rect 806 24872 852 24918
rect 806 24764 852 24810
rect 806 24656 852 24702
rect 806 24549 852 24595
rect 806 24442 852 24488
rect 806 24335 852 24381
rect 806 24228 852 24274
rect 806 24121 852 24167
rect 806 24014 852 24060
rect 1030 25304 1076 25350
rect 1030 25196 1076 25242
rect 1030 25088 1076 25134
rect 1030 24980 1076 25026
rect 1030 24872 1076 24918
rect 1030 24764 1076 24810
rect 1030 24656 1076 24702
rect 1426 25304 1472 25350
rect 1426 25196 1472 25242
rect 1426 25088 1472 25134
rect 1426 24980 1472 25026
rect 1426 24872 1472 24918
rect 1426 24764 1472 24810
rect 1030 24549 1076 24595
rect 1030 24442 1076 24488
rect 1426 24656 1472 24702
rect 1426 24549 1472 24595
rect 1426 24442 1472 24488
rect 1030 24335 1076 24381
rect 1030 24228 1076 24274
rect 1030 24121 1076 24167
rect 1030 24014 1076 24060
rect 1426 24335 1472 24381
rect 1426 24228 1472 24274
rect 1426 24121 1472 24167
rect 1426 24014 1472 24060
rect 1650 25304 1696 25350
rect 1650 25196 1696 25242
rect 1650 25088 1696 25134
rect 1650 24980 1696 25026
rect 1650 24872 1696 24918
rect 1650 24764 1696 24810
rect 1650 24656 1696 24702
rect 1650 24549 1696 24595
rect 1650 24442 1696 24488
rect 1650 24335 1696 24381
rect 1650 24228 1696 24274
rect 1650 24121 1696 24167
rect 1650 24014 1696 24060
rect 2045 25304 2091 25350
rect 2045 25196 2091 25242
rect 2045 25088 2091 25134
rect 2045 24980 2091 25026
rect 2045 24872 2091 24918
rect 2045 24764 2091 24810
rect 2045 24656 2091 24702
rect 2045 24549 2091 24595
rect 2045 24442 2091 24488
rect 2045 24335 2091 24381
rect 2045 24228 2091 24274
rect 2045 24121 2091 24167
rect 2045 24014 2091 24060
rect 2269 25304 2315 25350
rect 2269 25196 2315 25242
rect 2269 25088 2315 25134
rect 2269 24980 2315 25026
rect 2269 24872 2315 24918
rect 2269 24764 2315 24810
rect 2269 24656 2315 24702
rect 2665 25304 2711 25350
rect 2665 25196 2711 25242
rect 2665 25088 2711 25134
rect 2665 24980 2711 25026
rect 2665 24872 2711 24918
rect 2665 24764 2711 24810
rect 2269 24549 2315 24595
rect 2269 24442 2315 24488
rect 2665 24656 2711 24702
rect 2665 24549 2711 24595
rect 2665 24442 2711 24488
rect 2269 24335 2315 24381
rect 2269 24228 2315 24274
rect 2269 24121 2315 24167
rect 2269 24014 2315 24060
rect 2665 24335 2711 24381
rect 2665 24228 2711 24274
rect 2665 24121 2711 24167
rect 2665 24014 2711 24060
rect 2889 25304 2935 25350
rect 2889 25196 2935 25242
rect 2889 25088 2935 25134
rect 2889 24980 2935 25026
rect 2889 24872 2935 24918
rect 2889 24764 2935 24810
rect 2889 24656 2935 24702
rect 2889 24549 2935 24595
rect 2889 24442 2935 24488
rect 2889 24335 2935 24381
rect 2889 24228 2935 24274
rect 2889 24121 2935 24167
rect 2889 24014 2935 24060
rect 3283 25304 3329 25350
rect 3283 25196 3329 25242
rect 3283 25088 3329 25134
rect 3283 24980 3329 25026
rect 3283 24872 3329 24918
rect 3283 24764 3329 24810
rect 3283 24656 3329 24702
rect 3283 24549 3329 24595
rect 3283 24442 3329 24488
rect 3283 24335 3329 24381
rect 3283 24228 3329 24274
rect 3283 24121 3329 24167
rect 3283 24014 3329 24060
rect 3507 25304 3553 25350
rect 3507 25196 3553 25242
rect 3507 25088 3553 25134
rect 3507 24980 3553 25026
rect 3507 24872 3553 24918
rect 3507 24764 3553 24810
rect 3507 24656 3553 24702
rect 3903 25304 3949 25350
rect 3903 25196 3949 25242
rect 3903 25088 3949 25134
rect 3903 24980 3949 25026
rect 3903 24872 3949 24918
rect 3903 24764 3949 24810
rect 3507 24549 3553 24595
rect 3507 24442 3553 24488
rect 3903 24656 3949 24702
rect 3903 24549 3949 24595
rect 3903 24442 3949 24488
rect 3507 24335 3553 24381
rect 3507 24228 3553 24274
rect 3507 24121 3553 24167
rect 3507 24014 3553 24060
rect 3903 24335 3949 24381
rect 3903 24228 3949 24274
rect 3903 24121 3949 24167
rect 3903 24014 3949 24060
rect 4127 25304 4173 25350
rect 4127 25196 4173 25242
rect 4127 25088 4173 25134
rect 4127 24980 4173 25026
rect 4127 24872 4173 24918
rect 4127 24764 4173 24810
rect 4127 24656 4173 24702
rect 4127 24549 4173 24595
rect 4127 24442 4173 24488
rect 4127 24335 4173 24381
rect 4127 24228 4173 24274
rect 4127 24121 4173 24167
rect 4127 24014 4173 24060
rect 4522 25304 4568 25350
rect 4522 25196 4568 25242
rect 4522 25088 4568 25134
rect 4522 24980 4568 25026
rect 4522 24872 4568 24918
rect 4522 24764 4568 24810
rect 4522 24656 4568 24702
rect 4522 24549 4568 24595
rect 4522 24442 4568 24488
rect 4522 24335 4568 24381
rect 4522 24228 4568 24274
rect 4522 24121 4568 24167
rect 4522 24014 4568 24060
rect 4746 25304 4792 25350
rect 4746 25196 4792 25242
rect 4746 25088 4792 25134
rect 4746 24980 4792 25026
rect 4746 24872 4792 24918
rect 4746 24764 4792 24810
rect 4746 24656 4792 24702
rect 5142 25304 5188 25350
rect 5142 25196 5188 25242
rect 5142 25088 5188 25134
rect 5142 24980 5188 25026
rect 5142 24872 5188 24918
rect 5142 24764 5188 24810
rect 4746 24549 4792 24595
rect 4746 24442 4792 24488
rect 5142 24656 5188 24702
rect 5142 24549 5188 24595
rect 5142 24442 5188 24488
rect 4746 24335 4792 24381
rect 4746 24228 4792 24274
rect 4746 24121 4792 24167
rect 4746 24014 4792 24060
rect 5142 24335 5188 24381
rect 5142 24228 5188 24274
rect 5142 24121 5188 24167
rect 5142 24014 5188 24060
rect 5366 25304 5412 25350
rect 5366 25196 5412 25242
rect 5366 25088 5412 25134
rect 5366 24980 5412 25026
rect 5366 24872 5412 24918
rect 5366 24764 5412 24810
rect 5366 24656 5412 24702
rect 5366 24549 5412 24595
rect 5366 24442 5412 24488
rect 5366 24335 5412 24381
rect 5366 24228 5412 24274
rect 5366 24121 5412 24167
rect 5366 24014 5412 24060
rect 806 19754 852 19800
rect 806 19646 852 19692
rect 806 19538 852 19584
rect 806 19430 852 19476
rect 806 19322 852 19368
rect 806 19214 852 19260
rect 806 19106 852 19152
rect 806 18999 852 19045
rect 806 18892 852 18938
rect 806 18785 852 18831
rect 806 18678 852 18724
rect 806 18571 852 18617
rect 806 18464 852 18510
rect 1030 19754 1076 19800
rect 1030 19646 1076 19692
rect 1030 19538 1076 19584
rect 1030 19430 1076 19476
rect 1030 19322 1076 19368
rect 1030 19214 1076 19260
rect 1030 19106 1076 19152
rect 1030 18999 1076 19045
rect 1030 18892 1076 18938
rect 1030 18785 1076 18831
rect 1030 18678 1076 18724
rect 1030 18571 1076 18617
rect 1030 18464 1076 18510
rect 1426 19754 1472 19800
rect 1426 19646 1472 19692
rect 1426 19538 1472 19584
rect 1426 19430 1472 19476
rect 1426 19322 1472 19368
rect 1426 19214 1472 19260
rect 1426 19106 1472 19152
rect 1426 18999 1472 19045
rect 1426 18892 1472 18938
rect 1426 18785 1472 18831
rect 1426 18678 1472 18724
rect 1426 18571 1472 18617
rect 1426 18464 1472 18510
rect 1650 19754 1696 19800
rect 1650 19646 1696 19692
rect 1650 19538 1696 19584
rect 1650 19430 1696 19476
rect 1650 19322 1696 19368
rect 1650 19214 1696 19260
rect 1650 19106 1696 19152
rect 1650 18999 1696 19045
rect 1650 18892 1696 18938
rect 1650 18785 1696 18831
rect 1650 18678 1696 18724
rect 1650 18571 1696 18617
rect 1650 18464 1696 18510
rect 2045 19754 2091 19800
rect 2045 19646 2091 19692
rect 2045 19538 2091 19584
rect 2045 19430 2091 19476
rect 2045 19322 2091 19368
rect 2045 19214 2091 19260
rect 2045 19106 2091 19152
rect 2045 18999 2091 19045
rect 2045 18892 2091 18938
rect 2045 18785 2091 18831
rect 2045 18678 2091 18724
rect 2045 18571 2091 18617
rect 2045 18464 2091 18510
rect 2269 19754 2315 19800
rect 2269 19646 2315 19692
rect 2269 19538 2315 19584
rect 2269 19430 2315 19476
rect 2269 19322 2315 19368
rect 2269 19214 2315 19260
rect 2269 19106 2315 19152
rect 2269 18999 2315 19045
rect 2269 18892 2315 18938
rect 2269 18785 2315 18831
rect 2269 18678 2315 18724
rect 2269 18571 2315 18617
rect 2269 18464 2315 18510
rect 2665 19754 2711 19800
rect 2665 19646 2711 19692
rect 2665 19538 2711 19584
rect 2665 19430 2711 19476
rect 2665 19322 2711 19368
rect 2665 19214 2711 19260
rect 2665 19106 2711 19152
rect 2665 18999 2711 19045
rect 2665 18892 2711 18938
rect 2665 18785 2711 18831
rect 2665 18678 2711 18724
rect 2665 18571 2711 18617
rect 2665 18464 2711 18510
rect 2889 19754 2935 19800
rect 2889 19646 2935 19692
rect 2889 19538 2935 19584
rect 2889 19430 2935 19476
rect 2889 19322 2935 19368
rect 2889 19214 2935 19260
rect 2889 19106 2935 19152
rect 2889 18999 2935 19045
rect 2889 18892 2935 18938
rect 2889 18785 2935 18831
rect 2889 18678 2935 18724
rect 2889 18571 2935 18617
rect 2889 18464 2935 18510
rect 3283 19754 3329 19800
rect 3283 19646 3329 19692
rect 3283 19538 3329 19584
rect 3283 19430 3329 19476
rect 3283 19322 3329 19368
rect 3283 19214 3329 19260
rect 3283 19106 3329 19152
rect 3283 18999 3329 19045
rect 3283 18892 3329 18938
rect 3283 18785 3329 18831
rect 3283 18678 3329 18724
rect 3283 18571 3329 18617
rect 3283 18464 3329 18510
rect 3507 19754 3553 19800
rect 3507 19646 3553 19692
rect 3507 19538 3553 19584
rect 3507 19430 3553 19476
rect 3507 19322 3553 19368
rect 3507 19214 3553 19260
rect 3507 19106 3553 19152
rect 3507 18999 3553 19045
rect 3507 18892 3553 18938
rect 3507 18785 3553 18831
rect 3507 18678 3553 18724
rect 3507 18571 3553 18617
rect 3507 18464 3553 18510
rect 3903 19754 3949 19800
rect 3903 19646 3949 19692
rect 3903 19538 3949 19584
rect 3903 19430 3949 19476
rect 3903 19322 3949 19368
rect 3903 19214 3949 19260
rect 3903 19106 3949 19152
rect 3903 18999 3949 19045
rect 3903 18892 3949 18938
rect 3903 18785 3949 18831
rect 3903 18678 3949 18724
rect 3903 18571 3949 18617
rect 3903 18464 3949 18510
rect 4127 19754 4173 19800
rect 4127 19646 4173 19692
rect 4127 19538 4173 19584
rect 4127 19430 4173 19476
rect 4127 19322 4173 19368
rect 4127 19214 4173 19260
rect 4127 19106 4173 19152
rect 4127 18999 4173 19045
rect 4127 18892 4173 18938
rect 4127 18785 4173 18831
rect 4127 18678 4173 18724
rect 4127 18571 4173 18617
rect 4127 18464 4173 18510
rect 4522 19754 4568 19800
rect 4522 19646 4568 19692
rect 4522 19538 4568 19584
rect 4522 19430 4568 19476
rect 4522 19322 4568 19368
rect 4522 19214 4568 19260
rect 4522 19106 4568 19152
rect 4522 18999 4568 19045
rect 4522 18892 4568 18938
rect 4522 18785 4568 18831
rect 4522 18678 4568 18724
rect 4522 18571 4568 18617
rect 4522 18464 4568 18510
rect 4746 19754 4792 19800
rect 4746 19646 4792 19692
rect 4746 19538 4792 19584
rect 4746 19430 4792 19476
rect 4746 19322 4792 19368
rect 4746 19214 4792 19260
rect 4746 19106 4792 19152
rect 4746 18999 4792 19045
rect 4746 18892 4792 18938
rect 4746 18785 4792 18831
rect 4746 18678 4792 18724
rect 4746 18571 4792 18617
rect 4746 18464 4792 18510
rect 5142 19754 5188 19800
rect 5142 19646 5188 19692
rect 5142 19538 5188 19584
rect 5142 19430 5188 19476
rect 5142 19322 5188 19368
rect 5142 19214 5188 19260
rect 5142 19106 5188 19152
rect 5142 18999 5188 19045
rect 5142 18892 5188 18938
rect 5142 18785 5188 18831
rect 5142 18678 5188 18724
rect 5142 18571 5188 18617
rect 5142 18464 5188 18510
rect 5366 19754 5412 19800
rect 5366 19646 5412 19692
rect 5366 19538 5412 19584
rect 5366 19430 5412 19476
rect 5366 19322 5412 19368
rect 5366 19214 5412 19260
rect 5366 19106 5412 19152
rect 5366 18999 5412 19045
rect 5366 18892 5412 18938
rect 5366 18785 5412 18831
rect 5366 18678 5412 18724
rect 5366 18571 5412 18617
rect 5366 18464 5412 18510
rect 725 17667 771 17713
rect 975 17667 1021 17713
rect 1228 17667 1274 17713
rect 1481 17667 1527 17713
rect 1731 17667 1777 17713
rect 1964 17667 2010 17713
rect 2214 17667 2260 17713
rect 2467 17667 2513 17713
rect 2720 17667 2766 17713
rect 2970 17667 3016 17713
rect 3202 17667 3248 17713
rect 3452 17667 3498 17713
rect 3705 17667 3751 17713
rect 3958 17667 4004 17713
rect 4208 17667 4254 17713
rect 4441 17667 4487 17713
rect 4691 17667 4737 17713
rect 4944 17667 4990 17713
rect 5197 17667 5243 17713
rect 5447 17667 5493 17713
rect 300 13062 346 15758
rect 524 13062 570 15758
rect 1644 15258 1690 15304
rect 853 15019 899 15065
rect 1117 15019 1163 15065
rect 1350 15019 1396 15065
rect 1644 15154 1690 15200
rect 1644 15050 1690 15096
rect 1644 14946 1690 14992
rect 1644 14842 1690 14888
rect 1644 14738 1690 14784
rect 1644 14634 1690 14680
rect 1644 14530 1690 14576
rect 1644 14426 1690 14472
rect 748 14352 794 14398
rect 748 14245 794 14291
rect 748 14138 794 14184
rect 748 14031 794 14077
rect 748 13924 794 13970
rect 748 13817 794 13863
rect 748 13710 794 13756
rect 748 13602 794 13648
rect 748 13494 794 13540
rect 748 13386 794 13432
rect 748 13278 794 13324
rect 748 13170 794 13216
rect 748 13062 794 13108
rect 972 14352 1018 14398
rect 972 14245 1018 14291
rect 972 14138 1018 14184
rect 972 14031 1018 14077
rect 972 13924 1018 13970
rect 972 13817 1018 13863
rect 972 13710 1018 13756
rect 972 13602 1018 13648
rect 972 13494 1018 13540
rect 972 13386 1018 13432
rect 972 13278 1018 13324
rect 972 13170 1018 13216
rect 972 13062 1018 13108
rect 1196 14352 1242 14398
rect 1196 14245 1242 14291
rect 1196 14138 1242 14184
rect 1196 14031 1242 14077
rect 1196 13924 1242 13970
rect 1196 13817 1242 13863
rect 1196 13710 1242 13756
rect 1196 13602 1242 13648
rect 1196 13494 1242 13540
rect 1196 13386 1242 13432
rect 1196 13278 1242 13324
rect 1196 13170 1242 13216
rect 1196 13062 1242 13108
rect 1420 14352 1466 14398
rect 1420 14245 1466 14291
rect 1420 14138 1466 14184
rect 1420 14031 1466 14077
rect 1420 13924 1466 13970
rect 1420 13817 1466 13863
rect 1420 13710 1466 13756
rect 1420 13602 1466 13648
rect 1420 13494 1466 13540
rect 1420 13386 1466 13432
rect 1420 13278 1466 13324
rect 1420 13170 1466 13216
rect 1420 13062 1466 13108
rect 1644 14322 1690 14368
rect 1644 14217 1690 14263
rect 1644 14112 1690 14158
rect 1644 14007 1690 14053
rect 1644 13902 1690 13948
rect 1644 13797 1690 13843
rect 1644 13692 1690 13738
rect 1644 13587 1690 13633
rect 1644 13482 1690 13528
rect 1644 13377 1690 13423
rect 1644 13272 1690 13318
rect 1644 13167 1690 13213
rect 1644 13062 1690 13108
rect 1868 15258 1914 15304
rect 1868 15154 1914 15200
rect 1868 15050 1914 15096
rect 1868 14946 1914 14992
rect 1868 14842 1914 14888
rect 1868 14738 1914 14784
rect 1868 14634 1914 14680
rect 1868 14530 1914 14576
rect 1868 14426 1914 14472
rect 1868 14322 1914 14368
rect 1868 14217 1914 14263
rect 1868 14112 1914 14158
rect 1868 14007 1914 14053
rect 1868 13902 1914 13948
rect 1868 13797 1914 13843
rect 1868 13692 1914 13738
rect 1868 13587 1914 13633
rect 1868 13482 1914 13528
rect 1868 13377 1914 13423
rect 1868 13272 1914 13318
rect 1868 13167 1914 13213
rect 1868 13062 1914 13108
rect 1629 9374 1675 9420
rect 801 9181 847 9227
rect 801 9025 847 9071
rect 1025 9181 1071 9227
rect 1025 9025 1071 9071
rect 1249 9181 1295 9227
rect 1629 9218 1675 9264
rect 1853 9374 1899 9420
rect 1853 9218 1899 9264
rect 2077 9374 2123 9420
rect 2077 9218 2123 9264
rect 2481 9199 2527 9245
rect 1249 9025 1295 9071
rect 2481 9092 2527 9138
rect 2481 8985 2527 9031
rect 2481 8878 2527 8924
rect 2481 8771 2527 8817
rect 1629 8659 1675 8705
rect 801 8577 847 8623
rect 801 8457 847 8503
rect 1025 8577 1071 8623
rect 1025 8457 1071 8503
rect 1249 8577 1295 8623
rect 1629 8539 1675 8585
rect 1853 8659 1899 8705
rect 1853 8539 1899 8585
rect 2077 8659 2123 8705
rect 2077 8539 2123 8585
rect 2481 8664 2527 8710
rect 2481 8557 2527 8603
rect 1249 8457 1295 8503
rect 2481 8449 2527 8495
rect 2481 8341 2527 8387
rect 2481 8233 2527 8279
rect 2481 8125 2527 8171
rect 2481 8017 2527 8063
rect 2481 7909 2527 7955
rect 2705 9199 2751 9245
rect 2705 9092 2751 9138
rect 2705 8985 2751 9031
rect 2705 8878 2751 8924
rect 2705 8771 2751 8817
rect 2705 8664 2751 8710
rect 2705 8557 2751 8603
rect 2705 8449 2751 8495
rect 2705 8341 2751 8387
rect 2705 8233 2751 8279
rect 2705 8125 2751 8171
rect 2705 8017 2751 8063
rect 2705 7909 2751 7955
<< mvpsubdiff >>
rect 1171 22013 1331 22073
rect 1171 21967 1228 22013
rect 1274 21967 1331 22013
rect 1171 21907 1331 21967
rect 2410 22013 2570 22073
rect 2410 21967 2467 22013
rect 2513 21967 2570 22013
rect 2410 21907 2570 21967
rect 3648 22013 3808 22073
rect 3648 21967 3705 22013
rect 3751 21967 3808 22013
rect 3648 21907 3808 21967
rect 4887 22013 5047 22073
rect 4887 21967 4944 22013
rect 4990 21967 5047 22013
rect 4887 21907 5047 21967
rect 5507 22013 5667 22073
rect 5507 21967 5564 22013
rect 5610 21967 5667 22013
rect 5507 21907 5667 21967
rect 502 17245 586 17264
rect 502 17105 521 17245
rect 567 17105 586 17245
rect 1829 17245 1913 17264
rect 502 17086 586 17105
rect 1829 17105 1848 17245
rect 1894 17105 1913 17245
rect 3068 17245 3152 17264
rect 1829 17086 1913 17105
rect 3068 17105 3087 17245
rect 3133 17105 3152 17245
rect 4306 17245 4390 17264
rect 3068 17086 3152 17105
rect 4306 17105 4325 17245
rect 4371 17105 4390 17245
rect 5545 17245 5629 17264
rect 4306 17086 4390 17105
rect 5545 17105 5564 17245
rect 5610 17105 5629 17245
rect 5545 17086 5629 17105
rect 631 16849 5587 16908
rect 631 16803 754 16849
rect 800 16803 912 16849
rect 958 16803 1070 16849
rect 1116 16803 1228 16849
rect 1274 16803 1386 16849
rect 1432 16803 1544 16849
rect 1590 16803 1702 16849
rect 1748 16803 1993 16849
rect 2039 16803 2151 16849
rect 2197 16803 2309 16849
rect 2355 16803 2467 16849
rect 2513 16803 2625 16849
rect 2671 16803 2783 16849
rect 2829 16803 2941 16849
rect 2987 16803 3231 16849
rect 3277 16803 3389 16849
rect 3435 16803 3547 16849
rect 3593 16803 3705 16849
rect 3751 16803 3863 16849
rect 3909 16803 4021 16849
rect 4067 16803 4179 16849
rect 4225 16803 4470 16849
rect 4516 16803 4628 16849
rect 4674 16803 4786 16849
rect 4832 16803 4944 16849
rect 4990 16803 5102 16849
rect 5148 16803 5260 16849
rect 5306 16803 5418 16849
rect 5464 16803 5587 16849
rect 631 16743 5587 16803
rect 2309 15502 2469 15561
rect 2309 15456 2366 15502
rect 2412 15456 2469 15502
rect 2309 15338 2469 15456
rect 2309 15292 2366 15338
rect 2412 15292 2469 15338
rect 2309 15175 2469 15292
rect 2309 15129 2366 15175
rect 2412 15129 2469 15175
rect 2309 15012 2469 15129
rect 2309 14966 2366 15012
rect 2412 14966 2469 15012
rect 2309 14849 2469 14966
rect 2309 14803 2366 14849
rect 2412 14803 2469 14849
rect 2309 14686 2469 14803
rect 2309 14640 2366 14686
rect 2412 14640 2469 14686
rect 2309 14522 2469 14640
rect 2309 14476 2366 14522
rect 2412 14476 2469 14522
rect 2309 14359 2469 14476
rect 2309 14313 2366 14359
rect 2412 14313 2469 14359
rect 2309 14196 2469 14313
rect 2309 14150 2366 14196
rect 2412 14150 2469 14196
rect 2309 14033 2469 14150
rect 2309 13987 2366 14033
rect 2412 13987 2469 14033
rect 2309 13869 2469 13987
rect 2309 13823 2366 13869
rect 2412 13823 2469 13869
rect 2309 13706 2469 13823
rect 2309 13660 2366 13706
rect 2412 13660 2469 13706
rect 2309 13543 2469 13660
rect 2309 13497 2366 13543
rect 2412 13497 2469 13543
rect 2309 13380 2469 13497
rect 2309 13334 2366 13380
rect 2412 13334 2469 13380
rect 2309 13216 2469 13334
rect 2309 13170 2366 13216
rect 2412 13170 2469 13216
rect 2309 13053 2469 13170
rect 2309 13007 2366 13053
rect 2412 13007 2469 13053
rect 2309 12890 2469 13007
rect 2309 12844 2366 12890
rect 2412 12844 2469 12890
rect 2309 12726 2469 12844
rect 2309 12680 2366 12726
rect 2412 12680 2469 12726
rect 2309 12623 2469 12680
rect 2151 12564 2469 12623
rect 2151 12518 2208 12564
rect 2254 12563 2469 12564
rect 2254 12518 2366 12563
rect 2151 12517 2366 12518
rect 2412 12517 2469 12563
rect 2151 12400 2469 12517
rect 2151 12354 2208 12400
rect 2254 12354 2366 12400
rect 2412 12354 2469 12400
rect 2151 12237 2469 12354
rect 2151 12191 2208 12237
rect 2254 12191 2366 12237
rect 2412 12191 2469 12237
rect 2151 12074 2469 12191
rect 2151 12028 2208 12074
rect 2254 12073 2469 12074
rect 2254 12028 2366 12073
rect 2151 12027 2366 12028
rect 2412 12027 2469 12073
rect 2151 11911 2469 12027
rect 2151 11865 2208 11911
rect 2254 11910 2469 11911
rect 2254 11865 2366 11910
rect 2151 11864 2366 11865
rect 2412 11864 2469 11910
rect 2151 11747 2469 11864
rect 2151 11701 2208 11747
rect 2254 11701 2366 11747
rect 2412 11701 2469 11747
rect 2151 11584 2469 11701
rect 2151 11538 2208 11584
rect 2254 11538 2366 11584
rect 2412 11538 2469 11584
rect 2151 11421 2469 11538
rect 2151 11375 2208 11421
rect 2254 11420 2469 11421
rect 2254 11375 2366 11420
rect 2151 11374 2366 11375
rect 2412 11374 2469 11420
rect 2151 11257 2469 11374
rect 2151 11211 2208 11257
rect 2254 11211 2366 11257
rect 2412 11211 2469 11257
rect 2151 11094 2469 11211
rect 2151 11048 2208 11094
rect 2254 11048 2366 11094
rect 2412 11048 2469 11094
rect 2151 10931 2469 11048
rect 2151 10885 2208 10931
rect 2254 10885 2366 10931
rect 2412 10885 2469 10931
rect 2151 10768 2469 10885
rect 2151 10722 2208 10768
rect 2254 10722 2366 10768
rect 2412 10722 2469 10768
rect 2151 10604 2469 10722
rect 2151 10558 2208 10604
rect 2254 10558 2366 10604
rect 2412 10558 2469 10604
rect 2151 10500 2469 10558
rect 243 9519 403 9579
rect 243 9473 300 9519
rect 346 9473 403 9519
rect 243 9413 403 9473
rect 314 8124 398 8143
rect 314 7984 333 8124
rect 379 7984 398 8124
rect 314 7965 398 7984
<< mvnsubdiff >>
rect 601 28918 5618 28975
rect 601 28872 760 28918
rect 806 28872 918 28918
rect 964 28872 1076 28918
rect 1122 28872 1380 28918
rect 1426 28872 1538 28918
rect 1584 28872 1696 28918
rect 1742 28872 1999 28918
rect 2045 28872 2157 28918
rect 2203 28872 2315 28918
rect 2361 28872 2619 28918
rect 2665 28872 2777 28918
rect 2823 28872 2935 28918
rect 2981 28872 3237 28918
rect 3283 28872 3395 28918
rect 3441 28872 3553 28918
rect 3599 28872 3857 28918
rect 3903 28872 4015 28918
rect 4061 28872 4173 28918
rect 4219 28872 4476 28918
rect 4522 28872 4634 28918
rect 4680 28872 4792 28918
rect 4838 28872 5096 28918
rect 5142 28872 5254 28918
rect 5300 28872 5412 28918
rect 5458 28872 5618 28918
rect 601 28815 5618 28872
rect 1209 24650 1293 24669
rect 1209 24416 1228 24650
rect 1274 24416 1293 24650
rect 1209 24397 1293 24416
rect 2448 24650 2532 24669
rect 2448 24416 2467 24650
rect 2513 24416 2532 24650
rect 2448 24397 2532 24416
rect 3686 24650 3770 24669
rect 3686 24416 3705 24650
rect 3751 24416 3770 24650
rect 3686 24397 3770 24416
rect 4925 24650 5009 24669
rect 4925 24416 4944 24650
rect 4990 24416 5009 24650
rect 4925 24397 5009 24416
rect 631 18168 5587 18225
rect 631 18122 754 18168
rect 800 18122 912 18168
rect 958 18122 1070 18168
rect 1116 18122 1228 18168
rect 1274 18122 1386 18168
rect 1432 18122 1544 18168
rect 1590 18122 1702 18168
rect 1748 18122 1993 18168
rect 2039 18122 2151 18168
rect 2197 18122 2309 18168
rect 2355 18122 2467 18168
rect 2513 18122 2625 18168
rect 2671 18122 2783 18168
rect 2829 18122 2941 18168
rect 2987 18122 3231 18168
rect 3277 18122 3389 18168
rect 3435 18122 3547 18168
rect 3593 18122 3705 18168
rect 3751 18122 3863 18168
rect 3909 18122 4021 18168
rect 4067 18122 4179 18168
rect 4225 18122 4470 18168
rect 4516 18122 4628 18168
rect 4674 18122 4786 18168
rect 4832 18122 4944 18168
rect 4990 18122 5102 18168
rect 5148 18122 5260 18168
rect 5306 18122 5418 18168
rect 5464 18122 5587 18168
rect 631 18065 5587 18122
rect 1646 15555 1918 15574
rect 1646 15509 1665 15555
rect 1899 15509 1918 15555
rect 1646 15490 1918 15509
rect 245 8971 401 9028
rect 245 8925 300 8971
rect 346 8925 401 8971
rect 245 8807 401 8925
rect 245 8761 300 8807
rect 346 8761 401 8807
rect 245 8704 401 8761
<< mvpsubdiffcont >>
rect 1228 21967 1274 22013
rect 2467 21967 2513 22013
rect 3705 21967 3751 22013
rect 4944 21967 4990 22013
rect 5564 21967 5610 22013
rect 521 17105 567 17245
rect 1848 17105 1894 17245
rect 3087 17105 3133 17245
rect 4325 17105 4371 17245
rect 5564 17105 5610 17245
rect 754 16803 800 16849
rect 912 16803 958 16849
rect 1070 16803 1116 16849
rect 1228 16803 1274 16849
rect 1386 16803 1432 16849
rect 1544 16803 1590 16849
rect 1702 16803 1748 16849
rect 1993 16803 2039 16849
rect 2151 16803 2197 16849
rect 2309 16803 2355 16849
rect 2467 16803 2513 16849
rect 2625 16803 2671 16849
rect 2783 16803 2829 16849
rect 2941 16803 2987 16849
rect 3231 16803 3277 16849
rect 3389 16803 3435 16849
rect 3547 16803 3593 16849
rect 3705 16803 3751 16849
rect 3863 16803 3909 16849
rect 4021 16803 4067 16849
rect 4179 16803 4225 16849
rect 4470 16803 4516 16849
rect 4628 16803 4674 16849
rect 4786 16803 4832 16849
rect 4944 16803 4990 16849
rect 5102 16803 5148 16849
rect 5260 16803 5306 16849
rect 5418 16803 5464 16849
rect 2366 15456 2412 15502
rect 2366 15292 2412 15338
rect 2366 15129 2412 15175
rect 2366 14966 2412 15012
rect 2366 14803 2412 14849
rect 2366 14640 2412 14686
rect 2366 14476 2412 14522
rect 2366 14313 2412 14359
rect 2366 14150 2412 14196
rect 2366 13987 2412 14033
rect 2366 13823 2412 13869
rect 2366 13660 2412 13706
rect 2366 13497 2412 13543
rect 2366 13334 2412 13380
rect 2366 13170 2412 13216
rect 2366 13007 2412 13053
rect 2366 12844 2412 12890
rect 2366 12680 2412 12726
rect 2208 12518 2254 12564
rect 2366 12517 2412 12563
rect 2208 12354 2254 12400
rect 2366 12354 2412 12400
rect 2208 12191 2254 12237
rect 2366 12191 2412 12237
rect 2208 12028 2254 12074
rect 2366 12027 2412 12073
rect 2208 11865 2254 11911
rect 2366 11864 2412 11910
rect 2208 11701 2254 11747
rect 2366 11701 2412 11747
rect 2208 11538 2254 11584
rect 2366 11538 2412 11584
rect 2208 11375 2254 11421
rect 2366 11374 2412 11420
rect 2208 11211 2254 11257
rect 2366 11211 2412 11257
rect 2208 11048 2254 11094
rect 2366 11048 2412 11094
rect 2208 10885 2254 10931
rect 2366 10885 2412 10931
rect 2208 10722 2254 10768
rect 2366 10722 2412 10768
rect 2208 10558 2254 10604
rect 2366 10558 2412 10604
rect 300 9473 346 9519
rect 333 7984 379 8124
<< mvnsubdiffcont >>
rect 760 28872 806 28918
rect 918 28872 964 28918
rect 1076 28872 1122 28918
rect 1380 28872 1426 28918
rect 1538 28872 1584 28918
rect 1696 28872 1742 28918
rect 1999 28872 2045 28918
rect 2157 28872 2203 28918
rect 2315 28872 2361 28918
rect 2619 28872 2665 28918
rect 2777 28872 2823 28918
rect 2935 28872 2981 28918
rect 3237 28872 3283 28918
rect 3395 28872 3441 28918
rect 3553 28872 3599 28918
rect 3857 28872 3903 28918
rect 4015 28872 4061 28918
rect 4173 28872 4219 28918
rect 4476 28872 4522 28918
rect 4634 28872 4680 28918
rect 4792 28872 4838 28918
rect 5096 28872 5142 28918
rect 5254 28872 5300 28918
rect 5412 28872 5458 28918
rect 1228 24416 1274 24650
rect 2467 24416 2513 24650
rect 3705 24416 3751 24650
rect 4944 24416 4990 24650
rect 754 18122 800 18168
rect 912 18122 958 18168
rect 1070 18122 1116 18168
rect 1228 18122 1274 18168
rect 1386 18122 1432 18168
rect 1544 18122 1590 18168
rect 1702 18122 1748 18168
rect 1993 18122 2039 18168
rect 2151 18122 2197 18168
rect 2309 18122 2355 18168
rect 2467 18122 2513 18168
rect 2625 18122 2671 18168
rect 2783 18122 2829 18168
rect 2941 18122 2987 18168
rect 3231 18122 3277 18168
rect 3389 18122 3435 18168
rect 3547 18122 3593 18168
rect 3705 18122 3751 18168
rect 3863 18122 3909 18168
rect 4021 18122 4067 18168
rect 4179 18122 4225 18168
rect 4470 18122 4516 18168
rect 4628 18122 4674 18168
rect 4786 18122 4832 18168
rect 4944 18122 4990 18168
rect 5102 18122 5148 18168
rect 5260 18122 5306 18168
rect 5418 18122 5464 18168
rect 1665 15509 1899 15555
rect 300 8925 346 8971
rect 300 8761 346 8807
<< polysilicon >>
rect 769 28626 889 28699
rect 993 28626 1113 28699
rect 1389 28626 1509 28699
rect 1613 28626 1733 28699
rect 2008 28626 2128 28699
rect 2232 28626 2352 28699
rect 2628 28626 2748 28699
rect 2852 28626 2972 28699
rect 3246 28626 3366 28699
rect 3470 28626 3590 28699
rect 3866 28626 3986 28699
rect 4090 28626 4210 28699
rect 4485 28626 4605 28699
rect 4709 28626 4829 28699
rect 5069 28626 5189 28699
rect 5294 28626 5414 28699
rect 769 27851 889 27944
rect 993 27851 1113 27944
rect 1389 27851 1509 27944
rect 1613 27851 1733 27944
rect 2008 27851 2128 27944
rect 2232 27851 2352 27944
rect 2628 27851 2748 27944
rect 2852 27851 2972 27944
rect 3246 27851 3366 27944
rect 3470 27851 3590 27944
rect 3866 27851 3986 27944
rect 4090 27851 4210 27944
rect 4485 27851 4605 27944
rect 4709 27851 4829 27944
rect 5069 27851 5189 27944
rect 5294 27851 5414 27944
rect 769 27105 889 27169
rect 993 27105 1113 27169
rect 769 27086 1113 27105
rect 769 27040 847 27086
rect 1081 27040 1113 27086
rect 769 27021 1113 27040
rect 1389 27105 1509 27169
rect 1613 27105 1733 27169
rect 1389 27086 1733 27105
rect 1389 27040 1421 27086
rect 1655 27040 1733 27086
rect 1389 27021 1733 27040
rect 2008 27105 2128 27169
rect 2232 27105 2352 27169
rect 2008 27086 2352 27105
rect 2008 27040 2086 27086
rect 2320 27040 2352 27086
rect 2008 27021 2352 27040
rect 2628 27105 2748 27169
rect 2852 27105 2972 27169
rect 2628 27086 2972 27105
rect 2628 27040 2660 27086
rect 2894 27040 2972 27086
rect 2628 27021 2972 27040
rect 3246 27105 3366 27169
rect 3470 27105 3590 27169
rect 3246 27086 3590 27105
rect 3246 27040 3324 27086
rect 3558 27040 3590 27086
rect 3246 27021 3590 27040
rect 3866 27105 3986 27169
rect 4090 27105 4210 27169
rect 3866 27086 4210 27105
rect 3866 27040 3898 27086
rect 4132 27040 4210 27086
rect 3866 27021 4210 27040
rect 4485 27105 4605 27169
rect 4709 27105 4829 27169
rect 4485 27086 4829 27105
rect 4485 27040 4563 27086
rect 4797 27040 4829 27086
rect 4485 27021 4829 27040
rect 5069 27101 5189 27169
rect 5294 27101 5414 27169
rect 5069 27082 5414 27101
rect 5069 27036 5122 27082
rect 5356 27036 5414 27082
rect 883 26950 1003 27021
rect 1499 26950 1619 27021
rect 2122 26950 2242 27021
rect 2738 26950 2858 27021
rect 3360 26950 3480 27021
rect 3976 26950 4096 27021
rect 4599 26950 4719 27021
rect 5069 27017 5414 27036
rect 5215 26950 5335 27017
rect 883 25517 1003 25588
rect 1499 25517 1619 25588
rect 2122 25517 2242 25588
rect 2738 25517 2858 25588
rect 3360 25517 3480 25588
rect 3976 25517 4096 25588
rect 4599 25517 4719 25588
rect 5215 25517 5335 25588
rect 881 25363 1001 25437
rect 1501 25363 1621 25437
rect 2120 25363 2240 25437
rect 2740 25363 2860 25437
rect 3358 25363 3478 25437
rect 3978 25363 4098 25437
rect 4597 25363 4717 25437
rect 5217 25363 5337 25437
rect 881 23917 1001 24001
rect 881 23871 912 23917
rect 958 23871 1001 23917
rect 881 23852 1001 23871
rect 1501 23917 1621 24001
rect 1501 23871 1544 23917
rect 1590 23871 1621 23917
rect 1501 23852 1621 23871
rect 2120 23917 2240 24001
rect 2120 23871 2151 23917
rect 2197 23871 2240 23917
rect 2120 23852 2240 23871
rect 2740 23917 2860 24001
rect 2740 23871 2783 23917
rect 2829 23871 2860 23917
rect 2740 23852 2860 23871
rect 3358 23917 3478 24001
rect 3358 23871 3389 23917
rect 3435 23871 3478 23917
rect 3358 23852 3478 23871
rect 3978 23917 4098 24001
rect 3978 23871 4021 23917
rect 4067 23871 4098 23917
rect 3978 23852 4098 23871
rect 4597 23917 4717 24001
rect 4597 23871 4628 23917
rect 4674 23871 4717 23917
rect 4597 23852 4717 23871
rect 5217 23917 5337 24001
rect 5217 23871 5260 23917
rect 5306 23871 5337 23917
rect 5217 23852 5337 23871
rect 881 23672 1001 23746
rect 1501 23672 1621 23746
rect 2120 23672 2240 23746
rect 2740 23672 2860 23746
rect 3358 23672 3478 23746
rect 3978 23672 4098 23746
rect 4597 23672 4717 23746
rect 5217 23672 5337 23746
rect 881 22238 1001 22310
rect 882 21742 1001 22238
rect 1501 22238 1621 22310
rect 2120 22238 2240 22310
rect 881 21668 1001 21742
rect 1501 21742 1620 22238
rect 2121 21742 2240 22238
rect 2740 22238 2860 22310
rect 3358 22238 3478 22310
rect 1501 21668 1621 21742
rect 2120 21668 2240 21742
rect 2740 21742 2859 22238
rect 3359 21742 3478 22238
rect 3978 22238 4098 22310
rect 4597 22238 4717 22310
rect 2740 21668 2860 21742
rect 3358 21668 3478 21742
rect 3978 21742 4097 22238
rect 4598 21742 4717 22238
rect 3978 21668 4098 21742
rect 4597 21668 4717 21742
rect 5217 21668 5337 22310
rect 881 20222 1001 20306
rect 881 20176 918 20222
rect 964 20176 1001 20222
rect 881 20157 1001 20176
rect 1501 20222 1621 20306
rect 1501 20176 1538 20222
rect 1584 20176 1621 20222
rect 1501 20157 1621 20176
rect 2120 20222 2240 20306
rect 2120 20176 2157 20222
rect 2203 20176 2240 20222
rect 2120 20157 2240 20176
rect 2740 20222 2860 20306
rect 2740 20176 2777 20222
rect 2823 20176 2860 20222
rect 2740 20157 2860 20176
rect 3358 20222 3478 20306
rect 3358 20176 3395 20222
rect 3441 20176 3478 20222
rect 3358 20157 3478 20176
rect 3978 20222 4098 20306
rect 3978 20176 4015 20222
rect 4061 20176 4098 20222
rect 3978 20157 4098 20176
rect 4597 20222 4717 20306
rect 4597 20176 4634 20222
rect 4680 20176 4717 20222
rect 4597 20157 4717 20176
rect 5217 20222 5337 20306
rect 5217 20176 5254 20222
rect 5300 20176 5337 20222
rect 5217 20157 5337 20176
rect 881 19945 1001 19964
rect 881 19899 918 19945
rect 964 19899 1001 19945
rect 881 19813 1001 19899
rect 1501 19945 1621 19964
rect 1501 19899 1538 19945
rect 1584 19899 1621 19945
rect 1501 19813 1621 19899
rect 2120 19945 2240 19964
rect 2120 19899 2157 19945
rect 2203 19899 2240 19945
rect 2120 19813 2240 19899
rect 2740 19945 2860 19964
rect 2740 19899 2777 19945
rect 2823 19899 2860 19945
rect 2740 19813 2860 19899
rect 3358 19945 3478 19964
rect 3358 19899 3395 19945
rect 3441 19899 3478 19945
rect 3358 19813 3478 19899
rect 3978 19945 4098 19964
rect 3978 19899 4015 19945
rect 4061 19899 4098 19945
rect 3978 19813 4098 19899
rect 4597 19945 4717 19964
rect 4597 19899 4634 19945
rect 4680 19899 4717 19945
rect 4597 19813 4717 19899
rect 5217 19945 5337 19964
rect 5217 19899 5254 19945
rect 5300 19899 5337 19945
rect 5217 19813 5337 19899
rect 881 18380 1001 18451
rect 1501 18380 1621 18451
rect 2120 18380 2240 18451
rect 2740 18380 2860 18451
rect 3358 18380 3478 18451
rect 3978 18380 4098 18451
rect 4597 18380 4717 18451
rect 5217 18380 5337 18451
rect 812 17978 1184 17997
rect 812 17932 975 17978
rect 1021 17932 1184 17978
rect 812 17898 1184 17932
rect 812 17838 932 17898
rect 1064 17838 1184 17898
rect 1318 17978 1690 17997
rect 1318 17932 1481 17978
rect 1527 17932 1690 17978
rect 1318 17898 1690 17932
rect 1318 17838 1438 17898
rect 1570 17838 1690 17898
rect 2051 17978 2423 17997
rect 2051 17932 2214 17978
rect 2260 17932 2423 17978
rect 2051 17898 2423 17932
rect 2051 17838 2171 17898
rect 2303 17838 2423 17898
rect 2557 17978 2929 17997
rect 2557 17932 2720 17978
rect 2766 17932 2929 17978
rect 2557 17898 2929 17932
rect 2557 17838 2677 17898
rect 2809 17838 2929 17898
rect 3289 17978 3661 17997
rect 3289 17932 3452 17978
rect 3498 17932 3661 17978
rect 3289 17898 3661 17932
rect 3289 17838 3409 17898
rect 3541 17838 3661 17898
rect 3795 17978 4167 17997
rect 3795 17932 3958 17978
rect 4004 17932 4167 17978
rect 3795 17898 4167 17932
rect 3795 17838 3915 17898
rect 4047 17838 4167 17898
rect 4528 17978 4900 17997
rect 4528 17932 4691 17978
rect 4737 17932 4900 17978
rect 4528 17898 4900 17932
rect 4528 17838 4648 17898
rect 4780 17838 4900 17898
rect 5034 17978 5405 17997
rect 5034 17932 5197 17978
rect 5243 17932 5405 17978
rect 5034 17898 5405 17932
rect 5034 17838 5154 17898
rect 5285 17838 5405 17898
rect 812 17354 932 17541
rect 1064 17414 1184 17541
rect 855 17323 932 17354
rect 1079 17365 1184 17414
rect 1318 17414 1438 17541
rect 1318 17365 1423 17414
rect 855 17250 975 17323
rect 1079 17250 1199 17365
rect 1303 17250 1423 17365
rect 1570 17354 1690 17541
rect 2051 17354 2171 17541
rect 2303 17414 2423 17541
rect 1570 17323 1647 17354
rect 1527 17250 1647 17323
rect 2094 17323 2171 17354
rect 2318 17365 2423 17414
rect 2557 17414 2677 17541
rect 2557 17365 2662 17414
rect 2094 17250 2214 17323
rect 2318 17250 2438 17365
rect 2542 17250 2662 17365
rect 2809 17354 2929 17541
rect 3289 17354 3409 17541
rect 3541 17414 3661 17541
rect 2809 17323 2886 17354
rect 2766 17250 2886 17323
rect 3332 17323 3409 17354
rect 3556 17365 3661 17414
rect 3795 17414 3915 17541
rect 3795 17365 3900 17414
rect 855 17063 975 17136
rect 1079 17063 1199 17136
rect 1303 17063 1423 17136
rect 1527 17063 1647 17136
rect 3332 17250 3452 17323
rect 3556 17250 3676 17365
rect 3780 17250 3900 17365
rect 4047 17354 4167 17541
rect 4528 17354 4648 17541
rect 4780 17414 4900 17541
rect 4047 17323 4124 17354
rect 4004 17250 4124 17323
rect 4571 17323 4648 17354
rect 4795 17365 4900 17414
rect 5034 17388 5154 17541
rect 5285 17389 5405 17541
rect 2094 17063 2214 17136
rect 2318 17063 2438 17136
rect 2542 17063 2662 17136
rect 2766 17063 2886 17136
rect 4571 17250 4691 17323
rect 4795 17250 4915 17365
rect 5019 17351 5154 17388
rect 5243 17355 5405 17389
rect 5019 17250 5139 17351
rect 5243 17250 5363 17355
rect 3332 17063 3452 17136
rect 3556 17063 3676 17136
rect 3780 17063 3900 17136
rect 4004 17063 4124 17136
rect 4571 17063 4691 17136
rect 4795 17063 4915 17136
rect 5019 17063 5139 17136
rect 5243 17063 5363 17136
rect 375 15815 494 15843
rect 375 15771 495 15815
rect 1043 15697 1163 15770
rect 1043 15407 1163 15469
rect 916 15400 1163 15407
rect 916 15361 1321 15400
rect 916 15315 990 15361
rect 1036 15315 1321 15361
rect 1719 15317 1839 15361
rect 916 15270 1321 15315
rect 928 15260 1321 15270
rect 928 15190 1048 15260
rect 1201 15190 1321 15260
rect 928 14821 1048 14893
rect 1201 14821 1321 14893
rect 1034 14695 1228 14741
rect 1034 14649 1108 14695
rect 1154 14649 1228 14695
rect 1034 14531 1228 14649
rect 823 14471 1391 14531
rect 823 14411 943 14471
rect 1271 14411 1391 14471
rect 375 12613 495 13049
rect 823 12975 943 13049
rect 1271 12975 1391 13049
rect 1719 12898 1839 13049
rect 1574 12897 1839 12898
rect 1443 12852 1839 12897
rect 1443 12806 1516 12852
rect 1562 12806 1839 12852
rect 1443 12761 1839 12806
rect 1574 12760 1839 12761
rect 823 12612 943 12685
rect 1271 12612 1391 12685
rect 1719 12612 1839 12760
rect 823 10284 943 10344
rect 1271 10284 1391 10344
rect 823 10258 1391 10284
rect 1719 10271 1839 10344
rect 823 10212 976 10258
rect 1022 10212 1391 10258
rect 823 10193 1391 10212
rect 1704 10045 1824 10064
rect 1704 9999 1741 10045
rect 1787 9999 1824 10045
rect 1704 9904 1824 9999
rect 2556 9990 2676 10034
rect 375 9818 495 9891
rect 339 9773 531 9818
rect 986 9804 1106 9876
rect 339 9727 412 9773
rect 458 9727 531 9773
rect 339 9682 531 9727
rect 1704 9629 1824 9712
rect 986 9354 1106 9612
rect 1704 9569 2048 9629
rect 1704 9433 1824 9569
rect 1928 9433 2048 9569
rect 876 9300 1220 9354
rect 876 9240 996 9300
rect 1100 9240 1220 9300
rect 2556 9258 2676 9536
rect 1704 9133 1824 9205
rect 1928 9133 2048 9205
rect 1371 9020 1563 9065
rect 876 8925 996 9012
rect 1100 8940 1220 9012
rect 1371 8974 1444 9020
rect 1490 8989 1563 9020
rect 1490 8974 2048 8989
rect 1371 8929 2048 8974
rect 1927 8928 2048 8929
rect 802 8880 996 8925
rect 802 8834 875 8880
rect 921 8849 996 8880
rect 921 8834 1824 8849
rect 802 8789 1824 8834
rect 876 8788 1824 8789
rect 1704 8718 1824 8788
rect 1928 8718 2048 8928
rect 876 8636 996 8680
rect 1100 8636 1220 8680
rect 599 8334 793 8373
rect 876 8334 996 8444
rect 1100 8372 1220 8444
rect 1704 8373 1824 8526
rect 1928 8453 2048 8526
rect 599 8327 996 8334
rect 599 8281 673 8327
rect 719 8281 996 8327
rect 599 8274 996 8281
rect 599 8236 793 8274
rect 611 8235 793 8236
rect 876 8163 996 8274
rect 1044 8327 1236 8372
rect 1044 8281 1117 8327
rect 1163 8281 1236 8327
rect 1704 8312 2048 8373
rect 1044 8236 1236 8281
rect 1425 8262 1509 8271
rect 1425 8252 1824 8262
rect 1100 8163 1220 8236
rect 1425 8206 1444 8252
rect 1490 8206 1824 8252
rect 1425 8202 1824 8206
rect 1425 8187 1509 8202
rect 1704 8142 1824 8202
rect 1928 8142 2048 8312
rect 876 7927 996 7971
rect 1100 7927 1220 7971
rect 1704 7906 1824 7950
rect 1928 7906 2048 7950
rect 2556 7813 2676 7896
rect 2556 7767 2593 7813
rect 2639 7767 2676 7813
rect 2556 7748 2676 7767
<< polycontact >>
rect 847 27040 1081 27086
rect 1421 27040 1655 27086
rect 2086 27040 2320 27086
rect 2660 27040 2894 27086
rect 3324 27040 3558 27086
rect 3898 27040 4132 27086
rect 4563 27040 4797 27086
rect 5122 27036 5356 27082
rect 912 23871 958 23917
rect 1544 23871 1590 23917
rect 2151 23871 2197 23917
rect 2783 23871 2829 23917
rect 3389 23871 3435 23917
rect 4021 23871 4067 23917
rect 4628 23871 4674 23917
rect 5260 23871 5306 23917
rect 918 20176 964 20222
rect 1538 20176 1584 20222
rect 2157 20176 2203 20222
rect 2777 20176 2823 20222
rect 3395 20176 3441 20222
rect 4015 20176 4061 20222
rect 4634 20176 4680 20222
rect 5254 20176 5300 20222
rect 918 19899 964 19945
rect 1538 19899 1584 19945
rect 2157 19899 2203 19945
rect 2777 19899 2823 19945
rect 3395 19899 3441 19945
rect 4015 19899 4061 19945
rect 4634 19899 4680 19945
rect 5254 19899 5300 19945
rect 975 17932 1021 17978
rect 1481 17932 1527 17978
rect 2214 17932 2260 17978
rect 2720 17932 2766 17978
rect 3452 17932 3498 17978
rect 3958 17932 4004 17978
rect 4691 17932 4737 17978
rect 5197 17932 5243 17978
rect 990 15315 1036 15361
rect 1108 14649 1154 14695
rect 1516 12806 1562 12852
rect 976 10212 1022 10258
rect 1741 9999 1787 10045
rect 412 9727 458 9773
rect 1444 8974 1490 9020
rect 875 8834 921 8880
rect 673 8281 719 8327
rect 1117 8281 1163 8327
rect 1444 8206 1490 8252
rect 2593 7767 2639 7813
<< metal1 >>
rect 631 28956 5587 28980
rect 631 28918 918 28956
rect 970 28918 1532 28956
rect 1584 28918 2157 28956
rect 2209 28918 2771 28956
rect 2823 28918 3395 28956
rect 3447 28918 4009 28956
rect 4061 28918 4634 28956
rect 4686 28918 5248 28956
rect 5300 28918 5587 28956
rect 631 28872 760 28918
rect 806 28872 918 28918
rect 970 28904 1076 28918
rect 964 28872 1076 28904
rect 1122 28872 1380 28918
rect 1426 28904 1532 28918
rect 1426 28872 1538 28904
rect 1584 28872 1696 28918
rect 1742 28872 1999 28918
rect 2045 28872 2157 28918
rect 2209 28904 2315 28918
rect 2203 28872 2315 28904
rect 2361 28872 2619 28918
rect 2665 28904 2771 28918
rect 2665 28872 2777 28904
rect 2823 28872 2935 28918
rect 2981 28872 3237 28918
rect 3283 28872 3395 28918
rect 3447 28904 3553 28918
rect 3441 28872 3553 28904
rect 3599 28872 3857 28918
rect 3903 28904 4009 28918
rect 3903 28872 4015 28904
rect 4061 28872 4173 28918
rect 4219 28872 4476 28918
rect 4522 28872 4634 28918
rect 4686 28904 4792 28918
rect 4680 28872 4792 28904
rect 4838 28872 5096 28918
rect 5142 28904 5248 28918
rect 5142 28872 5254 28904
rect 5300 28872 5412 28918
rect 5458 28872 5587 28918
rect 631 28770 5587 28872
rect 631 28718 918 28770
rect 970 28718 1532 28770
rect 1584 28718 2157 28770
rect 2209 28718 2771 28770
rect 2823 28718 3395 28770
rect 3447 28718 4009 28770
rect 4061 28718 4634 28770
rect 4686 28718 5248 28770
rect 5300 28718 5587 28770
rect 631 28697 5587 28718
rect 631 28581 779 28697
rect 631 28535 692 28581
rect 738 28535 779 28581
rect 631 28399 779 28535
rect 631 28353 692 28399
rect 738 28353 779 28399
rect 631 28218 779 28353
rect 631 28172 692 28218
rect 738 28172 779 28218
rect 631 28036 779 28172
rect 631 27990 692 28036
rect 738 27990 779 28036
rect 631 27805 779 27990
rect 884 28581 999 28617
rect 884 28535 918 28581
rect 964 28535 999 28581
rect 884 28399 999 28535
rect 884 28386 918 28399
rect 964 28386 999 28399
rect 884 28230 914 28386
rect 966 28230 999 28386
rect 884 28218 999 28230
rect 884 28172 918 28218
rect 964 28172 999 28218
rect 884 28036 999 28172
rect 884 27990 918 28036
rect 964 27990 999 28036
rect 884 27953 999 27990
rect 1104 28581 1398 28697
rect 1104 28535 1228 28581
rect 1274 28535 1398 28581
rect 1104 28399 1398 28535
rect 1104 28353 1228 28399
rect 1274 28353 1398 28399
rect 1104 28218 1398 28353
rect 1104 28172 1228 28218
rect 1274 28172 1398 28218
rect 1104 28036 1398 28172
rect 1104 27990 1228 28036
rect 1274 27990 1398 28036
rect 631 27759 692 27805
rect 738 27759 779 27805
rect 631 27624 779 27759
rect 631 27578 692 27624
rect 738 27578 779 27624
rect 631 27443 779 27578
rect 631 27397 692 27443
rect 738 27397 779 27443
rect 631 27261 779 27397
rect 631 27215 692 27261
rect 738 27215 779 27261
rect 631 27178 779 27215
rect 884 27805 999 27842
rect 884 27759 918 27805
rect 964 27759 999 27805
rect 884 27624 999 27759
rect 884 27611 918 27624
rect 964 27611 999 27624
rect 884 27455 914 27611
rect 966 27455 999 27611
rect 884 27443 999 27455
rect 884 27397 918 27443
rect 964 27397 999 27443
rect 884 27261 999 27397
rect 884 27215 918 27261
rect 964 27215 999 27261
rect 884 27178 999 27215
rect 1104 27805 1398 27990
rect 1503 28581 1618 28617
rect 1503 28535 1538 28581
rect 1584 28535 1618 28581
rect 1503 28399 1618 28535
rect 1503 28386 1538 28399
rect 1584 28386 1618 28399
rect 1503 28230 1536 28386
rect 1588 28230 1618 28386
rect 1503 28218 1618 28230
rect 1503 28172 1538 28218
rect 1584 28172 1618 28218
rect 1503 28036 1618 28172
rect 1503 27990 1538 28036
rect 1584 27990 1618 28036
rect 1503 27953 1618 27990
rect 1723 28581 2018 28697
rect 1723 28535 1764 28581
rect 1810 28535 1931 28581
rect 1977 28535 2018 28581
rect 1723 28399 2018 28535
rect 1723 28353 1764 28399
rect 1810 28353 1931 28399
rect 1977 28353 2018 28399
rect 1723 28218 2018 28353
rect 1723 28172 1764 28218
rect 1810 28172 1931 28218
rect 1977 28172 2018 28218
rect 1723 28036 2018 28172
rect 1723 27990 1764 28036
rect 1810 27990 1931 28036
rect 1977 27990 2018 28036
rect 1104 27759 1228 27805
rect 1274 27759 1398 27805
rect 1104 27624 1398 27759
rect 1104 27578 1228 27624
rect 1274 27578 1398 27624
rect 1104 27443 1398 27578
rect 1104 27397 1228 27443
rect 1274 27397 1398 27443
rect 1104 27261 1398 27397
rect 1104 27215 1228 27261
rect 1274 27215 1398 27261
rect 1104 27178 1398 27215
rect 1503 27805 1618 27842
rect 1503 27759 1538 27805
rect 1584 27759 1618 27805
rect 1503 27624 1618 27759
rect 1503 27611 1538 27624
rect 1584 27611 1618 27624
rect 1503 27455 1536 27611
rect 1588 27455 1618 27611
rect 1503 27443 1618 27455
rect 1503 27397 1538 27443
rect 1584 27397 1618 27443
rect 1503 27261 1618 27397
rect 1503 27215 1538 27261
rect 1584 27215 1618 27261
rect 1503 27178 1618 27215
rect 1723 27805 2018 27990
rect 2123 28581 2238 28617
rect 2123 28535 2157 28581
rect 2203 28535 2238 28581
rect 2123 28399 2238 28535
rect 2123 28386 2157 28399
rect 2203 28386 2238 28399
rect 2123 28230 2153 28386
rect 2205 28230 2238 28386
rect 2123 28218 2238 28230
rect 2123 28172 2157 28218
rect 2203 28172 2238 28218
rect 2123 28036 2238 28172
rect 2123 27990 2157 28036
rect 2203 27990 2238 28036
rect 2123 27953 2238 27990
rect 2343 28581 2637 28697
rect 2343 28535 2467 28581
rect 2513 28535 2637 28581
rect 2343 28399 2637 28535
rect 2343 28353 2467 28399
rect 2513 28353 2637 28399
rect 2343 28218 2637 28353
rect 2343 28172 2467 28218
rect 2513 28172 2637 28218
rect 2343 28036 2637 28172
rect 2343 27990 2467 28036
rect 2513 27990 2637 28036
rect 1723 27759 1764 27805
rect 1810 27759 1931 27805
rect 1977 27759 2018 27805
rect 1723 27624 2018 27759
rect 1723 27578 1764 27624
rect 1810 27578 1931 27624
rect 1977 27578 2018 27624
rect 1723 27443 2018 27578
rect 1723 27397 1764 27443
rect 1810 27397 1931 27443
rect 1977 27397 2018 27443
rect 1723 27261 2018 27397
rect 1723 27215 1764 27261
rect 1810 27215 1931 27261
rect 1977 27215 2018 27261
rect 1723 27178 2018 27215
rect 2123 27805 2238 27842
rect 2123 27759 2157 27805
rect 2203 27759 2238 27805
rect 2123 27624 2238 27759
rect 2123 27611 2157 27624
rect 2203 27611 2238 27624
rect 2123 27455 2153 27611
rect 2205 27455 2238 27611
rect 2123 27443 2238 27455
rect 2123 27397 2157 27443
rect 2203 27397 2238 27443
rect 2123 27261 2238 27397
rect 2123 27215 2157 27261
rect 2203 27215 2238 27261
rect 2123 27178 2238 27215
rect 2343 27805 2637 27990
rect 2742 28581 2857 28617
rect 2742 28535 2777 28581
rect 2823 28535 2857 28581
rect 2742 28399 2857 28535
rect 2742 28386 2777 28399
rect 2823 28386 2857 28399
rect 2742 28230 2775 28386
rect 2827 28230 2857 28386
rect 2742 28218 2857 28230
rect 2742 28172 2777 28218
rect 2823 28172 2857 28218
rect 2742 28036 2857 28172
rect 2742 27990 2777 28036
rect 2823 27990 2857 28036
rect 2742 27953 2857 27990
rect 2962 28581 3256 28697
rect 2962 28535 3003 28581
rect 3049 28535 3169 28581
rect 3215 28535 3256 28581
rect 2962 28399 3256 28535
rect 2962 28353 3003 28399
rect 3049 28353 3169 28399
rect 3215 28353 3256 28399
rect 2962 28218 3256 28353
rect 2962 28172 3003 28218
rect 3049 28172 3169 28218
rect 3215 28172 3256 28218
rect 2962 28036 3256 28172
rect 2962 27990 3003 28036
rect 3049 27990 3169 28036
rect 3215 27990 3256 28036
rect 2343 27759 2467 27805
rect 2513 27759 2637 27805
rect 2343 27624 2637 27759
rect 2343 27578 2467 27624
rect 2513 27578 2637 27624
rect 2343 27443 2637 27578
rect 2343 27397 2467 27443
rect 2513 27397 2637 27443
rect 2343 27261 2637 27397
rect 2343 27215 2467 27261
rect 2513 27215 2637 27261
rect 2343 27178 2637 27215
rect 2742 27805 2857 27842
rect 2742 27759 2777 27805
rect 2823 27759 2857 27805
rect 2742 27624 2857 27759
rect 2742 27611 2777 27624
rect 2823 27611 2857 27624
rect 2742 27455 2775 27611
rect 2827 27455 2857 27611
rect 2742 27443 2857 27455
rect 2742 27397 2777 27443
rect 2823 27397 2857 27443
rect 2742 27261 2857 27397
rect 2742 27215 2777 27261
rect 2823 27215 2857 27261
rect 2742 27178 2857 27215
rect 2962 27805 3256 27990
rect 3361 28581 3476 28617
rect 3361 28535 3395 28581
rect 3441 28535 3476 28581
rect 3361 28399 3476 28535
rect 3361 28386 3395 28399
rect 3441 28386 3476 28399
rect 3361 28230 3391 28386
rect 3443 28230 3476 28386
rect 3361 28218 3476 28230
rect 3361 28172 3395 28218
rect 3441 28172 3476 28218
rect 3361 28036 3476 28172
rect 3361 27990 3395 28036
rect 3441 27990 3476 28036
rect 3361 27953 3476 27990
rect 3581 28581 3875 28697
rect 3581 28535 3705 28581
rect 3751 28535 3875 28581
rect 3581 28399 3875 28535
rect 3581 28353 3705 28399
rect 3751 28353 3875 28399
rect 3581 28218 3875 28353
rect 3581 28172 3705 28218
rect 3751 28172 3875 28218
rect 3581 28036 3875 28172
rect 3581 27990 3705 28036
rect 3751 27990 3875 28036
rect 2962 27759 3003 27805
rect 3049 27759 3169 27805
rect 3215 27759 3256 27805
rect 2962 27624 3256 27759
rect 2962 27578 3003 27624
rect 3049 27578 3169 27624
rect 3215 27578 3256 27624
rect 2962 27443 3256 27578
rect 2962 27397 3003 27443
rect 3049 27397 3169 27443
rect 3215 27397 3256 27443
rect 2962 27261 3256 27397
rect 2962 27215 3003 27261
rect 3049 27215 3169 27261
rect 3215 27215 3256 27261
rect 2962 27178 3256 27215
rect 3361 27805 3476 27842
rect 3361 27759 3395 27805
rect 3441 27759 3476 27805
rect 3361 27624 3476 27759
rect 3361 27611 3395 27624
rect 3441 27611 3476 27624
rect 3361 27455 3391 27611
rect 3443 27455 3476 27611
rect 3361 27443 3476 27455
rect 3361 27397 3395 27443
rect 3441 27397 3476 27443
rect 3361 27261 3476 27397
rect 3361 27215 3395 27261
rect 3441 27215 3476 27261
rect 3361 27178 3476 27215
rect 3581 27805 3875 27990
rect 3980 28581 4095 28617
rect 3980 28535 4015 28581
rect 4061 28535 4095 28581
rect 3980 28399 4095 28535
rect 3980 28386 4015 28399
rect 4061 28386 4095 28399
rect 3980 28230 4013 28386
rect 4065 28230 4095 28386
rect 3980 28218 4095 28230
rect 3980 28172 4015 28218
rect 4061 28172 4095 28218
rect 3980 28036 4095 28172
rect 3980 27990 4015 28036
rect 4061 27990 4095 28036
rect 3980 27953 4095 27990
rect 4200 28581 4495 28697
rect 4200 28535 4241 28581
rect 4287 28535 4408 28581
rect 4454 28535 4495 28581
rect 4200 28399 4495 28535
rect 4200 28353 4241 28399
rect 4287 28353 4408 28399
rect 4454 28353 4495 28399
rect 4200 28218 4495 28353
rect 4200 28172 4241 28218
rect 4287 28172 4408 28218
rect 4454 28172 4495 28218
rect 4200 28036 4495 28172
rect 4200 27990 4241 28036
rect 4287 27990 4408 28036
rect 4454 27990 4495 28036
rect 3581 27759 3705 27805
rect 3751 27759 3875 27805
rect 3581 27624 3875 27759
rect 3581 27578 3705 27624
rect 3751 27578 3875 27624
rect 3581 27443 3875 27578
rect 3581 27397 3705 27443
rect 3751 27397 3875 27443
rect 3581 27261 3875 27397
rect 3581 27215 3705 27261
rect 3751 27215 3875 27261
rect 3581 27178 3875 27215
rect 3980 27805 4095 27842
rect 3980 27759 4015 27805
rect 4061 27759 4095 27805
rect 3980 27624 4095 27759
rect 3980 27611 4015 27624
rect 4061 27611 4095 27624
rect 3980 27455 4013 27611
rect 4065 27455 4095 27611
rect 3980 27443 4095 27455
rect 3980 27397 4015 27443
rect 4061 27397 4095 27443
rect 3980 27261 4095 27397
rect 3980 27215 4015 27261
rect 4061 27215 4095 27261
rect 3980 27178 4095 27215
rect 4200 27805 4495 27990
rect 4600 28581 4715 28617
rect 4600 28535 4634 28581
rect 4680 28535 4715 28581
rect 4600 28399 4715 28535
rect 4600 28386 4634 28399
rect 4680 28386 4715 28399
rect 4600 28230 4630 28386
rect 4682 28230 4715 28386
rect 4600 28218 4715 28230
rect 4600 28172 4634 28218
rect 4680 28172 4715 28218
rect 4600 28036 4715 28172
rect 4600 27990 4634 28036
rect 4680 27990 4715 28036
rect 4600 27953 4715 27990
rect 4820 28581 5025 28697
rect 4820 28535 4944 28581
rect 4990 28535 5025 28581
rect 4820 28399 5025 28535
rect 4820 28353 4944 28399
rect 4990 28353 5025 28399
rect 4820 28218 5025 28353
rect 4820 28172 4944 28218
rect 4990 28172 5025 28218
rect 4820 28036 5025 28172
rect 4820 27990 4944 28036
rect 4990 27990 5025 28036
rect 4200 27759 4241 27805
rect 4287 27759 4408 27805
rect 4454 27759 4495 27805
rect 4200 27624 4495 27759
rect 4200 27578 4241 27624
rect 4287 27578 4408 27624
rect 4454 27578 4495 27624
rect 4200 27443 4495 27578
rect 4200 27397 4241 27443
rect 4287 27397 4408 27443
rect 4454 27397 4495 27443
rect 4200 27261 4495 27397
rect 4200 27215 4241 27261
rect 4287 27215 4408 27261
rect 4454 27215 4495 27261
rect 4200 27178 4495 27215
rect 4600 27805 4715 27842
rect 4600 27759 4634 27805
rect 4680 27759 4715 27805
rect 4600 27624 4715 27759
rect 4600 27611 4634 27624
rect 4680 27611 4715 27624
rect 4600 27455 4630 27611
rect 4682 27455 4715 27611
rect 4600 27443 4715 27455
rect 4600 27397 4634 27443
rect 4680 27397 4715 27443
rect 4600 27261 4715 27397
rect 4600 27215 4634 27261
rect 4680 27215 4715 27261
rect 4600 27178 4715 27215
rect 4820 27805 5025 27990
rect 5184 28581 5300 28617
rect 5184 28535 5219 28581
rect 5265 28535 5300 28581
rect 5184 28399 5300 28535
rect 5184 28353 5219 28399
rect 5265 28386 5300 28399
rect 5184 28334 5226 28353
rect 5278 28334 5300 28386
rect 5184 28218 5300 28334
rect 5184 28172 5219 28218
rect 5265 28200 5300 28218
rect 5184 28148 5226 28172
rect 5278 28148 5300 28200
rect 5184 28036 5300 28148
rect 5184 27990 5219 28036
rect 5265 27990 5300 28036
rect 5184 27953 5300 27990
rect 5445 28581 5587 28697
rect 5445 28535 5480 28581
rect 5526 28535 5587 28581
rect 5445 28399 5587 28535
rect 5445 28353 5480 28399
rect 5526 28353 5587 28399
rect 5445 28218 5587 28353
rect 5445 28172 5480 28218
rect 5526 28172 5587 28218
rect 5445 28036 5587 28172
rect 5445 27990 5480 28036
rect 5526 27990 5587 28036
rect 4820 27759 4944 27805
rect 4990 27759 5025 27805
rect 4820 27624 5025 27759
rect 4820 27578 4944 27624
rect 4990 27578 5025 27624
rect 4820 27443 5025 27578
rect 4820 27397 4944 27443
rect 4990 27397 5025 27443
rect 4820 27261 5025 27397
rect 4820 27215 4944 27261
rect 4990 27215 5025 27261
rect 4820 27178 5025 27215
rect 5184 27805 5300 27842
rect 5184 27759 5219 27805
rect 5265 27759 5300 27805
rect 5184 27624 5300 27759
rect 5184 27611 5219 27624
rect 5265 27611 5300 27624
rect 5184 27455 5216 27611
rect 5268 27455 5300 27611
rect 5184 27443 5300 27455
rect 5184 27397 5219 27443
rect 5265 27397 5300 27443
rect 5184 27261 5300 27397
rect 5184 27215 5219 27261
rect 5265 27215 5300 27261
rect 5184 27178 5300 27215
rect 5445 27805 5587 27990
rect 5445 27759 5480 27805
rect 5526 27759 5587 27805
rect 5445 27624 5587 27759
rect 5445 27578 5480 27624
rect 5526 27578 5587 27624
rect 5445 27443 5587 27578
rect 5445 27397 5480 27443
rect 5526 27397 5587 27443
rect 5445 27261 5587 27397
rect 5445 27215 5480 27261
rect 5526 27215 5587 27261
rect 5445 27178 5587 27215
rect 412 27098 540 27118
rect 412 27097 5519 27098
rect 412 27045 448 27097
rect 500 27086 5519 27097
rect 500 27045 847 27086
rect 412 27040 847 27045
rect 1081 27040 1421 27086
rect 1655 27040 2086 27086
rect 2320 27040 2660 27086
rect 2894 27040 3324 27086
rect 3558 27040 3898 27086
rect 4132 27040 4563 27086
rect 4797 27082 5519 27086
rect 4797 27040 5122 27082
rect 412 27036 5122 27040
rect 5356 27036 5519 27082
rect 412 27025 5519 27036
rect 530 27024 5519 27025
rect 808 26937 854 26950
rect 808 26829 854 26891
rect 808 26721 854 26783
rect 808 26613 854 26675
rect 808 26505 854 26567
rect 808 26403 854 26459
rect 687 26397 854 26403
rect 687 26391 808 26397
rect 687 26235 699 26391
rect 751 26351 808 26391
rect 751 26289 854 26351
rect 751 26243 808 26289
rect 751 26235 854 26243
rect 687 26223 854 26235
rect 808 26182 854 26223
rect 808 26075 854 26136
rect 808 25968 854 26029
rect 808 25861 854 25922
rect 808 25754 854 25815
rect 808 25647 854 25708
rect 808 25588 854 25601
rect 1032 26937 1078 26950
rect 1032 26829 1078 26891
rect 1032 26721 1078 26783
rect 1032 26613 1078 26675
rect 1032 26505 1078 26567
rect 1032 26403 1078 26459
rect 1424 26937 1470 26950
rect 1424 26829 1470 26891
rect 1424 26721 1470 26783
rect 1424 26613 1470 26675
rect 1424 26505 1470 26567
rect 1424 26403 1470 26459
rect 1032 26397 1193 26403
rect 1078 26391 1193 26397
rect 1078 26351 1129 26391
rect 1032 26289 1129 26351
rect 1078 26243 1129 26289
rect 1032 26235 1129 26243
rect 1181 26235 1193 26391
rect 1032 26223 1193 26235
rect 1309 26397 1470 26403
rect 1309 26391 1424 26397
rect 1309 26235 1321 26391
rect 1373 26351 1424 26391
rect 1373 26289 1470 26351
rect 1373 26243 1424 26289
rect 1373 26235 1470 26243
rect 1309 26223 1470 26235
rect 1032 26182 1078 26223
rect 1032 26075 1078 26136
rect 1032 25968 1078 26029
rect 1032 25861 1078 25922
rect 1032 25754 1078 25815
rect 1032 25647 1078 25708
rect 1032 25588 1078 25601
rect 1424 26182 1470 26223
rect 1424 26075 1470 26136
rect 1424 25968 1470 26029
rect 1424 25861 1470 25922
rect 1424 25754 1470 25815
rect 1424 25647 1470 25708
rect 1424 25588 1470 25601
rect 1648 26937 1694 26950
rect 1648 26829 1694 26891
rect 1648 26721 1694 26783
rect 1648 26613 1694 26675
rect 1648 26505 1694 26567
rect 1648 26403 1694 26459
rect 2047 26937 2093 26950
rect 2047 26829 2093 26891
rect 2047 26721 2093 26783
rect 2047 26613 2093 26675
rect 2047 26505 2093 26567
rect 2047 26403 2093 26459
rect 1648 26397 1815 26403
rect 1694 26391 1815 26397
rect 1694 26351 1751 26391
rect 1648 26289 1751 26351
rect 1694 26243 1751 26289
rect 1648 26235 1751 26243
rect 1803 26235 1815 26391
rect 1648 26223 1815 26235
rect 1926 26397 2093 26403
rect 1926 26391 2047 26397
rect 1926 26235 1938 26391
rect 1990 26351 2047 26391
rect 1990 26289 2093 26351
rect 1990 26243 2047 26289
rect 1990 26235 2093 26243
rect 1926 26223 2093 26235
rect 1648 26182 1694 26223
rect 1648 26075 1694 26136
rect 1648 25968 1694 26029
rect 1648 25861 1694 25922
rect 1648 25754 1694 25815
rect 1648 25647 1694 25708
rect 1648 25588 1694 25601
rect 2047 26182 2093 26223
rect 2047 26075 2093 26136
rect 2047 25968 2093 26029
rect 2047 25861 2093 25922
rect 2047 25754 2093 25815
rect 2047 25647 2093 25708
rect 2047 25588 2093 25601
rect 2271 26937 2317 26950
rect 2271 26829 2317 26891
rect 2271 26721 2317 26783
rect 2271 26613 2317 26675
rect 2271 26505 2317 26567
rect 2271 26403 2317 26459
rect 2663 26937 2709 26950
rect 2663 26829 2709 26891
rect 2663 26721 2709 26783
rect 2663 26613 2709 26675
rect 2663 26505 2709 26567
rect 2663 26403 2709 26459
rect 2271 26397 2432 26403
rect 2317 26391 2432 26397
rect 2317 26351 2368 26391
rect 2271 26289 2368 26351
rect 2317 26243 2368 26289
rect 2271 26235 2368 26243
rect 2420 26235 2432 26391
rect 2271 26223 2432 26235
rect 2548 26397 2709 26403
rect 2548 26391 2663 26397
rect 2548 26235 2560 26391
rect 2612 26351 2663 26391
rect 2612 26289 2709 26351
rect 2612 26243 2663 26289
rect 2612 26235 2709 26243
rect 2548 26223 2709 26235
rect 2271 26182 2317 26223
rect 2271 26075 2317 26136
rect 2271 25968 2317 26029
rect 2271 25861 2317 25922
rect 2271 25754 2317 25815
rect 2271 25647 2317 25708
rect 2271 25588 2317 25601
rect 2663 26182 2709 26223
rect 2663 26075 2709 26136
rect 2663 25968 2709 26029
rect 2663 25861 2709 25922
rect 2663 25754 2709 25815
rect 2663 25647 2709 25708
rect 2663 25588 2709 25601
rect 2887 26937 2933 26950
rect 2887 26829 2933 26891
rect 2887 26721 2933 26783
rect 2887 26613 2933 26675
rect 2887 26505 2933 26567
rect 2887 26403 2933 26459
rect 3285 26937 3331 26950
rect 3285 26829 3331 26891
rect 3285 26721 3331 26783
rect 3285 26613 3331 26675
rect 3285 26505 3331 26567
rect 3285 26403 3331 26459
rect 2887 26397 3054 26403
rect 2933 26391 3054 26397
rect 2933 26351 2990 26391
rect 2887 26289 2990 26351
rect 2933 26243 2990 26289
rect 2887 26235 2990 26243
rect 3042 26235 3054 26391
rect 2887 26223 3054 26235
rect 3164 26397 3331 26403
rect 3164 26391 3285 26397
rect 3164 26235 3176 26391
rect 3228 26351 3285 26391
rect 3228 26289 3331 26351
rect 3228 26243 3285 26289
rect 3228 26235 3331 26243
rect 3164 26223 3331 26235
rect 2887 26182 2933 26223
rect 2887 26075 2933 26136
rect 2887 25968 2933 26029
rect 2887 25861 2933 25922
rect 2887 25754 2933 25815
rect 2887 25647 2933 25708
rect 2887 25588 2933 25601
rect 3285 26182 3331 26223
rect 3285 26075 3331 26136
rect 3285 25968 3331 26029
rect 3285 25861 3331 25922
rect 3285 25754 3331 25815
rect 3285 25647 3331 25708
rect 3285 25588 3331 25601
rect 3509 26937 3555 26950
rect 3509 26829 3555 26891
rect 3509 26721 3555 26783
rect 3509 26613 3555 26675
rect 3509 26505 3555 26567
rect 3509 26403 3555 26459
rect 3901 26937 3947 26950
rect 3901 26829 3947 26891
rect 3901 26721 3947 26783
rect 3901 26613 3947 26675
rect 3901 26505 3947 26567
rect 3901 26403 3947 26459
rect 3509 26397 3670 26403
rect 3555 26391 3670 26397
rect 3555 26351 3606 26391
rect 3509 26289 3606 26351
rect 3555 26243 3606 26289
rect 3509 26235 3606 26243
rect 3658 26235 3670 26391
rect 3509 26223 3670 26235
rect 3786 26397 3947 26403
rect 3786 26391 3901 26397
rect 3786 26235 3798 26391
rect 3850 26351 3901 26391
rect 3850 26289 3947 26351
rect 3850 26243 3901 26289
rect 3850 26235 3947 26243
rect 3786 26223 3947 26235
rect 3509 26182 3555 26223
rect 3509 26075 3555 26136
rect 3509 25968 3555 26029
rect 3509 25861 3555 25922
rect 3509 25754 3555 25815
rect 3509 25647 3555 25708
rect 3509 25588 3555 25601
rect 3901 26182 3947 26223
rect 3901 26075 3947 26136
rect 3901 25968 3947 26029
rect 3901 25861 3947 25922
rect 3901 25754 3947 25815
rect 3901 25647 3947 25708
rect 3901 25588 3947 25601
rect 4125 26937 4171 26950
rect 4125 26829 4171 26891
rect 4125 26721 4171 26783
rect 4125 26613 4171 26675
rect 4125 26505 4171 26567
rect 4125 26403 4171 26459
rect 4524 26937 4570 26950
rect 4524 26829 4570 26891
rect 4524 26721 4570 26783
rect 4524 26613 4570 26675
rect 4524 26505 4570 26567
rect 4524 26403 4570 26459
rect 4125 26397 4292 26403
rect 4171 26391 4292 26397
rect 4171 26351 4228 26391
rect 4125 26289 4228 26351
rect 4171 26243 4228 26289
rect 4125 26235 4228 26243
rect 4280 26235 4292 26391
rect 4125 26223 4292 26235
rect 4403 26397 4570 26403
rect 4403 26391 4524 26397
rect 4403 26235 4415 26391
rect 4467 26351 4524 26391
rect 4467 26289 4570 26351
rect 4467 26243 4524 26289
rect 4467 26235 4570 26243
rect 4403 26223 4570 26235
rect 4125 26182 4171 26223
rect 4125 26075 4171 26136
rect 4125 25968 4171 26029
rect 4125 25861 4171 25922
rect 4125 25754 4171 25815
rect 4125 25647 4171 25708
rect 4125 25588 4171 25601
rect 4524 26182 4570 26223
rect 4524 26075 4570 26136
rect 4524 25968 4570 26029
rect 4524 25861 4570 25922
rect 4524 25754 4570 25815
rect 4524 25647 4570 25708
rect 4524 25588 4570 25601
rect 4748 26937 4794 26950
rect 4748 26829 4794 26891
rect 4748 26721 4794 26783
rect 4748 26613 4794 26675
rect 4748 26505 4794 26567
rect 4748 26403 4794 26459
rect 5140 26937 5186 26950
rect 5140 26829 5186 26891
rect 5140 26721 5186 26783
rect 5140 26613 5186 26675
rect 5140 26505 5186 26567
rect 5140 26403 5186 26459
rect 4748 26397 4909 26403
rect 4794 26391 4909 26397
rect 4794 26351 4845 26391
rect 4748 26289 4845 26351
rect 4794 26243 4845 26289
rect 4748 26235 4845 26243
rect 4897 26235 4909 26391
rect 4748 26223 4909 26235
rect 5029 26397 5186 26403
rect 5029 26391 5140 26397
rect 5029 26235 5041 26391
rect 5093 26351 5140 26391
rect 5093 26289 5186 26351
rect 5093 26243 5140 26289
rect 5093 26235 5186 26243
rect 5029 26223 5186 26235
rect 4748 26182 4794 26223
rect 4748 26075 4794 26136
rect 4748 25968 4794 26029
rect 4748 25861 4794 25922
rect 4748 25754 4794 25815
rect 4748 25647 4794 25708
rect 4748 25588 4794 25601
rect 5140 26182 5186 26223
rect 5140 26075 5186 26136
rect 5140 25968 5186 26029
rect 5140 25861 5186 25922
rect 5140 25754 5186 25815
rect 5140 25647 5186 25708
rect 5140 25588 5186 25601
rect 5364 26937 5410 26950
rect 5364 26829 5410 26891
rect 5364 26721 5410 26783
rect 5364 26613 5410 26675
rect 5364 26505 5410 26567
rect 5364 26403 5410 26459
rect 5364 26397 5523 26403
rect 5410 26391 5523 26397
rect 5410 26351 5459 26391
rect 5364 26289 5459 26351
rect 5410 26243 5459 26289
rect 5364 26235 5459 26243
rect 5511 26235 5523 26391
rect 5364 26223 5523 26235
rect 5364 26182 5410 26223
rect 5364 26075 5410 26136
rect 5364 25968 5410 26029
rect 5364 25861 5410 25922
rect 5364 25754 5410 25815
rect 5364 25647 5410 25708
rect 5364 25588 5410 25601
rect 702 25350 852 25363
rect 702 25304 806 25350
rect 702 25242 852 25304
rect 702 25196 806 25242
rect 702 25134 852 25196
rect 702 25088 806 25134
rect 702 25026 852 25088
rect 702 24980 806 25026
rect 702 24918 852 24980
rect 702 24872 806 24918
rect 702 24810 852 24872
rect 702 24764 806 24810
rect 702 24702 852 24764
rect 702 24656 806 24702
rect 702 24595 852 24656
rect 702 24549 806 24595
rect 702 24488 852 24549
rect 702 24442 806 24488
rect 702 24381 852 24442
rect 702 24335 806 24381
rect 702 24274 852 24335
rect 702 24228 806 24274
rect 702 24167 852 24228
rect 702 24121 806 24167
rect 702 24060 852 24121
rect 702 24014 806 24060
rect 702 24001 852 24014
rect 1030 25351 1181 25363
rect 1030 25350 1117 25351
rect 1076 25304 1117 25350
rect 1030 25242 1117 25304
rect 1076 25196 1117 25242
rect 1030 25195 1117 25196
rect 1169 25195 1181 25351
rect 1030 25134 1181 25195
rect 1076 25088 1181 25134
rect 1030 25026 1181 25088
rect 1076 24980 1181 25026
rect 1030 24918 1181 24980
rect 1076 24872 1181 24918
rect 1030 24810 1181 24872
rect 1076 24798 1181 24810
rect 1321 25351 1472 25363
rect 1321 25195 1333 25351
rect 1385 25350 1472 25351
rect 1385 25304 1426 25350
rect 1385 25242 1472 25304
rect 1385 25196 1426 25242
rect 1385 25195 1472 25196
rect 1321 25134 1472 25195
rect 1321 25088 1426 25134
rect 1321 25026 1472 25088
rect 1321 24980 1426 25026
rect 1321 24918 1472 24980
rect 1321 24872 1426 24918
rect 1321 24810 1472 24872
rect 1321 24798 1426 24810
rect 1076 24764 1137 24798
rect 1030 24702 1137 24764
rect 1076 24656 1137 24702
rect 1365 24764 1426 24798
rect 1365 24702 1472 24764
rect 1030 24595 1137 24656
rect 1076 24549 1137 24595
rect 1030 24488 1137 24549
rect 1076 24442 1137 24488
rect 1030 24381 1137 24442
rect 1213 24677 1289 24689
rect 1213 24417 1225 24677
rect 1277 24417 1289 24677
rect 1213 24416 1228 24417
rect 1274 24416 1289 24417
rect 1213 24405 1289 24416
rect 1365 24656 1426 24702
rect 1365 24595 1472 24656
rect 1365 24549 1426 24595
rect 1365 24488 1472 24549
rect 1365 24442 1426 24488
rect 1076 24335 1137 24381
rect 1030 24278 1137 24335
rect 1365 24381 1472 24442
rect 1365 24335 1426 24381
rect 1365 24278 1472 24335
rect 1030 24274 1181 24278
rect 1076 24228 1181 24274
rect 1030 24167 1181 24228
rect 1076 24121 1181 24167
rect 1030 24060 1181 24121
rect 1076 24014 1181 24060
rect 1030 24001 1181 24014
rect 702 23672 772 24001
rect 851 23919 1032 23931
rect 851 23763 909 23919
rect 961 23763 1032 23919
rect 851 23748 1032 23763
rect 1110 23672 1181 24001
rect 702 23659 852 23672
rect 702 23613 806 23659
rect 702 23551 852 23613
rect 702 23505 806 23551
rect 702 23443 852 23505
rect 702 23397 806 23443
rect 702 23335 852 23397
rect 702 23289 806 23335
rect 702 23227 852 23289
rect 702 23181 806 23227
rect 702 23119 852 23181
rect 702 23073 806 23119
rect 702 23011 852 23073
rect 702 22965 806 23011
rect 702 22904 852 22965
rect 702 22858 806 22904
rect 702 22797 852 22858
rect 702 22751 806 22797
rect 702 22690 852 22751
rect 702 22644 806 22690
rect 702 22583 852 22644
rect 702 22537 806 22583
rect 702 22476 852 22537
rect 702 22430 806 22476
rect 702 22369 852 22430
rect 702 22323 806 22369
rect 702 22320 852 22323
rect 806 22240 852 22320
rect 1030 23659 1181 23672
rect 1076 23613 1181 23659
rect 1030 23551 1181 23613
rect 1076 23505 1181 23551
rect 1030 23443 1181 23505
rect 1076 23397 1181 23443
rect 1030 23335 1181 23397
rect 1076 23289 1181 23335
rect 1030 23227 1181 23289
rect 1076 23181 1181 23227
rect 1030 23119 1181 23181
rect 1076 23073 1181 23119
rect 1030 23011 1181 23073
rect 1076 22965 1181 23011
rect 1030 22904 1181 22965
rect 1076 22858 1181 22904
rect 1030 22797 1181 22858
rect 1076 22751 1181 22797
rect 1030 22690 1181 22751
rect 1076 22644 1181 22690
rect 1030 22583 1181 22644
rect 1076 22537 1181 22583
rect 1030 22476 1181 22537
rect 1076 22430 1181 22476
rect 1030 22369 1181 22430
rect 1076 22323 1181 22369
rect 1030 22310 1181 22323
rect 1321 24274 1472 24278
rect 1321 24228 1426 24274
rect 1321 24167 1472 24228
rect 1321 24121 1426 24167
rect 1321 24060 1472 24121
rect 1321 24014 1426 24060
rect 1321 24001 1472 24014
rect 1650 25350 1800 25363
rect 1696 25304 1800 25350
rect 1650 25242 1800 25304
rect 1696 25196 1800 25242
rect 1650 25134 1800 25196
rect 1696 25088 1800 25134
rect 1650 25026 1800 25088
rect 1696 24980 1800 25026
rect 1650 24918 1800 24980
rect 1696 24872 1800 24918
rect 1650 24810 1800 24872
rect 1696 24764 1800 24810
rect 1650 24702 1800 24764
rect 1696 24656 1800 24702
rect 1650 24595 1800 24656
rect 1696 24549 1800 24595
rect 1650 24488 1800 24549
rect 1696 24442 1800 24488
rect 1650 24381 1800 24442
rect 1696 24335 1800 24381
rect 1650 24274 1800 24335
rect 1696 24228 1800 24274
rect 1650 24167 1800 24228
rect 1696 24121 1800 24167
rect 1650 24060 1800 24121
rect 1696 24014 1800 24060
rect 1650 24001 1800 24014
rect 1321 23672 1392 24001
rect 1470 23919 1651 23931
rect 1470 23763 1541 23919
rect 1593 23763 1651 23919
rect 1470 23748 1651 23763
rect 1730 23672 1800 24001
rect 1321 23659 1472 23672
rect 1321 23613 1426 23659
rect 1321 23551 1472 23613
rect 1321 23505 1426 23551
rect 1321 23443 1472 23505
rect 1321 23397 1426 23443
rect 1321 23335 1472 23397
rect 1321 23289 1426 23335
rect 1321 23227 1472 23289
rect 1321 23181 1426 23227
rect 1321 23119 1472 23181
rect 1321 23073 1426 23119
rect 1321 23011 1472 23073
rect 1321 22965 1426 23011
rect 1321 22904 1472 22965
rect 1321 22858 1426 22904
rect 1321 22797 1472 22858
rect 1321 22751 1426 22797
rect 1321 22690 1472 22751
rect 1321 22644 1426 22690
rect 1321 22583 1472 22644
rect 1321 22537 1426 22583
rect 1321 22476 1472 22537
rect 1321 22430 1426 22476
rect 1321 22369 1472 22430
rect 1321 22323 1426 22369
rect 1321 22310 1472 22323
rect 1650 23659 1800 23672
rect 1696 23613 1800 23659
rect 1650 23551 1800 23613
rect 1696 23505 1800 23551
rect 1650 23443 1800 23505
rect 1696 23397 1800 23443
rect 1650 23335 1800 23397
rect 1696 23289 1800 23335
rect 1650 23227 1800 23289
rect 1696 23181 1800 23227
rect 1650 23119 1800 23181
rect 1696 23073 1800 23119
rect 1650 23011 1800 23073
rect 1696 22965 1800 23011
rect 1650 22904 1800 22965
rect 1696 22858 1800 22904
rect 1650 22797 1800 22858
rect 1696 22751 1800 22797
rect 1650 22690 1800 22751
rect 1696 22644 1800 22690
rect 1650 22583 1800 22644
rect 1696 22537 1800 22583
rect 1650 22476 1800 22537
rect 1696 22430 1800 22476
rect 1650 22369 1800 22430
rect 1696 22323 1800 22369
rect 1650 22320 1800 22323
rect 1941 25350 2091 25363
rect 1941 25304 2045 25350
rect 1941 25242 2091 25304
rect 1941 25196 2045 25242
rect 1941 25134 2091 25196
rect 1941 25088 2045 25134
rect 1941 25026 2091 25088
rect 1941 24980 2045 25026
rect 1941 24918 2091 24980
rect 1941 24872 2045 24918
rect 1941 24810 2091 24872
rect 1941 24764 2045 24810
rect 1941 24702 2091 24764
rect 1941 24656 2045 24702
rect 1941 24595 2091 24656
rect 1941 24549 2045 24595
rect 1941 24488 2091 24549
rect 1941 24442 2045 24488
rect 1941 24381 2091 24442
rect 1941 24335 2045 24381
rect 1941 24274 2091 24335
rect 1941 24228 2045 24274
rect 1941 24167 2091 24228
rect 1941 24121 2045 24167
rect 1941 24060 2091 24121
rect 1941 24014 2045 24060
rect 1941 24001 2091 24014
rect 2269 25351 2420 25363
rect 2269 25350 2356 25351
rect 2315 25304 2356 25350
rect 2269 25242 2356 25304
rect 2315 25196 2356 25242
rect 2269 25195 2356 25196
rect 2408 25195 2420 25351
rect 2269 25134 2420 25195
rect 2315 25088 2420 25134
rect 2269 25026 2420 25088
rect 2315 24980 2420 25026
rect 2269 24918 2420 24980
rect 2315 24872 2420 24918
rect 2269 24810 2420 24872
rect 2315 24798 2420 24810
rect 2560 25351 2711 25363
rect 2560 25195 2572 25351
rect 2624 25350 2711 25351
rect 2624 25304 2665 25350
rect 2624 25242 2711 25304
rect 2624 25196 2665 25242
rect 2624 25195 2711 25196
rect 2560 25134 2711 25195
rect 2560 25088 2665 25134
rect 2560 25026 2711 25088
rect 2560 24980 2665 25026
rect 2560 24918 2711 24980
rect 2560 24872 2665 24918
rect 2560 24810 2711 24872
rect 2560 24798 2665 24810
rect 2315 24764 2376 24798
rect 2269 24702 2376 24764
rect 2315 24656 2376 24702
rect 2604 24764 2665 24798
rect 2604 24702 2711 24764
rect 2269 24595 2376 24656
rect 2315 24549 2376 24595
rect 2269 24488 2376 24549
rect 2315 24442 2376 24488
rect 2269 24381 2376 24442
rect 2452 24677 2528 24689
rect 2452 24417 2464 24677
rect 2516 24417 2528 24677
rect 2452 24416 2467 24417
rect 2513 24416 2528 24417
rect 2452 24405 2528 24416
rect 2604 24656 2665 24702
rect 2604 24595 2711 24656
rect 2604 24549 2665 24595
rect 2604 24488 2711 24549
rect 2604 24442 2665 24488
rect 2315 24335 2376 24381
rect 2269 24278 2376 24335
rect 2604 24381 2711 24442
rect 2604 24335 2665 24381
rect 2604 24278 2711 24335
rect 2269 24274 2420 24278
rect 2315 24228 2420 24274
rect 2269 24167 2420 24228
rect 2315 24121 2420 24167
rect 2269 24060 2420 24121
rect 2315 24014 2420 24060
rect 2269 24001 2420 24014
rect 1941 23672 2011 24001
rect 2090 23919 2271 23931
rect 2090 23763 2148 23919
rect 2200 23763 2271 23919
rect 2090 23748 2271 23763
rect 2349 23672 2420 24001
rect 1941 23659 2091 23672
rect 1941 23613 2045 23659
rect 1941 23551 2091 23613
rect 1941 23505 2045 23551
rect 1941 23443 2091 23505
rect 1941 23397 2045 23443
rect 1941 23335 2091 23397
rect 1941 23289 2045 23335
rect 1941 23227 2091 23289
rect 1941 23181 2045 23227
rect 1941 23119 2091 23181
rect 1941 23073 2045 23119
rect 1941 23011 2091 23073
rect 1941 22965 2045 23011
rect 1941 22904 2091 22965
rect 1941 22858 2045 22904
rect 1941 22797 2091 22858
rect 1941 22751 2045 22797
rect 1941 22690 2091 22751
rect 1941 22644 2045 22690
rect 1941 22583 2091 22644
rect 1941 22537 2045 22583
rect 1941 22476 2091 22537
rect 1941 22430 2045 22476
rect 1941 22369 2091 22430
rect 1941 22323 2045 22369
rect 1941 22320 2091 22323
rect 1650 22240 1696 22320
rect 806 22218 1206 22240
rect 806 22166 1124 22218
rect 1176 22166 1206 22218
rect 806 22143 1206 22166
rect 1296 22218 1696 22240
rect 1296 22166 1326 22218
rect 1378 22166 1696 22218
rect 1296 22143 1696 22166
rect 2045 22240 2091 22320
rect 2269 23659 2420 23672
rect 2315 23613 2420 23659
rect 2269 23551 2420 23613
rect 2315 23505 2420 23551
rect 2269 23443 2420 23505
rect 2315 23397 2420 23443
rect 2269 23335 2420 23397
rect 2315 23289 2420 23335
rect 2269 23227 2420 23289
rect 2315 23181 2420 23227
rect 2269 23119 2420 23181
rect 2315 23073 2420 23119
rect 2269 23011 2420 23073
rect 2315 22965 2420 23011
rect 2269 22904 2420 22965
rect 2315 22858 2420 22904
rect 2269 22797 2420 22858
rect 2315 22751 2420 22797
rect 2269 22690 2420 22751
rect 2315 22644 2420 22690
rect 2269 22583 2420 22644
rect 2315 22537 2420 22583
rect 2269 22476 2420 22537
rect 2315 22430 2420 22476
rect 2269 22369 2420 22430
rect 2315 22323 2420 22369
rect 2269 22310 2420 22323
rect 2560 24274 2711 24278
rect 2560 24228 2665 24274
rect 2560 24167 2711 24228
rect 2560 24121 2665 24167
rect 2560 24060 2711 24121
rect 2560 24014 2665 24060
rect 2560 24001 2711 24014
rect 2889 25350 3039 25363
rect 2935 25304 3039 25350
rect 2889 25242 3039 25304
rect 2935 25196 3039 25242
rect 2889 25134 3039 25196
rect 2935 25088 3039 25134
rect 2889 25026 3039 25088
rect 2935 24980 3039 25026
rect 2889 24918 3039 24980
rect 2935 24872 3039 24918
rect 2889 24810 3039 24872
rect 2935 24764 3039 24810
rect 2889 24702 3039 24764
rect 2935 24656 3039 24702
rect 2889 24595 3039 24656
rect 2935 24549 3039 24595
rect 2889 24488 3039 24549
rect 2935 24442 3039 24488
rect 2889 24381 3039 24442
rect 2935 24335 3039 24381
rect 2889 24274 3039 24335
rect 2935 24228 3039 24274
rect 2889 24167 3039 24228
rect 2935 24121 3039 24167
rect 2889 24060 3039 24121
rect 2935 24014 3039 24060
rect 2889 24001 3039 24014
rect 2560 23672 2631 24001
rect 2709 23919 2890 23931
rect 2709 23763 2780 23919
rect 2832 23763 2890 23919
rect 2709 23748 2890 23763
rect 2969 23672 3039 24001
rect 2560 23659 2711 23672
rect 2560 23613 2665 23659
rect 2560 23551 2711 23613
rect 2560 23505 2665 23551
rect 2560 23443 2711 23505
rect 2560 23397 2665 23443
rect 2560 23335 2711 23397
rect 2560 23289 2665 23335
rect 2560 23227 2711 23289
rect 2560 23181 2665 23227
rect 2560 23119 2711 23181
rect 2560 23073 2665 23119
rect 2560 23011 2711 23073
rect 2560 22965 2665 23011
rect 2560 22904 2711 22965
rect 2560 22858 2665 22904
rect 2560 22797 2711 22858
rect 2560 22751 2665 22797
rect 2560 22690 2711 22751
rect 2560 22644 2665 22690
rect 2560 22583 2711 22644
rect 2560 22537 2665 22583
rect 2560 22476 2711 22537
rect 2560 22430 2665 22476
rect 2560 22369 2711 22430
rect 2560 22323 2665 22369
rect 2560 22310 2711 22323
rect 2889 23659 3039 23672
rect 2935 23613 3039 23659
rect 2889 23551 3039 23613
rect 2935 23505 3039 23551
rect 2889 23443 3039 23505
rect 2935 23397 3039 23443
rect 2889 23335 3039 23397
rect 2935 23289 3039 23335
rect 2889 23227 3039 23289
rect 2935 23181 3039 23227
rect 2889 23119 3039 23181
rect 2935 23073 3039 23119
rect 2889 23011 3039 23073
rect 2935 22965 3039 23011
rect 2889 22904 3039 22965
rect 2935 22858 3039 22904
rect 2889 22797 3039 22858
rect 2935 22751 3039 22797
rect 2889 22690 3039 22751
rect 2935 22644 3039 22690
rect 2889 22583 3039 22644
rect 2935 22537 3039 22583
rect 2889 22476 3039 22537
rect 2935 22430 3039 22476
rect 2889 22369 3039 22430
rect 2935 22323 3039 22369
rect 2889 22320 3039 22323
rect 3179 25350 3329 25363
rect 3179 25304 3283 25350
rect 3179 25242 3329 25304
rect 3179 25196 3283 25242
rect 3179 25134 3329 25196
rect 3179 25088 3283 25134
rect 3179 25026 3329 25088
rect 3179 24980 3283 25026
rect 3179 24918 3329 24980
rect 3179 24872 3283 24918
rect 3179 24810 3329 24872
rect 3179 24764 3283 24810
rect 3179 24702 3329 24764
rect 3179 24656 3283 24702
rect 3179 24595 3329 24656
rect 3179 24549 3283 24595
rect 3179 24488 3329 24549
rect 3179 24442 3283 24488
rect 3179 24381 3329 24442
rect 3179 24335 3283 24381
rect 3179 24274 3329 24335
rect 3179 24228 3283 24274
rect 3179 24167 3329 24228
rect 3179 24121 3283 24167
rect 3179 24060 3329 24121
rect 3179 24014 3283 24060
rect 3179 24001 3329 24014
rect 3507 25351 3658 25363
rect 3507 25350 3594 25351
rect 3553 25304 3594 25350
rect 3507 25242 3594 25304
rect 3553 25196 3594 25242
rect 3507 25195 3594 25196
rect 3646 25195 3658 25351
rect 3507 25134 3658 25195
rect 3553 25088 3658 25134
rect 3507 25026 3658 25088
rect 3553 24980 3658 25026
rect 3507 24918 3658 24980
rect 3553 24872 3658 24918
rect 3507 24810 3658 24872
rect 3553 24798 3658 24810
rect 3798 25351 3949 25363
rect 3798 25195 3810 25351
rect 3862 25350 3949 25351
rect 3862 25304 3903 25350
rect 3862 25242 3949 25304
rect 3862 25196 3903 25242
rect 3862 25195 3949 25196
rect 3798 25134 3949 25195
rect 3798 25088 3903 25134
rect 3798 25026 3949 25088
rect 3798 24980 3903 25026
rect 3798 24918 3949 24980
rect 3798 24872 3903 24918
rect 3798 24810 3949 24872
rect 3798 24798 3903 24810
rect 3553 24764 3614 24798
rect 3507 24702 3614 24764
rect 3553 24656 3614 24702
rect 3842 24764 3903 24798
rect 3842 24702 3949 24764
rect 3507 24595 3614 24656
rect 3553 24549 3614 24595
rect 3507 24488 3614 24549
rect 3553 24442 3614 24488
rect 3507 24381 3614 24442
rect 3690 24677 3766 24689
rect 3690 24417 3702 24677
rect 3754 24417 3766 24677
rect 3690 24416 3705 24417
rect 3751 24416 3766 24417
rect 3690 24405 3766 24416
rect 3842 24656 3903 24702
rect 3842 24595 3949 24656
rect 3842 24549 3903 24595
rect 3842 24488 3949 24549
rect 3842 24442 3903 24488
rect 3553 24335 3614 24381
rect 3507 24278 3614 24335
rect 3842 24381 3949 24442
rect 3842 24335 3903 24381
rect 3842 24278 3949 24335
rect 3507 24274 3658 24278
rect 3553 24228 3658 24274
rect 3507 24167 3658 24228
rect 3553 24121 3658 24167
rect 3507 24060 3658 24121
rect 3553 24014 3658 24060
rect 3507 24001 3658 24014
rect 3179 23672 3249 24001
rect 3328 23919 3509 23931
rect 3328 23763 3386 23919
rect 3438 23763 3509 23919
rect 3328 23748 3509 23763
rect 3587 23672 3658 24001
rect 3179 23659 3329 23672
rect 3179 23613 3283 23659
rect 3179 23551 3329 23613
rect 3179 23505 3283 23551
rect 3179 23443 3329 23505
rect 3179 23397 3283 23443
rect 3179 23335 3329 23397
rect 3179 23289 3283 23335
rect 3179 23227 3329 23289
rect 3179 23181 3283 23227
rect 3179 23119 3329 23181
rect 3179 23073 3283 23119
rect 3179 23011 3329 23073
rect 3179 22965 3283 23011
rect 3179 22904 3329 22965
rect 3179 22858 3283 22904
rect 3179 22797 3329 22858
rect 3179 22751 3283 22797
rect 3179 22690 3329 22751
rect 3179 22644 3283 22690
rect 3179 22583 3329 22644
rect 3179 22537 3283 22583
rect 3179 22476 3329 22537
rect 3179 22430 3283 22476
rect 3179 22369 3329 22430
rect 3179 22323 3283 22369
rect 3179 22320 3329 22323
rect 2889 22240 2935 22320
rect 2045 22218 2445 22240
rect 2045 22166 2363 22218
rect 2415 22166 2445 22218
rect 2045 22143 2445 22166
rect 2535 22218 2935 22240
rect 2535 22166 2565 22218
rect 2617 22166 2935 22218
rect 2535 22143 2935 22166
rect 3283 22240 3329 22320
rect 3507 23659 3658 23672
rect 3553 23613 3658 23659
rect 3507 23551 3658 23613
rect 3553 23505 3658 23551
rect 3507 23443 3658 23505
rect 3553 23397 3658 23443
rect 3507 23335 3658 23397
rect 3553 23289 3658 23335
rect 3507 23227 3658 23289
rect 3553 23181 3658 23227
rect 3507 23119 3658 23181
rect 3553 23073 3658 23119
rect 3507 23011 3658 23073
rect 3553 22965 3658 23011
rect 3507 22904 3658 22965
rect 3553 22858 3658 22904
rect 3507 22797 3658 22858
rect 3553 22751 3658 22797
rect 3507 22690 3658 22751
rect 3553 22644 3658 22690
rect 3507 22583 3658 22644
rect 3553 22537 3658 22583
rect 3507 22476 3658 22537
rect 3553 22430 3658 22476
rect 3507 22369 3658 22430
rect 3553 22323 3658 22369
rect 3507 22310 3658 22323
rect 3798 24274 3949 24278
rect 3798 24228 3903 24274
rect 3798 24167 3949 24228
rect 3798 24121 3903 24167
rect 3798 24060 3949 24121
rect 3798 24014 3903 24060
rect 3798 24001 3949 24014
rect 4127 25350 4277 25363
rect 4173 25304 4277 25350
rect 4127 25242 4277 25304
rect 4173 25196 4277 25242
rect 4127 25134 4277 25196
rect 4173 25088 4277 25134
rect 4127 25026 4277 25088
rect 4173 24980 4277 25026
rect 4127 24918 4277 24980
rect 4173 24872 4277 24918
rect 4127 24810 4277 24872
rect 4173 24764 4277 24810
rect 4127 24702 4277 24764
rect 4173 24656 4277 24702
rect 4127 24595 4277 24656
rect 4173 24549 4277 24595
rect 4127 24488 4277 24549
rect 4173 24442 4277 24488
rect 4127 24381 4277 24442
rect 4173 24335 4277 24381
rect 4127 24274 4277 24335
rect 4173 24228 4277 24274
rect 4127 24167 4277 24228
rect 4173 24121 4277 24167
rect 4127 24060 4277 24121
rect 4173 24014 4277 24060
rect 4127 24001 4277 24014
rect 3798 23672 3869 24001
rect 3947 23919 4128 23931
rect 3947 23763 4018 23919
rect 4070 23763 4128 23919
rect 3947 23748 4128 23763
rect 4207 23672 4277 24001
rect 3798 23659 3949 23672
rect 3798 23613 3903 23659
rect 3798 23551 3949 23613
rect 3798 23505 3903 23551
rect 3798 23443 3949 23505
rect 3798 23397 3903 23443
rect 3798 23335 3949 23397
rect 3798 23289 3903 23335
rect 3798 23227 3949 23289
rect 3798 23181 3903 23227
rect 3798 23119 3949 23181
rect 3798 23073 3903 23119
rect 3798 23011 3949 23073
rect 3798 22965 3903 23011
rect 3798 22904 3949 22965
rect 3798 22858 3903 22904
rect 3798 22797 3949 22858
rect 3798 22751 3903 22797
rect 3798 22690 3949 22751
rect 3798 22644 3903 22690
rect 3798 22583 3949 22644
rect 3798 22537 3903 22583
rect 3798 22476 3949 22537
rect 3798 22430 3903 22476
rect 3798 22369 3949 22430
rect 3798 22323 3903 22369
rect 3798 22310 3949 22323
rect 4127 23659 4277 23672
rect 4173 23613 4277 23659
rect 4127 23551 4277 23613
rect 4173 23505 4277 23551
rect 4127 23443 4277 23505
rect 4173 23397 4277 23443
rect 4127 23335 4277 23397
rect 4173 23289 4277 23335
rect 4127 23227 4277 23289
rect 4173 23181 4277 23227
rect 4127 23119 4277 23181
rect 4173 23073 4277 23119
rect 4127 23011 4277 23073
rect 4173 22965 4277 23011
rect 4127 22904 4277 22965
rect 4173 22858 4277 22904
rect 4127 22797 4277 22858
rect 4173 22751 4277 22797
rect 4127 22690 4277 22751
rect 4173 22644 4277 22690
rect 4127 22583 4277 22644
rect 4173 22537 4277 22583
rect 4127 22476 4277 22537
rect 4173 22430 4277 22476
rect 4127 22369 4277 22430
rect 4173 22323 4277 22369
rect 4127 22320 4277 22323
rect 4418 25350 4568 25363
rect 4418 25304 4522 25350
rect 4418 25242 4568 25304
rect 4418 25196 4522 25242
rect 4418 25134 4568 25196
rect 4418 25088 4522 25134
rect 4418 25026 4568 25088
rect 4418 24980 4522 25026
rect 4418 24918 4568 24980
rect 4418 24872 4522 24918
rect 4418 24810 4568 24872
rect 4418 24764 4522 24810
rect 4418 24702 4568 24764
rect 4418 24656 4522 24702
rect 4418 24595 4568 24656
rect 4418 24549 4522 24595
rect 4418 24488 4568 24549
rect 4418 24442 4522 24488
rect 4418 24381 4568 24442
rect 4418 24335 4522 24381
rect 4418 24274 4568 24335
rect 4418 24228 4522 24274
rect 4418 24167 4568 24228
rect 4418 24121 4522 24167
rect 4418 24060 4568 24121
rect 4418 24014 4522 24060
rect 4418 24001 4568 24014
rect 4746 25351 4897 25363
rect 4746 25350 4833 25351
rect 4792 25304 4833 25350
rect 4746 25242 4833 25304
rect 4792 25196 4833 25242
rect 4746 25195 4833 25196
rect 4885 25195 4897 25351
rect 4746 25134 4897 25195
rect 4792 25088 4897 25134
rect 4746 25026 4897 25088
rect 4792 24980 4897 25026
rect 4746 24918 4897 24980
rect 4792 24872 4897 24918
rect 4746 24810 4897 24872
rect 4792 24798 4897 24810
rect 5041 25351 5188 25363
rect 5041 25195 5053 25351
rect 5105 25350 5188 25351
rect 5105 25304 5142 25350
rect 5105 25242 5188 25304
rect 5105 25196 5142 25242
rect 5105 25195 5188 25196
rect 5041 25134 5188 25195
rect 5041 25088 5142 25134
rect 5041 25026 5188 25088
rect 5041 24980 5142 25026
rect 5041 24918 5188 24980
rect 5041 24872 5142 24918
rect 5041 24810 5188 24872
rect 5041 24798 5142 24810
rect 4792 24764 4853 24798
rect 4746 24702 4853 24764
rect 4792 24656 4853 24702
rect 5081 24764 5142 24798
rect 5081 24702 5188 24764
rect 4746 24595 4853 24656
rect 4792 24549 4853 24595
rect 4746 24488 4853 24549
rect 4792 24442 4853 24488
rect 4746 24381 4853 24442
rect 4929 24677 5005 24689
rect 4929 24417 4941 24677
rect 4993 24417 5005 24677
rect 4929 24416 4944 24417
rect 4990 24416 5005 24417
rect 4929 24405 5005 24416
rect 5081 24656 5142 24702
rect 5081 24595 5188 24656
rect 5081 24549 5142 24595
rect 5081 24488 5188 24549
rect 5081 24442 5142 24488
rect 4792 24335 4853 24381
rect 4746 24278 4853 24335
rect 5081 24381 5188 24442
rect 5081 24335 5142 24381
rect 5081 24278 5188 24335
rect 4746 24274 4897 24278
rect 4792 24228 4897 24274
rect 4746 24167 4897 24228
rect 4792 24121 4897 24167
rect 4746 24060 4897 24121
rect 4792 24014 4897 24060
rect 4746 24001 4897 24014
rect 4418 23672 4488 24001
rect 4567 23919 4748 23931
rect 4567 23763 4625 23919
rect 4677 23763 4748 23919
rect 4567 23748 4748 23763
rect 4826 23672 4897 24001
rect 4418 23659 4568 23672
rect 4418 23613 4522 23659
rect 4418 23551 4568 23613
rect 4418 23505 4522 23551
rect 4418 23443 4568 23505
rect 4418 23397 4522 23443
rect 4418 23335 4568 23397
rect 4418 23289 4522 23335
rect 4418 23227 4568 23289
rect 4418 23181 4522 23227
rect 4418 23119 4568 23181
rect 4418 23073 4522 23119
rect 4418 23011 4568 23073
rect 4418 22965 4522 23011
rect 4418 22904 4568 22965
rect 4418 22858 4522 22904
rect 4418 22797 4568 22858
rect 4418 22751 4522 22797
rect 4418 22690 4568 22751
rect 4418 22644 4522 22690
rect 4418 22583 4568 22644
rect 4418 22537 4522 22583
rect 4418 22476 4568 22537
rect 4418 22430 4522 22476
rect 4418 22369 4568 22430
rect 4418 22323 4522 22369
rect 4418 22320 4568 22323
rect 4127 22240 4173 22320
rect 3283 22218 3683 22240
rect 3283 22166 3601 22218
rect 3653 22166 3683 22218
rect 3283 22143 3683 22166
rect 3773 22218 4173 22240
rect 3773 22166 3803 22218
rect 3855 22166 4173 22218
rect 3773 22143 4173 22166
rect 4522 22240 4568 22320
rect 4746 23659 4897 23672
rect 4792 23613 4897 23659
rect 4746 23551 4897 23613
rect 4792 23505 4897 23551
rect 4746 23443 4897 23505
rect 4792 23397 4897 23443
rect 4746 23335 4897 23397
rect 4792 23289 4897 23335
rect 4746 23227 4897 23289
rect 4792 23181 4897 23227
rect 4746 23119 4897 23181
rect 4792 23073 4897 23119
rect 4746 23011 4897 23073
rect 4792 22965 4897 23011
rect 4746 22904 4897 22965
rect 4792 22858 4897 22904
rect 4746 22797 4897 22858
rect 4792 22751 4897 22797
rect 4746 22690 4897 22751
rect 4792 22644 4897 22690
rect 4746 22583 4897 22644
rect 4792 22537 4897 22583
rect 4746 22476 4897 22537
rect 4792 22430 4897 22476
rect 4746 22369 4897 22430
rect 4792 22323 4897 22369
rect 4746 22310 4897 22323
rect 5041 24274 5188 24278
rect 5041 24228 5142 24274
rect 5041 24167 5188 24228
rect 5041 24121 5142 24167
rect 5041 24060 5188 24121
rect 5041 24014 5142 24060
rect 5041 24001 5188 24014
rect 5366 25355 5412 25363
rect 5366 25350 5517 25355
rect 5412 25304 5517 25350
rect 5366 25242 5517 25304
rect 5412 25196 5517 25242
rect 5366 25134 5517 25196
rect 5412 25088 5517 25134
rect 5366 25026 5517 25088
rect 5412 24980 5517 25026
rect 5366 24918 5517 24980
rect 5412 24872 5517 24918
rect 5366 24810 5517 24872
rect 5412 24764 5517 24810
rect 5366 24702 5517 24764
rect 5412 24656 5517 24702
rect 5366 24595 5517 24656
rect 5412 24549 5517 24595
rect 5366 24488 5517 24549
rect 5412 24442 5517 24488
rect 5366 24381 5517 24442
rect 5412 24335 5517 24381
rect 5366 24274 5517 24335
rect 5412 24228 5517 24274
rect 5366 24167 5517 24228
rect 5412 24121 5517 24167
rect 5366 24060 5517 24121
rect 5412 24014 5517 24060
rect 5366 24001 5517 24014
rect 5041 23672 5129 24001
rect 5186 23919 5368 23931
rect 5186 23763 5257 23919
rect 5309 23763 5368 23919
rect 5186 23748 5368 23763
rect 5425 23672 5517 24001
rect 5041 23659 5188 23672
rect 5041 23613 5142 23659
rect 5041 23551 5188 23613
rect 5041 23505 5142 23551
rect 5041 23443 5188 23505
rect 5041 23397 5142 23443
rect 5041 23335 5188 23397
rect 5041 23289 5142 23335
rect 5041 23227 5188 23289
rect 5041 23181 5142 23227
rect 5041 23119 5188 23181
rect 5041 23073 5142 23119
rect 5041 23011 5188 23073
rect 5041 22965 5142 23011
rect 5041 22904 5188 22965
rect 5041 22858 5142 22904
rect 5041 22797 5188 22858
rect 5041 22751 5142 22797
rect 5041 22690 5188 22751
rect 5041 22644 5142 22690
rect 5041 22583 5188 22644
rect 5041 22537 5142 22583
rect 5041 22476 5188 22537
rect 5041 22430 5142 22476
rect 5041 22369 5188 22430
rect 5041 22323 5142 22369
rect 5041 22320 5188 22323
rect 5142 22310 5188 22320
rect 5366 23659 5517 23672
rect 5412 23613 5517 23659
rect 5366 23551 5517 23613
rect 5412 23505 5517 23551
rect 5366 23443 5517 23505
rect 5412 23397 5517 23443
rect 5366 23335 5517 23397
rect 5412 23289 5517 23335
rect 5366 23227 5517 23289
rect 5412 23181 5517 23227
rect 5366 23119 5517 23181
rect 5412 23073 5517 23119
rect 5366 23011 5517 23073
rect 5412 22965 5517 23011
rect 5366 22904 5517 22965
rect 5412 22858 5517 22904
rect 5366 22797 5517 22858
rect 5412 22751 5517 22797
rect 5366 22690 5517 22751
rect 5412 22644 5517 22690
rect 5366 22583 5517 22644
rect 5412 22537 5517 22583
rect 5366 22476 5517 22537
rect 5412 22430 5517 22476
rect 5366 22369 5517 22430
rect 5412 22323 5517 22369
rect 5366 22320 5517 22323
rect 5366 22240 5412 22320
rect 4522 22218 4922 22240
rect 4522 22166 4840 22218
rect 4892 22166 4922 22218
rect 4522 22143 4922 22166
rect 5012 22218 5412 22240
rect 5012 22166 5042 22218
rect 5094 22166 5412 22218
rect 5012 22143 5412 22166
rect 1180 22059 1322 22064
rect 2419 22059 2561 22064
rect 3657 22059 3799 22064
rect 4896 22059 5038 22064
rect 5516 22059 5658 22064
rect 631 22027 5658 22059
rect 631 22020 5327 22027
rect 631 21968 831 22020
rect 883 22013 1619 22020
rect 883 21968 1228 22013
rect 631 21967 1228 21968
rect 1274 21968 1619 22013
rect 1671 21968 2070 22020
rect 2122 22013 2858 22020
rect 2122 21968 2467 22013
rect 1274 21967 2467 21968
rect 2513 21968 2858 22013
rect 2910 21968 3308 22020
rect 3360 22013 4096 22020
rect 3360 21968 3705 22013
rect 2513 21967 3705 21968
rect 3751 21968 4096 22013
rect 4148 21968 4547 22020
rect 4599 22013 5327 22020
rect 4599 21968 4944 22013
rect 3751 21967 4944 21968
rect 4990 21975 5327 22013
rect 5379 22013 5658 22027
rect 5379 21975 5564 22013
rect 4990 21967 5564 21975
rect 5610 21967 5658 22013
rect 631 21925 5658 21967
rect 1180 21916 1322 21925
rect 2419 21916 2561 21925
rect 3657 21916 3799 21925
rect 4896 21916 5038 21925
rect 5516 21916 5658 21925
rect 686 21812 1203 21837
rect 686 21760 699 21812
rect 751 21760 1203 21812
rect 686 21740 1203 21760
rect 1110 21668 1203 21740
rect 806 21660 852 21668
rect 702 21655 852 21660
rect 702 21609 806 21655
rect 702 21547 852 21609
rect 702 21501 806 21547
rect 702 21439 852 21501
rect 702 21393 806 21439
rect 702 21331 852 21393
rect 702 21285 806 21331
rect 702 21223 852 21285
rect 702 21177 806 21223
rect 702 21115 852 21177
rect 702 21069 806 21115
rect 702 21007 852 21069
rect 702 20961 806 21007
rect 702 20900 852 20961
rect 702 20854 806 20900
rect 702 20793 852 20854
rect 702 20747 806 20793
rect 702 20686 852 20747
rect 702 20640 806 20686
rect 702 20579 852 20640
rect 702 20533 806 20579
rect 702 20472 852 20533
rect 702 20426 806 20472
rect 702 20365 852 20426
rect 702 20319 806 20365
rect 702 20306 852 20319
rect 1030 21655 1203 21668
rect 1076 21609 1203 21655
rect 1030 21547 1203 21609
rect 1076 21501 1203 21547
rect 1030 21439 1203 21501
rect 1076 21393 1203 21439
rect 1030 21331 1203 21393
rect 1076 21285 1203 21331
rect 1030 21223 1203 21285
rect 1076 21177 1203 21223
rect 1030 21115 1203 21177
rect 1076 21069 1203 21115
rect 1030 21007 1203 21069
rect 1076 20961 1203 21007
rect 1030 20900 1203 20961
rect 1076 20854 1203 20900
rect 1030 20793 1203 20854
rect 1076 20747 1203 20793
rect 1030 20686 1203 20747
rect 1076 20640 1203 20686
rect 1030 20579 1203 20640
rect 1076 20533 1203 20579
rect 1030 20472 1203 20533
rect 1076 20426 1203 20472
rect 1030 20365 1203 20426
rect 1076 20319 1203 20365
rect 1030 20306 1203 20319
rect 702 19813 772 20306
rect 851 20222 1032 20236
rect 851 20212 918 20222
rect 964 20212 1032 20222
rect 851 20160 913 20212
rect 965 20160 1032 20212
rect 851 20101 1032 20160
rect 851 19948 1032 20021
rect 851 19896 915 19948
rect 967 19896 1032 19948
rect 851 19885 1032 19896
rect 903 19884 979 19885
rect 1110 19813 1203 20306
rect 702 19800 852 19813
rect 702 19754 806 19800
rect 702 19692 852 19754
rect 702 19646 806 19692
rect 702 19584 852 19646
rect 702 19538 806 19584
rect 702 19476 852 19538
rect 702 19430 806 19476
rect 702 19368 852 19430
rect 702 19322 806 19368
rect 702 19260 852 19322
rect 702 19214 806 19260
rect 702 19152 852 19214
rect 702 19106 806 19152
rect 702 19045 852 19106
rect 702 18999 806 19045
rect 702 18938 852 18999
rect 702 18892 806 18938
rect 702 18831 852 18892
rect 702 18785 806 18831
rect 702 18724 852 18785
rect 702 18678 806 18724
rect 702 18617 852 18678
rect 702 18571 806 18617
rect 702 18510 852 18571
rect 702 18464 806 18510
rect 702 18463 852 18464
rect 1030 19800 1203 19813
rect 1076 19754 1203 19800
rect 1030 19692 1203 19754
rect 1076 19646 1203 19692
rect 1030 19584 1203 19646
rect 1076 19538 1203 19584
rect 1030 19476 1203 19538
rect 1076 19430 1203 19476
rect 1030 19368 1203 19430
rect 1076 19322 1203 19368
rect 1030 19260 1203 19322
rect 1076 19214 1203 19260
rect 1030 19152 1203 19214
rect 1076 19106 1203 19152
rect 1030 19045 1203 19106
rect 1076 18999 1203 19045
rect 1030 18938 1203 18999
rect 1076 18892 1203 18938
rect 1030 18831 1203 18892
rect 1076 18785 1203 18831
rect 1030 18724 1203 18785
rect 1076 18678 1203 18724
rect 1030 18617 1203 18678
rect 1076 18571 1203 18617
rect 1030 18510 1203 18571
rect 1076 18464 1203 18510
rect 702 18401 887 18463
rect 1030 18461 1203 18464
rect 1299 21812 1816 21837
rect 1299 21760 1751 21812
rect 1803 21760 1816 21812
rect 1299 21740 1816 21760
rect 1925 21812 2442 21837
rect 1925 21760 1938 21812
rect 1990 21760 2442 21812
rect 1925 21740 2442 21760
rect 1299 21668 1392 21740
rect 2349 21668 2442 21740
rect 1299 21655 1472 21668
rect 1299 21609 1426 21655
rect 1299 21547 1472 21609
rect 1299 21501 1426 21547
rect 1299 21439 1472 21501
rect 1299 21393 1426 21439
rect 1299 21331 1472 21393
rect 1299 21285 1426 21331
rect 1299 21223 1472 21285
rect 1299 21177 1426 21223
rect 1299 21115 1472 21177
rect 1299 21069 1426 21115
rect 1299 21007 1472 21069
rect 1299 20961 1426 21007
rect 1299 20900 1472 20961
rect 1299 20854 1426 20900
rect 1299 20793 1472 20854
rect 1299 20747 1426 20793
rect 1299 20686 1472 20747
rect 1299 20640 1426 20686
rect 1299 20579 1472 20640
rect 1299 20533 1426 20579
rect 1299 20472 1472 20533
rect 1299 20426 1426 20472
rect 1299 20365 1472 20426
rect 1299 20319 1426 20365
rect 1299 20306 1472 20319
rect 1650 21660 1696 21668
rect 2045 21660 2091 21668
rect 1650 21655 1800 21660
rect 1696 21609 1800 21655
rect 1650 21547 1800 21609
rect 1696 21501 1800 21547
rect 1650 21439 1800 21501
rect 1696 21393 1800 21439
rect 1650 21331 1800 21393
rect 1696 21285 1800 21331
rect 1650 21223 1800 21285
rect 1696 21177 1800 21223
rect 1650 21115 1800 21177
rect 1696 21069 1800 21115
rect 1650 21007 1800 21069
rect 1696 20961 1800 21007
rect 1650 20900 1800 20961
rect 1696 20854 1800 20900
rect 1650 20793 1800 20854
rect 1696 20747 1800 20793
rect 1650 20686 1800 20747
rect 1696 20640 1800 20686
rect 1650 20579 1800 20640
rect 1696 20533 1800 20579
rect 1650 20472 1800 20533
rect 1696 20426 1800 20472
rect 1650 20365 1800 20426
rect 1696 20319 1800 20365
rect 1650 20306 1800 20319
rect 1299 19813 1392 20306
rect 1470 20222 1651 20236
rect 1470 20212 1538 20222
rect 1584 20212 1651 20222
rect 1470 20160 1537 20212
rect 1589 20160 1651 20212
rect 1470 20101 1651 20160
rect 1470 19948 1651 20021
rect 1470 19896 1535 19948
rect 1587 19896 1651 19948
rect 1470 19885 1651 19896
rect 1523 19884 1599 19885
rect 1730 19813 1800 20306
rect 1299 19800 1472 19813
rect 1299 19754 1426 19800
rect 1299 19692 1472 19754
rect 1299 19646 1426 19692
rect 1299 19584 1472 19646
rect 1299 19538 1426 19584
rect 1299 19476 1472 19538
rect 1299 19430 1426 19476
rect 1299 19368 1472 19430
rect 1299 19322 1426 19368
rect 1299 19260 1472 19322
rect 1299 19214 1426 19260
rect 1299 19152 1472 19214
rect 1299 19106 1426 19152
rect 1299 19045 1472 19106
rect 1299 18999 1426 19045
rect 1299 18938 1472 18999
rect 1299 18892 1426 18938
rect 1299 18831 1472 18892
rect 1299 18785 1426 18831
rect 1299 18724 1472 18785
rect 1299 18678 1426 18724
rect 1299 18617 1472 18678
rect 1299 18571 1426 18617
rect 1299 18510 1472 18571
rect 1299 18464 1426 18510
rect 1299 18461 1472 18464
rect 1650 19800 1800 19813
rect 1696 19754 1800 19800
rect 1650 19692 1800 19754
rect 1696 19646 1800 19692
rect 1650 19584 1800 19646
rect 1696 19538 1800 19584
rect 1650 19476 1800 19538
rect 1696 19430 1800 19476
rect 1650 19368 1800 19430
rect 1696 19322 1800 19368
rect 1650 19260 1800 19322
rect 1696 19214 1800 19260
rect 1650 19152 1800 19214
rect 1696 19106 1800 19152
rect 1650 19045 1800 19106
rect 1696 18999 1800 19045
rect 1650 18938 1800 18999
rect 1696 18892 1800 18938
rect 1650 18831 1800 18892
rect 1696 18785 1800 18831
rect 1650 18724 1800 18785
rect 1696 18678 1800 18724
rect 1650 18617 1800 18678
rect 1696 18571 1800 18617
rect 1650 18510 1800 18571
rect 1696 18464 1800 18510
rect 1650 18463 1800 18464
rect 1030 18451 1076 18461
rect 1426 18451 1472 18461
rect 698 18380 887 18401
rect 698 18328 734 18380
rect 786 18328 887 18380
rect 698 18308 887 18328
rect 702 18307 887 18308
rect 1615 18400 1800 18463
rect 1941 21655 2091 21660
rect 1941 21609 2045 21655
rect 1941 21547 2091 21609
rect 1941 21501 2045 21547
rect 1941 21439 2091 21501
rect 1941 21393 2045 21439
rect 1941 21331 2091 21393
rect 1941 21285 2045 21331
rect 1941 21223 2091 21285
rect 1941 21177 2045 21223
rect 1941 21115 2091 21177
rect 1941 21069 2045 21115
rect 1941 21007 2091 21069
rect 1941 20961 2045 21007
rect 1941 20900 2091 20961
rect 1941 20854 2045 20900
rect 1941 20793 2091 20854
rect 1941 20747 2045 20793
rect 1941 20686 2091 20747
rect 1941 20640 2045 20686
rect 1941 20579 2091 20640
rect 1941 20533 2045 20579
rect 1941 20472 2091 20533
rect 1941 20426 2045 20472
rect 1941 20365 2091 20426
rect 1941 20319 2045 20365
rect 1941 20306 2091 20319
rect 2269 21655 2442 21668
rect 2315 21609 2442 21655
rect 2269 21547 2442 21609
rect 2315 21501 2442 21547
rect 2269 21439 2442 21501
rect 2315 21393 2442 21439
rect 2269 21331 2442 21393
rect 2315 21285 2442 21331
rect 2269 21223 2442 21285
rect 2315 21177 2442 21223
rect 2269 21115 2442 21177
rect 2315 21069 2442 21115
rect 2269 21007 2442 21069
rect 2315 20961 2442 21007
rect 2269 20900 2442 20961
rect 2315 20854 2442 20900
rect 2269 20793 2442 20854
rect 2315 20747 2442 20793
rect 2269 20686 2442 20747
rect 2315 20640 2442 20686
rect 2269 20579 2442 20640
rect 2315 20533 2442 20579
rect 2269 20472 2442 20533
rect 2315 20426 2442 20472
rect 2269 20365 2442 20426
rect 2315 20319 2442 20365
rect 2269 20306 2442 20319
rect 1941 19813 2011 20306
rect 2090 20222 2271 20236
rect 2090 20212 2157 20222
rect 2203 20212 2271 20222
rect 2090 20160 2152 20212
rect 2204 20160 2271 20212
rect 2090 20101 2271 20160
rect 2090 19948 2271 20021
rect 2090 19896 2154 19948
rect 2206 19896 2271 19948
rect 2090 19885 2271 19896
rect 2142 19884 2218 19885
rect 2349 19813 2442 20306
rect 1941 19800 2091 19813
rect 1941 19754 2045 19800
rect 1941 19692 2091 19754
rect 1941 19646 2045 19692
rect 1941 19584 2091 19646
rect 1941 19538 2045 19584
rect 1941 19476 2091 19538
rect 1941 19430 2045 19476
rect 1941 19368 2091 19430
rect 1941 19322 2045 19368
rect 1941 19260 2091 19322
rect 1941 19214 2045 19260
rect 1941 19152 2091 19214
rect 1941 19106 2045 19152
rect 1941 19045 2091 19106
rect 1941 18999 2045 19045
rect 1941 18938 2091 18999
rect 1941 18892 2045 18938
rect 1941 18831 2091 18892
rect 1941 18785 2045 18831
rect 1941 18724 2091 18785
rect 1941 18678 2045 18724
rect 1941 18617 2091 18678
rect 1941 18571 2045 18617
rect 1941 18510 2091 18571
rect 1941 18464 2045 18510
rect 1941 18463 2091 18464
rect 2269 19800 2442 19813
rect 2315 19754 2442 19800
rect 2269 19692 2442 19754
rect 2315 19646 2442 19692
rect 2269 19584 2442 19646
rect 2315 19538 2442 19584
rect 2269 19476 2442 19538
rect 2315 19430 2442 19476
rect 2269 19368 2442 19430
rect 2315 19322 2442 19368
rect 2269 19260 2442 19322
rect 2315 19214 2442 19260
rect 2269 19152 2442 19214
rect 2315 19106 2442 19152
rect 2269 19045 2442 19106
rect 2315 18999 2442 19045
rect 2269 18938 2442 18999
rect 2315 18892 2442 18938
rect 2269 18831 2442 18892
rect 2315 18785 2442 18831
rect 2269 18724 2442 18785
rect 2315 18678 2442 18724
rect 2269 18617 2442 18678
rect 2315 18571 2442 18617
rect 2269 18510 2442 18571
rect 2315 18464 2442 18510
rect 1941 18400 2126 18463
rect 2269 18461 2442 18464
rect 2538 21812 3055 21837
rect 2538 21760 2990 21812
rect 3042 21760 3055 21812
rect 2538 21740 3055 21760
rect 3163 21812 3680 21837
rect 3163 21760 3176 21812
rect 3228 21760 3680 21812
rect 3163 21740 3680 21760
rect 2538 21668 2631 21740
rect 3587 21668 3680 21740
rect 2538 21655 2711 21668
rect 2538 21609 2665 21655
rect 2538 21547 2711 21609
rect 2538 21501 2665 21547
rect 2538 21439 2711 21501
rect 2538 21393 2665 21439
rect 2538 21331 2711 21393
rect 2538 21285 2665 21331
rect 2538 21223 2711 21285
rect 2538 21177 2665 21223
rect 2538 21115 2711 21177
rect 2538 21069 2665 21115
rect 2538 21007 2711 21069
rect 2538 20961 2665 21007
rect 2538 20900 2711 20961
rect 2538 20854 2665 20900
rect 2538 20793 2711 20854
rect 2538 20747 2665 20793
rect 2538 20686 2711 20747
rect 2538 20640 2665 20686
rect 2538 20579 2711 20640
rect 2538 20533 2665 20579
rect 2538 20472 2711 20533
rect 2538 20426 2665 20472
rect 2538 20365 2711 20426
rect 2538 20319 2665 20365
rect 2538 20306 2711 20319
rect 2889 21660 2935 21668
rect 3283 21660 3329 21668
rect 2889 21655 3039 21660
rect 2935 21609 3039 21655
rect 2889 21547 3039 21609
rect 2935 21501 3039 21547
rect 2889 21439 3039 21501
rect 2935 21393 3039 21439
rect 2889 21331 3039 21393
rect 2935 21285 3039 21331
rect 2889 21223 3039 21285
rect 2935 21177 3039 21223
rect 2889 21115 3039 21177
rect 2935 21069 3039 21115
rect 2889 21007 3039 21069
rect 2935 20961 3039 21007
rect 2889 20900 3039 20961
rect 2935 20854 3039 20900
rect 2889 20793 3039 20854
rect 2935 20747 3039 20793
rect 2889 20686 3039 20747
rect 2935 20640 3039 20686
rect 2889 20579 3039 20640
rect 2935 20533 3039 20579
rect 2889 20472 3039 20533
rect 2935 20426 3039 20472
rect 2889 20365 3039 20426
rect 2935 20319 3039 20365
rect 2889 20306 3039 20319
rect 2538 19813 2631 20306
rect 2709 20222 2890 20236
rect 2709 20212 2777 20222
rect 2823 20212 2890 20222
rect 2709 20160 2776 20212
rect 2828 20160 2890 20212
rect 2709 20101 2890 20160
rect 2709 19948 2890 20021
rect 2709 19896 2774 19948
rect 2826 19896 2890 19948
rect 2709 19885 2890 19896
rect 2762 19884 2838 19885
rect 2969 19813 3039 20306
rect 2538 19800 2711 19813
rect 2538 19754 2665 19800
rect 2538 19692 2711 19754
rect 2538 19646 2665 19692
rect 2538 19584 2711 19646
rect 2538 19538 2665 19584
rect 2538 19476 2711 19538
rect 2538 19430 2665 19476
rect 2538 19368 2711 19430
rect 2538 19322 2665 19368
rect 2538 19260 2711 19322
rect 2538 19214 2665 19260
rect 2538 19152 2711 19214
rect 2538 19106 2665 19152
rect 2538 19045 2711 19106
rect 2538 18999 2665 19045
rect 2538 18938 2711 18999
rect 2538 18892 2665 18938
rect 2538 18831 2711 18892
rect 2538 18785 2665 18831
rect 2538 18724 2711 18785
rect 2538 18678 2665 18724
rect 2538 18617 2711 18678
rect 2538 18571 2665 18617
rect 2538 18510 2711 18571
rect 2538 18464 2665 18510
rect 2538 18461 2711 18464
rect 2889 19800 3039 19813
rect 2935 19754 3039 19800
rect 2889 19692 3039 19754
rect 2935 19646 3039 19692
rect 2889 19584 3039 19646
rect 2935 19538 3039 19584
rect 2889 19476 3039 19538
rect 2935 19430 3039 19476
rect 2889 19368 3039 19430
rect 2935 19322 3039 19368
rect 2889 19260 3039 19322
rect 2935 19214 3039 19260
rect 2889 19152 3039 19214
rect 2935 19106 3039 19152
rect 2889 19045 3039 19106
rect 2935 18999 3039 19045
rect 2889 18938 3039 18999
rect 2935 18892 3039 18938
rect 2889 18831 3039 18892
rect 2935 18785 3039 18831
rect 2889 18724 3039 18785
rect 2935 18678 3039 18724
rect 2889 18617 3039 18678
rect 2935 18571 3039 18617
rect 2889 18510 3039 18571
rect 2935 18464 3039 18510
rect 2889 18463 3039 18464
rect 2269 18451 2315 18461
rect 2665 18451 2711 18461
rect 1615 18380 2126 18400
rect 1615 18328 1747 18380
rect 1799 18328 1933 18380
rect 1985 18328 2126 18380
rect 1615 18308 2126 18328
rect 1615 18307 1800 18308
rect 1941 18307 2126 18308
rect 2854 18400 3039 18463
rect 3179 21655 3329 21660
rect 3179 21609 3283 21655
rect 3179 21547 3329 21609
rect 3179 21501 3283 21547
rect 3179 21439 3329 21501
rect 3179 21393 3283 21439
rect 3179 21331 3329 21393
rect 3179 21285 3283 21331
rect 3179 21223 3329 21285
rect 3179 21177 3283 21223
rect 3179 21115 3329 21177
rect 3179 21069 3283 21115
rect 3179 21007 3329 21069
rect 3179 20961 3283 21007
rect 3179 20900 3329 20961
rect 3179 20854 3283 20900
rect 3179 20793 3329 20854
rect 3179 20747 3283 20793
rect 3179 20686 3329 20747
rect 3179 20640 3283 20686
rect 3179 20579 3329 20640
rect 3179 20533 3283 20579
rect 3179 20472 3329 20533
rect 3179 20426 3283 20472
rect 3179 20365 3329 20426
rect 3179 20319 3283 20365
rect 3179 20306 3329 20319
rect 3507 21655 3680 21668
rect 3553 21609 3680 21655
rect 3507 21547 3680 21609
rect 3553 21501 3680 21547
rect 3507 21439 3680 21501
rect 3553 21393 3680 21439
rect 3507 21331 3680 21393
rect 3553 21285 3680 21331
rect 3507 21223 3680 21285
rect 3553 21177 3680 21223
rect 3507 21115 3680 21177
rect 3553 21069 3680 21115
rect 3507 21007 3680 21069
rect 3553 20961 3680 21007
rect 3507 20900 3680 20961
rect 3553 20854 3680 20900
rect 3507 20793 3680 20854
rect 3553 20747 3680 20793
rect 3507 20686 3680 20747
rect 3553 20640 3680 20686
rect 3507 20579 3680 20640
rect 3553 20533 3680 20579
rect 3507 20472 3680 20533
rect 3553 20426 3680 20472
rect 3507 20365 3680 20426
rect 3553 20319 3680 20365
rect 3507 20306 3680 20319
rect 3179 19813 3249 20306
rect 3328 20222 3509 20236
rect 3328 20212 3395 20222
rect 3441 20212 3509 20222
rect 3328 20160 3390 20212
rect 3442 20160 3509 20212
rect 3328 20101 3509 20160
rect 3328 19948 3509 20021
rect 3328 19896 3392 19948
rect 3444 19896 3509 19948
rect 3328 19885 3509 19896
rect 3380 19884 3456 19885
rect 3587 19813 3680 20306
rect 3179 19800 3329 19813
rect 3179 19754 3283 19800
rect 3179 19692 3329 19754
rect 3179 19646 3283 19692
rect 3179 19584 3329 19646
rect 3179 19538 3283 19584
rect 3179 19476 3329 19538
rect 3179 19430 3283 19476
rect 3179 19368 3329 19430
rect 3179 19322 3283 19368
rect 3179 19260 3329 19322
rect 3179 19214 3283 19260
rect 3179 19152 3329 19214
rect 3179 19106 3283 19152
rect 3179 19045 3329 19106
rect 3179 18999 3283 19045
rect 3179 18938 3329 18999
rect 3179 18892 3283 18938
rect 3179 18831 3329 18892
rect 3179 18785 3283 18831
rect 3179 18724 3329 18785
rect 3179 18678 3283 18724
rect 3179 18617 3329 18678
rect 3179 18571 3283 18617
rect 3179 18510 3329 18571
rect 3179 18464 3283 18510
rect 3179 18463 3329 18464
rect 3507 19800 3680 19813
rect 3553 19754 3680 19800
rect 3507 19692 3680 19754
rect 3553 19646 3680 19692
rect 3507 19584 3680 19646
rect 3553 19538 3680 19584
rect 3507 19476 3680 19538
rect 3553 19430 3680 19476
rect 3507 19368 3680 19430
rect 3553 19322 3680 19368
rect 3507 19260 3680 19322
rect 3553 19214 3680 19260
rect 3507 19152 3680 19214
rect 3553 19106 3680 19152
rect 3507 19045 3680 19106
rect 3553 18999 3680 19045
rect 3507 18938 3680 18999
rect 3553 18892 3680 18938
rect 3507 18831 3680 18892
rect 3553 18785 3680 18831
rect 3507 18724 3680 18785
rect 3553 18678 3680 18724
rect 3507 18617 3680 18678
rect 3553 18571 3680 18617
rect 3507 18510 3680 18571
rect 3553 18464 3680 18510
rect 3179 18400 3364 18463
rect 3507 18461 3680 18464
rect 3776 21812 4293 21837
rect 3776 21760 4228 21812
rect 4280 21760 4293 21812
rect 3776 21740 4293 21760
rect 4402 21812 4919 21837
rect 4402 21760 4415 21812
rect 4467 21760 4919 21812
rect 4402 21740 4919 21760
rect 3776 21668 3869 21740
rect 4826 21668 4919 21740
rect 3776 21655 3949 21668
rect 3776 21609 3903 21655
rect 3776 21547 3949 21609
rect 3776 21501 3903 21547
rect 3776 21439 3949 21501
rect 3776 21393 3903 21439
rect 3776 21331 3949 21393
rect 3776 21285 3903 21331
rect 3776 21223 3949 21285
rect 3776 21177 3903 21223
rect 3776 21115 3949 21177
rect 3776 21069 3903 21115
rect 3776 21007 3949 21069
rect 3776 20961 3903 21007
rect 3776 20900 3949 20961
rect 3776 20854 3903 20900
rect 3776 20793 3949 20854
rect 3776 20747 3903 20793
rect 3776 20686 3949 20747
rect 3776 20640 3903 20686
rect 3776 20579 3949 20640
rect 3776 20533 3903 20579
rect 3776 20472 3949 20533
rect 3776 20426 3903 20472
rect 3776 20365 3949 20426
rect 3776 20319 3903 20365
rect 3776 20306 3949 20319
rect 4127 21660 4173 21668
rect 4522 21660 4568 21668
rect 4127 21655 4277 21660
rect 4173 21609 4277 21655
rect 4127 21547 4277 21609
rect 4173 21501 4277 21547
rect 4127 21439 4277 21501
rect 4173 21393 4277 21439
rect 4127 21331 4277 21393
rect 4173 21285 4277 21331
rect 4127 21223 4277 21285
rect 4173 21177 4277 21223
rect 4127 21115 4277 21177
rect 4173 21069 4277 21115
rect 4127 21007 4277 21069
rect 4173 20961 4277 21007
rect 4127 20900 4277 20961
rect 4173 20854 4277 20900
rect 4127 20793 4277 20854
rect 4173 20747 4277 20793
rect 4127 20686 4277 20747
rect 4173 20640 4277 20686
rect 4127 20579 4277 20640
rect 4173 20533 4277 20579
rect 4127 20472 4277 20533
rect 4173 20426 4277 20472
rect 4127 20365 4277 20426
rect 4173 20319 4277 20365
rect 4127 20306 4277 20319
rect 3776 19813 3869 20306
rect 3947 20222 4128 20236
rect 3947 20212 4015 20222
rect 4061 20212 4128 20222
rect 3947 20160 4014 20212
rect 4066 20160 4128 20212
rect 3947 20101 4128 20160
rect 3947 19948 4128 20021
rect 3947 19896 4012 19948
rect 4064 19896 4128 19948
rect 3947 19885 4128 19896
rect 4000 19884 4076 19885
rect 4207 19813 4277 20306
rect 3776 19800 3949 19813
rect 3776 19754 3903 19800
rect 3776 19692 3949 19754
rect 3776 19646 3903 19692
rect 3776 19584 3949 19646
rect 3776 19538 3903 19584
rect 3776 19476 3949 19538
rect 3776 19430 3903 19476
rect 3776 19368 3949 19430
rect 3776 19322 3903 19368
rect 3776 19260 3949 19322
rect 3776 19214 3903 19260
rect 3776 19152 3949 19214
rect 3776 19106 3903 19152
rect 3776 19045 3949 19106
rect 3776 18999 3903 19045
rect 3776 18938 3949 18999
rect 3776 18892 3903 18938
rect 3776 18831 3949 18892
rect 3776 18785 3903 18831
rect 3776 18724 3949 18785
rect 3776 18678 3903 18724
rect 3776 18617 3949 18678
rect 3776 18571 3903 18617
rect 3776 18510 3949 18571
rect 3776 18464 3903 18510
rect 3776 18461 3949 18464
rect 4127 19800 4277 19813
rect 4173 19754 4277 19800
rect 4127 19692 4277 19754
rect 4173 19646 4277 19692
rect 4127 19584 4277 19646
rect 4173 19538 4277 19584
rect 4127 19476 4277 19538
rect 4173 19430 4277 19476
rect 4127 19368 4277 19430
rect 4173 19322 4277 19368
rect 4127 19260 4277 19322
rect 4173 19214 4277 19260
rect 4127 19152 4277 19214
rect 4173 19106 4277 19152
rect 4127 19045 4277 19106
rect 4173 18999 4277 19045
rect 4127 18938 4277 18999
rect 4173 18892 4277 18938
rect 4127 18831 4277 18892
rect 4173 18785 4277 18831
rect 4127 18724 4277 18785
rect 4173 18678 4277 18724
rect 4127 18617 4277 18678
rect 4173 18571 4277 18617
rect 4127 18510 4277 18571
rect 4173 18464 4277 18510
rect 4127 18463 4277 18464
rect 3507 18451 3553 18461
rect 3903 18451 3949 18461
rect 2854 18380 3364 18400
rect 2854 18328 2985 18380
rect 3037 18328 3171 18380
rect 3223 18328 3364 18380
rect 2854 18308 3364 18328
rect 2854 18307 3039 18308
rect 3179 18307 3364 18308
rect 4092 18400 4277 18463
rect 4418 21655 4568 21660
rect 4418 21609 4522 21655
rect 4418 21547 4568 21609
rect 4418 21501 4522 21547
rect 4418 21439 4568 21501
rect 4418 21393 4522 21439
rect 4418 21331 4568 21393
rect 4418 21285 4522 21331
rect 4418 21223 4568 21285
rect 4418 21177 4522 21223
rect 4418 21115 4568 21177
rect 4418 21069 4522 21115
rect 4418 21007 4568 21069
rect 4418 20961 4522 21007
rect 4418 20900 4568 20961
rect 4418 20854 4522 20900
rect 4418 20793 4568 20854
rect 4418 20747 4522 20793
rect 4418 20686 4568 20747
rect 4418 20640 4522 20686
rect 4418 20579 4568 20640
rect 4418 20533 4522 20579
rect 4418 20472 4568 20533
rect 4418 20426 4522 20472
rect 4418 20365 4568 20426
rect 4418 20319 4522 20365
rect 4418 20306 4568 20319
rect 4746 21655 4919 21668
rect 4792 21609 4919 21655
rect 4746 21547 4919 21609
rect 4792 21501 4919 21547
rect 4746 21439 4919 21501
rect 4792 21393 4919 21439
rect 4746 21331 4919 21393
rect 4792 21285 4919 21331
rect 4746 21223 4919 21285
rect 4792 21177 4919 21223
rect 4746 21115 4919 21177
rect 4792 21069 4919 21115
rect 4746 21007 4919 21069
rect 4792 20961 4919 21007
rect 4746 20900 4919 20961
rect 4792 20854 4919 20900
rect 4746 20793 4919 20854
rect 4792 20747 4919 20793
rect 4746 20686 4919 20747
rect 4792 20640 4919 20686
rect 4746 20579 4919 20640
rect 4792 20533 4919 20579
rect 4746 20472 4919 20533
rect 4792 20426 4919 20472
rect 4746 20365 4919 20426
rect 4792 20319 4919 20365
rect 4746 20306 4919 20319
rect 4418 19813 4488 20306
rect 4567 20222 4748 20236
rect 4567 20212 4634 20222
rect 4680 20212 4748 20222
rect 4567 20160 4629 20212
rect 4681 20160 4748 20212
rect 4567 20101 4748 20160
rect 4567 19948 4748 20021
rect 4567 19896 4631 19948
rect 4683 19896 4748 19948
rect 4567 19885 4748 19896
rect 4619 19884 4695 19885
rect 4826 19813 4919 20306
rect 4418 19800 4568 19813
rect 4418 19754 4522 19800
rect 4418 19692 4568 19754
rect 4418 19646 4522 19692
rect 4418 19584 4568 19646
rect 4418 19538 4522 19584
rect 4418 19476 4568 19538
rect 4418 19430 4522 19476
rect 4418 19368 4568 19430
rect 4418 19322 4522 19368
rect 4418 19260 4568 19322
rect 4418 19214 4522 19260
rect 4418 19152 4568 19214
rect 4418 19106 4522 19152
rect 4418 19045 4568 19106
rect 4418 18999 4522 19045
rect 4418 18938 4568 18999
rect 4418 18892 4522 18938
rect 4418 18831 4568 18892
rect 4418 18785 4522 18831
rect 4418 18724 4568 18785
rect 4418 18678 4522 18724
rect 4418 18617 4568 18678
rect 4418 18571 4522 18617
rect 4418 18510 4568 18571
rect 4418 18464 4522 18510
rect 4418 18463 4568 18464
rect 4746 19800 4919 19813
rect 4792 19754 4919 19800
rect 4746 19692 4919 19754
rect 4792 19646 4919 19692
rect 4746 19584 4919 19646
rect 4792 19538 4919 19584
rect 4746 19476 4919 19538
rect 4792 19430 4919 19476
rect 4746 19368 4919 19430
rect 4792 19322 4919 19368
rect 4746 19260 4919 19322
rect 4792 19214 4919 19260
rect 4746 19152 4919 19214
rect 4792 19106 4919 19152
rect 4746 19045 4919 19106
rect 4792 18999 4919 19045
rect 4746 18938 4919 18999
rect 4792 18892 4919 18938
rect 4746 18831 4919 18892
rect 4792 18785 4919 18831
rect 4746 18724 4919 18785
rect 4792 18678 4919 18724
rect 4746 18617 4919 18678
rect 4792 18571 4919 18617
rect 4746 18510 4919 18571
rect 4792 18464 4919 18510
rect 4418 18400 4603 18463
rect 4746 18461 4919 18464
rect 5015 21811 5528 21837
rect 5015 21759 5459 21811
rect 5511 21759 5528 21811
rect 5015 21740 5528 21759
rect 5015 21668 5155 21740
rect 5015 21655 5188 21668
rect 5015 21609 5142 21655
rect 5015 21547 5188 21609
rect 5015 21501 5142 21547
rect 5015 21439 5188 21501
rect 5015 21393 5142 21439
rect 5015 21331 5188 21393
rect 5015 21285 5142 21331
rect 5015 21223 5188 21285
rect 5015 21177 5142 21223
rect 5015 21115 5188 21177
rect 5015 21069 5142 21115
rect 5015 21007 5188 21069
rect 5015 20961 5142 21007
rect 5015 20900 5188 20961
rect 5015 20854 5142 20900
rect 5015 20793 5188 20854
rect 5015 20747 5142 20793
rect 5015 20686 5188 20747
rect 5015 20640 5142 20686
rect 5015 20579 5188 20640
rect 5015 20533 5142 20579
rect 5015 20472 5188 20533
rect 5015 20426 5142 20472
rect 5015 20365 5188 20426
rect 5015 20319 5142 20365
rect 5015 20306 5188 20319
rect 5366 21660 5412 21668
rect 5366 21655 5517 21660
rect 5412 21609 5517 21655
rect 5366 21547 5517 21609
rect 5412 21501 5517 21547
rect 5366 21439 5517 21501
rect 5412 21393 5517 21439
rect 5366 21331 5517 21393
rect 5412 21285 5517 21331
rect 5366 21223 5517 21285
rect 5412 21177 5517 21223
rect 5366 21115 5517 21177
rect 5412 21069 5517 21115
rect 5366 21007 5517 21069
rect 5412 20961 5517 21007
rect 5366 20900 5517 20961
rect 5412 20854 5517 20900
rect 5366 20793 5517 20854
rect 5412 20747 5517 20793
rect 5366 20686 5517 20747
rect 5412 20640 5517 20686
rect 5366 20579 5517 20640
rect 5412 20533 5517 20579
rect 5366 20472 5517 20533
rect 5412 20426 5517 20472
rect 5366 20365 5517 20426
rect 5412 20319 5517 20365
rect 5366 20306 5517 20319
rect 5015 19813 5112 20306
rect 5186 20222 5368 20236
rect 5186 20212 5254 20222
rect 5300 20212 5368 20222
rect 5186 20160 5253 20212
rect 5305 20160 5368 20212
rect 5186 20101 5368 20160
rect 5186 19949 5368 20021
rect 5186 19897 5251 19949
rect 5303 19897 5368 19949
rect 5186 19885 5368 19897
rect 5431 19813 5517 20306
rect 5015 19800 5188 19813
rect 5015 19754 5142 19800
rect 5015 19692 5188 19754
rect 5015 19646 5142 19692
rect 5015 19584 5188 19646
rect 5015 19538 5142 19584
rect 5015 19476 5188 19538
rect 5015 19430 5142 19476
rect 5015 19368 5188 19430
rect 5015 19322 5142 19368
rect 5015 19260 5188 19322
rect 5015 19214 5142 19260
rect 5015 19152 5188 19214
rect 5015 19106 5142 19152
rect 5015 19045 5188 19106
rect 5015 18999 5142 19045
rect 5015 18938 5188 18999
rect 5015 18892 5142 18938
rect 5015 18831 5188 18892
rect 5015 18785 5142 18831
rect 5015 18724 5188 18785
rect 5015 18678 5142 18724
rect 5015 18617 5188 18678
rect 5015 18571 5142 18617
rect 5015 18510 5188 18571
rect 5015 18464 5142 18510
rect 5015 18461 5188 18464
rect 4746 18451 4792 18461
rect 5142 18451 5188 18461
rect 5366 19800 5517 19813
rect 5412 19754 5517 19800
rect 5366 19692 5517 19754
rect 5412 19646 5517 19692
rect 5366 19584 5517 19646
rect 5412 19538 5517 19584
rect 5366 19476 5517 19538
rect 5412 19430 5517 19476
rect 5366 19368 5517 19430
rect 5412 19322 5517 19368
rect 5366 19260 5517 19322
rect 5412 19214 5517 19260
rect 5366 19152 5517 19214
rect 5412 19106 5517 19152
rect 5366 19045 5517 19106
rect 5412 18999 5517 19045
rect 5366 18938 5517 18999
rect 5412 18892 5517 18938
rect 5366 18831 5517 18892
rect 5412 18785 5517 18831
rect 5366 18724 5517 18785
rect 5412 18678 5517 18724
rect 5366 18617 5517 18678
rect 5412 18571 5517 18617
rect 5366 18510 5517 18571
rect 5412 18464 5517 18510
rect 5366 18451 5517 18464
rect 4092 18380 4603 18400
rect 4092 18328 4224 18380
rect 4276 18328 4410 18380
rect 4462 18328 4603 18380
rect 4092 18308 4603 18328
rect 4092 18307 4277 18308
rect 4418 18307 4603 18308
rect 5388 18380 5517 18451
rect 5388 18328 5429 18380
rect 5481 18328 5517 18380
rect 5388 18307 5517 18328
rect 631 18171 5587 18205
rect 631 18168 1699 18171
rect 631 18122 754 18168
rect 800 18122 912 18168
rect 958 18122 1070 18168
rect 1116 18122 1228 18168
rect 1274 18122 1386 18168
rect 1432 18122 1544 18168
rect 1590 18122 1699 18168
rect 631 18119 1699 18122
rect 1751 18119 1990 18171
rect 2042 18168 2938 18171
rect 2042 18122 2151 18168
rect 2197 18122 2309 18168
rect 2355 18122 2467 18168
rect 2513 18122 2625 18168
rect 2671 18122 2783 18168
rect 2829 18122 2938 18168
rect 2042 18119 2938 18122
rect 2990 18119 3229 18171
rect 3281 18168 4176 18171
rect 3281 18122 3389 18168
rect 3435 18122 3547 18168
rect 3593 18122 3705 18168
rect 3751 18122 3863 18168
rect 3909 18122 4021 18168
rect 4067 18122 4176 18168
rect 3281 18119 4176 18122
rect 4228 18119 4467 18171
rect 4519 18168 5587 18171
rect 4519 18122 4628 18168
rect 4674 18122 4786 18168
rect 4832 18122 4944 18168
rect 4990 18122 5102 18168
rect 5148 18122 5260 18168
rect 5306 18122 5418 18168
rect 5464 18122 5587 18168
rect 4519 18119 5587 18122
rect 631 18085 5587 18119
rect 631 17829 702 18085
rect 847 17980 1115 18005
rect 847 17928 913 17980
rect 965 17978 1115 17980
rect 965 17932 975 17978
rect 1021 17932 1115 17978
rect 965 17928 1115 17932
rect 847 17908 1115 17928
rect 631 17713 805 17829
rect 631 17667 725 17713
rect 771 17667 805 17713
rect 631 17550 805 17667
rect 948 17817 1056 17829
rect 948 17661 973 17817
rect 1025 17661 1056 17817
rect 510 17253 578 17256
rect 510 17245 826 17253
rect 510 17105 521 17245
rect 567 17216 826 17245
rect 567 17170 780 17216
rect 567 17105 826 17170
rect 948 17216 1056 17661
rect 1194 17713 1308 18085
rect 1387 17980 1655 18005
rect 1387 17978 1537 17980
rect 1387 17932 1481 17978
rect 1527 17932 1537 17978
rect 1387 17928 1537 17932
rect 1589 17928 1655 17980
rect 1387 17908 1655 17928
rect 1800 17829 1941 18085
rect 2086 17980 2354 18005
rect 2086 17928 2152 17980
rect 2204 17978 2354 17980
rect 2204 17932 2214 17978
rect 2260 17932 2354 17978
rect 2204 17928 2354 17932
rect 2086 17908 2354 17928
rect 1194 17667 1228 17713
rect 1274 17667 1308 17713
rect 1194 17550 1308 17667
rect 1446 17817 1554 17829
rect 1446 17661 1477 17817
rect 1529 17661 1554 17817
rect 948 17170 1004 17216
rect 1050 17170 1056 17216
rect 948 17133 1056 17170
rect 1194 17216 1308 17253
rect 1194 17170 1228 17216
rect 1274 17170 1308 17216
rect 510 17024 826 17105
rect 1194 17024 1308 17170
rect 1446 17216 1554 17661
rect 1697 17713 2044 17829
rect 1697 17667 1731 17713
rect 1777 17667 1964 17713
rect 2010 17667 2044 17713
rect 1697 17550 2044 17667
rect 2187 17817 2295 17829
rect 2187 17661 2212 17817
rect 2264 17661 2295 17817
rect 1837 17253 1905 17256
rect 1446 17170 1452 17216
rect 1498 17170 1554 17216
rect 1446 17133 1554 17170
rect 1676 17245 2065 17253
rect 1676 17216 1848 17245
rect 1722 17170 1848 17216
rect 1676 17105 1848 17170
rect 1894 17216 2065 17245
rect 1894 17170 2019 17216
rect 1894 17105 2065 17170
rect 2187 17216 2295 17661
rect 2433 17713 2547 18085
rect 2626 17980 2894 18005
rect 2626 17978 2776 17980
rect 2626 17932 2720 17978
rect 2766 17932 2776 17978
rect 2626 17928 2776 17932
rect 2828 17928 2894 17980
rect 2626 17908 2894 17928
rect 3039 17829 3179 18085
rect 3324 17980 3592 18005
rect 3324 17928 3390 17980
rect 3442 17978 3592 17980
rect 3442 17932 3452 17978
rect 3498 17932 3592 17978
rect 3442 17928 3592 17932
rect 3324 17908 3592 17928
rect 2433 17667 2467 17713
rect 2513 17667 2547 17713
rect 2433 17550 2547 17667
rect 2685 17817 2793 17829
rect 2685 17661 2716 17817
rect 2768 17661 2793 17817
rect 2187 17170 2243 17216
rect 2289 17170 2295 17216
rect 2187 17133 2295 17170
rect 2433 17216 2547 17253
rect 2433 17170 2467 17216
rect 2513 17170 2547 17216
rect 1676 17024 2065 17105
rect 2433 17024 2547 17170
rect 2685 17216 2793 17661
rect 2936 17713 3282 17829
rect 2936 17667 2970 17713
rect 3016 17667 3202 17713
rect 3248 17667 3282 17713
rect 2936 17550 3282 17667
rect 3425 17817 3533 17829
rect 3425 17661 3450 17817
rect 3502 17661 3533 17817
rect 3076 17253 3144 17256
rect 2685 17170 2691 17216
rect 2737 17170 2793 17216
rect 2685 17133 2793 17170
rect 2915 17245 3303 17253
rect 2915 17216 3087 17245
rect 2961 17170 3087 17216
rect 2915 17105 3087 17170
rect 3133 17216 3303 17245
rect 3133 17170 3257 17216
rect 3133 17105 3303 17170
rect 3425 17216 3533 17661
rect 3671 17713 3785 18085
rect 3864 17980 4132 18005
rect 3864 17978 4014 17980
rect 3864 17932 3958 17978
rect 4004 17932 4014 17978
rect 3864 17928 4014 17932
rect 4066 17928 4132 17980
rect 3864 17908 4132 17928
rect 4277 17829 4418 18085
rect 4563 17980 4831 18005
rect 4563 17928 4629 17980
rect 4681 17978 4831 17980
rect 4681 17932 4691 17978
rect 4737 17932 4831 17978
rect 4681 17928 4831 17932
rect 4563 17908 4831 17928
rect 3671 17667 3705 17713
rect 3751 17667 3785 17713
rect 3671 17550 3785 17667
rect 3923 17817 4031 17829
rect 3923 17661 3954 17817
rect 4006 17661 4031 17817
rect 3425 17170 3481 17216
rect 3527 17170 3533 17216
rect 3425 17133 3533 17170
rect 3671 17216 3785 17253
rect 3671 17170 3705 17216
rect 3751 17170 3785 17216
rect 2915 17024 3303 17105
rect 3671 17024 3785 17170
rect 3923 17216 4031 17661
rect 4174 17713 4521 17829
rect 4174 17667 4208 17713
rect 4254 17667 4441 17713
rect 4487 17667 4521 17713
rect 4174 17550 4521 17667
rect 4664 17817 4772 17829
rect 4664 17661 4689 17817
rect 4741 17661 4772 17817
rect 4314 17253 4382 17256
rect 3923 17170 3929 17216
rect 3975 17170 4031 17216
rect 3923 17133 4031 17170
rect 4153 17245 4542 17253
rect 4153 17216 4325 17245
rect 4199 17170 4325 17216
rect 4153 17105 4325 17170
rect 4371 17216 4542 17245
rect 4371 17170 4496 17216
rect 4371 17105 4542 17170
rect 4664 17216 4772 17661
rect 4909 17713 5025 18085
rect 5103 17981 5372 18005
rect 5103 17978 5254 17981
rect 5103 17932 5197 17978
rect 5243 17932 5254 17978
rect 5103 17929 5254 17932
rect 5306 17929 5372 17981
rect 5103 17908 5372 17929
rect 5515 17829 5587 18085
rect 4909 17667 4944 17713
rect 4990 17667 5025 17713
rect 4909 17550 5025 17667
rect 5162 17817 5291 17829
rect 5162 17661 5174 17817
rect 5226 17713 5291 17817
rect 5243 17667 5291 17713
rect 5226 17661 5291 17667
rect 5162 17550 5291 17661
rect 5412 17713 5587 17829
rect 5412 17667 5447 17713
rect 5493 17667 5587 17713
rect 5412 17550 5587 17667
rect 5184 17253 5256 17550
rect 5553 17253 5621 17256
rect 4664 17170 4720 17216
rect 4766 17170 4772 17216
rect 4664 17133 4772 17170
rect 4909 17216 5025 17253
rect 4909 17170 4944 17216
rect 4990 17170 5025 17216
rect 4153 17024 4542 17105
rect 4909 17024 5025 17170
rect 5159 17216 5256 17253
rect 5159 17170 5168 17216
rect 5214 17170 5256 17216
rect 5159 17133 5256 17170
rect 5392 17245 5621 17253
rect 5392 17216 5564 17245
rect 5438 17170 5564 17216
rect 5392 17105 5564 17170
rect 5610 17105 5621 17245
rect 5392 17094 5621 17105
rect 5392 17024 5587 17094
rect 510 16933 5587 17024
rect 510 16881 915 16933
rect 967 16881 1535 16933
rect 1587 16881 2154 16933
rect 2206 16881 2774 16933
rect 2826 16881 3392 16933
rect 3444 16881 4012 16933
rect 4064 16881 4631 16933
rect 4683 16881 5251 16933
rect 5303 16881 5587 16933
rect 510 16849 5587 16881
rect 510 16803 754 16849
rect 800 16803 912 16849
rect 958 16803 1070 16849
rect 1116 16803 1228 16849
rect 1274 16803 1386 16849
rect 1432 16803 1544 16849
rect 1590 16803 1702 16849
rect 1748 16803 1993 16849
rect 2039 16803 2151 16849
rect 2197 16803 2309 16849
rect 2355 16803 2467 16849
rect 2513 16803 2625 16849
rect 2671 16803 2783 16849
rect 2829 16803 2941 16849
rect 2987 16803 3231 16849
rect 3277 16803 3389 16849
rect 3435 16803 3547 16849
rect 3593 16803 3705 16849
rect 3751 16803 3863 16849
rect 3909 16803 4021 16849
rect 4067 16803 4179 16849
rect 4225 16803 4470 16849
rect 4516 16803 4628 16849
rect 4674 16803 4786 16849
rect 4832 16803 4944 16849
rect 4990 16803 5102 16849
rect 5148 16803 5260 16849
rect 5306 16803 5418 16849
rect 5464 16803 5587 16849
rect 510 16752 5587 16803
rect 678 16616 2390 16641
rect 678 16564 728 16616
rect 780 16564 914 16616
rect 966 16564 1745 16616
rect 1797 16564 1931 16616
rect 1983 16564 2390 16616
rect 678 16544 2390 16564
rect 678 16428 2390 16432
rect 678 16408 2624 16428
rect 678 16356 1108 16408
rect 1160 16356 1294 16408
rect 1346 16356 2346 16408
rect 2398 16356 2532 16408
rect 2584 16356 2624 16408
rect 678 16336 2624 16356
rect 4824 16408 5132 16428
rect 4824 16356 4854 16408
rect 4906 16356 5040 16408
rect 5092 16356 5132 16408
rect 4824 16336 5132 16356
rect 678 16335 2390 16336
rect 929 16223 1058 16224
rect 368 16220 2390 16223
rect 368 16183 3373 16220
rect 368 16131 967 16183
rect 1019 16180 3373 16183
rect 1019 16131 1806 16180
rect 368 16128 1806 16131
rect 1858 16128 2017 16180
rect 2069 16128 2227 16180
rect 2279 16128 2438 16180
rect 2490 16128 2650 16180
rect 2702 16128 2861 16180
rect 2913 16128 3071 16180
rect 3123 16128 3282 16180
rect 3334 16128 3373 16180
rect 368 16087 3373 16128
rect 3720 16180 4482 16220
rect 3720 16128 3758 16180
rect 3810 16128 3969 16180
rect 4021 16128 4181 16180
rect 4233 16128 4392 16180
rect 4444 16128 4482 16180
rect 3720 16087 4482 16128
rect 368 16086 2390 16087
rect 487 15946 1903 15969
rect 487 15894 536 15946
rect 588 15894 1903 15946
rect 487 15873 1903 15894
rect 2258 15929 2350 15970
rect 2258 15877 2278 15929
rect 2330 15877 2350 15929
rect 913 15774 1413 15775
rect 300 15758 346 15771
rect 277 15605 300 15635
rect 524 15758 570 15771
rect 346 15605 369 15635
rect 277 15553 297 15605
rect 349 15553 369 15605
rect 277 15419 300 15553
rect 346 15419 369 15553
rect 277 15367 297 15419
rect 349 15367 369 15419
rect 277 15327 300 15367
rect 277 15006 300 15036
rect 346 15327 369 15367
rect 346 15006 369 15036
rect 277 14954 297 15006
rect 349 14954 369 15006
rect 277 14820 300 14954
rect 346 14820 369 14954
rect 277 14768 297 14820
rect 349 14768 369 14820
rect 277 14728 300 14768
rect 277 13549 300 13579
rect 346 14728 369 14768
rect 346 13549 369 13579
rect 277 13497 297 13549
rect 349 13497 369 13549
rect 277 13363 300 13497
rect 346 13363 369 13497
rect 277 13311 297 13363
rect 349 13311 369 13363
rect 277 13271 300 13311
rect 346 13271 369 13311
rect 300 13049 346 13062
rect 489 13062 524 13324
rect 913 15734 1491 15774
rect 913 15700 1419 15734
rect 913 15584 1009 15700
rect 1399 15682 1419 15700
rect 1471 15682 1491 15734
rect 913 15538 948 15584
rect 994 15538 1009 15584
rect 913 15478 1009 15538
rect 1126 15584 1292 15620
rect 1126 15538 1211 15584
rect 1257 15538 1292 15584
rect 1126 15501 1292 15538
rect 1399 15548 1491 15682
rect 2258 15743 2350 15877
rect 2258 15691 2278 15743
rect 2330 15691 2350 15743
rect 2258 15651 2350 15691
rect 790 15361 1048 15398
rect 790 15358 990 15361
rect 790 15306 967 15358
rect 1036 15315 1048 15361
rect 1019 15306 1048 15315
rect 790 15265 1048 15306
rect 1126 15181 1198 15501
rect 1399 15496 1419 15548
rect 1471 15496 1491 15548
rect 1399 15455 1491 15496
rect 1627 15558 1935 15578
rect 1627 15506 1657 15558
rect 1709 15555 1843 15558
rect 1895 15555 1935 15558
rect 1899 15509 1935 15555
rect 1709 15506 1843 15509
rect 1895 15506 1935 15509
rect 1627 15486 1935 15506
rect 2318 15502 2478 15552
rect 1644 15304 1690 15317
rect 1644 15200 1690 15258
rect 818 15065 915 15169
rect 818 15019 853 15065
rect 899 15019 915 15065
rect 818 14902 915 15019
rect 1082 15065 1198 15181
rect 1082 15019 1117 15065
rect 1163 15019 1198 15065
rect 1082 14902 1198 15019
rect 842 14555 915 14902
rect 1126 14709 1198 14902
rect 1074 14695 1198 14709
rect 1074 14649 1108 14695
rect 1154 14649 1198 14695
rect 1074 14635 1198 14649
rect 1315 15170 1431 15181
rect 1315 15140 1449 15170
rect 1315 15088 1377 15140
rect 1429 15088 1449 15140
rect 1315 15065 1449 15088
rect 1315 15019 1350 15065
rect 1396 15019 1449 15065
rect 1315 14954 1449 15019
rect 1315 14902 1377 14954
rect 1429 14902 1449 14954
rect 1315 14862 1449 14902
rect 1644 15096 1690 15154
rect 1868 15304 1914 15486
rect 1868 15200 1914 15258
rect 1868 15096 1914 15154
rect 1644 14992 1690 15050
rect 1644 14888 1690 14946
rect 1315 14555 1387 14862
rect 842 14481 1387 14555
rect 1644 14784 1690 14842
rect 1847 15050 1868 15070
rect 2318 15456 2366 15502
rect 2412 15456 2478 15502
rect 2318 15338 2478 15456
rect 2318 15292 2366 15338
rect 2412 15292 2478 15338
rect 2318 15175 2478 15292
rect 2318 15129 2366 15175
rect 2412 15129 2478 15175
rect 1914 15050 1939 15070
rect 1847 15040 1939 15050
rect 1847 14988 1867 15040
rect 1919 14988 1939 15040
rect 1847 14946 1868 14988
rect 1914 14946 1939 14988
rect 1847 14888 1939 14946
rect 1847 14854 1868 14888
rect 1914 14854 1939 14888
rect 1847 14802 1867 14854
rect 1919 14802 1939 14854
rect 1847 14784 1939 14802
rect 1847 14762 1868 14784
rect 1644 14680 1690 14738
rect 1644 14576 1690 14634
rect 1644 14472 1690 14530
rect 748 14398 794 14411
rect 720 14352 748 14391
rect 972 14398 1018 14411
rect 794 14352 812 14391
rect 720 14351 812 14352
rect 720 14299 740 14351
rect 792 14299 812 14351
rect 720 14291 812 14299
rect 720 14245 748 14291
rect 794 14245 812 14291
rect 720 14184 812 14245
rect 720 14165 748 14184
rect 720 14113 740 14165
rect 794 14138 812 14184
rect 792 14113 812 14138
rect 720 14077 812 14113
rect 720 14072 748 14077
rect 794 14072 812 14077
rect 1196 14398 1242 14411
rect 972 14291 1018 14352
rect 972 14184 1018 14245
rect 972 14077 1018 14138
rect 748 13970 794 14031
rect 748 13863 794 13924
rect 748 13756 794 13817
rect 748 13648 794 13710
rect 748 13540 794 13602
rect 748 13432 794 13494
rect 748 13324 794 13386
rect 1173 14352 1196 14391
rect 1420 14398 1466 14411
rect 1242 14352 1265 14391
rect 1173 14351 1265 14352
rect 1173 14299 1193 14351
rect 1245 14299 1265 14351
rect 1173 14291 1265 14299
rect 1173 14245 1196 14291
rect 1242 14245 1265 14291
rect 1173 14184 1265 14245
rect 1173 14165 1196 14184
rect 1242 14165 1265 14184
rect 1173 14113 1193 14165
rect 1245 14113 1265 14165
rect 1173 14077 1265 14113
rect 1173 14072 1196 14077
rect 972 13970 1018 14031
rect 972 13863 1018 13924
rect 972 13756 1018 13817
rect 972 13648 1018 13710
rect 972 13540 1018 13602
rect 972 13432 1018 13494
rect 972 13324 1018 13386
rect 1242 14072 1265 14077
rect 1420 14291 1466 14352
rect 1420 14184 1466 14245
rect 1420 14077 1466 14138
rect 1196 13970 1242 14031
rect 1196 13863 1242 13924
rect 1196 13756 1242 13817
rect 1196 13648 1242 13710
rect 1196 13540 1242 13602
rect 1196 13432 1242 13494
rect 1196 13324 1242 13386
rect 570 13062 605 13324
rect 489 12889 605 13062
rect 748 13216 794 13278
rect 748 13108 794 13170
rect 748 13049 794 13062
rect 937 13278 972 13324
rect 1018 13278 1053 13324
rect 937 13216 1053 13278
rect 937 13170 972 13216
rect 1018 13170 1053 13216
rect 937 13108 1053 13170
rect 937 13062 972 13108
rect 1018 13062 1053 13108
rect 937 12889 1053 13062
rect 1196 13216 1242 13278
rect 1420 13970 1466 14031
rect 1420 13863 1466 13924
rect 1420 13756 1466 13817
rect 1420 13648 1466 13710
rect 1420 13540 1466 13602
rect 1420 13432 1466 13494
rect 1420 13324 1466 13386
rect 1420 13216 1466 13278
rect 1196 13108 1242 13170
rect 1196 13049 1242 13062
rect 1385 13170 1420 13177
rect 1644 14368 1690 14426
rect 1644 14263 1690 14322
rect 1644 14158 1690 14217
rect 1644 14053 1690 14112
rect 1644 13948 1690 14007
rect 1644 13843 1690 13902
rect 1644 13738 1690 13797
rect 1644 13633 1690 13692
rect 1644 13528 1690 13587
rect 1914 14762 1939 14784
rect 2318 15012 2478 15129
rect 2318 14966 2366 15012
rect 2412 14966 2478 15012
rect 2318 14849 2478 14966
rect 2318 14803 2366 14849
rect 2412 14803 2478 14849
rect 1868 14680 1914 14738
rect 1868 14576 1914 14634
rect 1868 14472 1914 14530
rect 1868 14368 1914 14426
rect 1868 14263 1914 14322
rect 1868 14158 1914 14217
rect 1868 14053 1914 14112
rect 1868 13948 1914 14007
rect 1868 13843 1914 13902
rect 1868 13738 1914 13797
rect 1868 13633 1914 13692
rect 1868 13579 1914 13587
rect 2318 14686 2478 14803
rect 2318 14640 2366 14686
rect 2412 14640 2478 14686
rect 2318 14522 2478 14640
rect 2318 14476 2366 14522
rect 2412 14476 2478 14522
rect 2318 14359 2478 14476
rect 2318 14313 2366 14359
rect 2412 14313 2478 14359
rect 2318 14196 2478 14313
rect 2318 14150 2366 14196
rect 2412 14150 2478 14196
rect 2318 14033 2478 14150
rect 2318 13987 2366 14033
rect 2412 13987 2478 14033
rect 2318 13869 2478 13987
rect 2318 13823 2366 13869
rect 2412 13823 2478 13869
rect 2318 13706 2478 13823
rect 2318 13660 2366 13706
rect 2412 13660 2478 13706
rect 1644 13423 1690 13482
rect 1644 13324 1690 13377
rect 1847 13549 1939 13579
rect 1847 13497 1867 13549
rect 1919 13497 1939 13549
rect 1847 13482 1868 13497
rect 1914 13482 1939 13497
rect 1847 13423 1939 13482
rect 1847 13377 1868 13423
rect 1914 13377 1939 13423
rect 1847 13363 1939 13377
rect 1644 13318 1725 13324
rect 1690 13272 1725 13318
rect 1644 13213 1725 13272
rect 1847 13311 1867 13363
rect 1919 13311 1939 13363
rect 1847 13272 1868 13311
rect 1914 13272 1939 13311
rect 1847 13271 1939 13272
rect 2318 13543 2478 13660
rect 2318 13497 2366 13543
rect 2412 13497 2478 13543
rect 2318 13380 2478 13497
rect 2318 13334 2366 13380
rect 2412 13334 2478 13380
rect 1466 13170 1644 13177
rect 1385 13167 1644 13170
rect 1690 13167 1725 13213
rect 1385 13108 1725 13167
rect 1385 13062 1420 13108
rect 1466 13062 1644 13108
rect 1690 13062 1725 13108
rect 1385 13057 1725 13062
rect 1420 13049 1466 13057
rect 1644 13049 1725 13057
rect 1868 13213 1914 13271
rect 1868 13108 1914 13167
rect 1868 13049 1914 13062
rect 2318 13216 2478 13334
rect 2318 13170 2366 13216
rect 2412 13170 2478 13216
rect 2318 13053 2478 13170
rect 489 12852 1576 12889
rect 489 12806 1516 12852
rect 1562 12806 1576 12852
rect 489 12769 1576 12806
rect 300 12600 346 12613
rect 277 12554 300 12584
rect 489 12600 605 12769
rect 748 12600 794 12612
rect 346 12554 369 12584
rect 277 12502 297 12554
rect 349 12502 369 12554
rect 489 12513 524 12600
rect 277 12368 300 12502
rect 346 12368 369 12502
rect 277 12316 297 12368
rect 349 12316 369 12368
rect 277 12276 300 12316
rect 277 11606 300 11636
rect 346 12276 369 12316
rect 346 11606 369 11636
rect 277 11554 297 11606
rect 349 11554 369 11606
rect 277 11420 300 11554
rect 346 11420 369 11554
rect 277 11368 297 11420
rect 349 11368 369 11420
rect 277 11328 300 11368
rect 277 10690 300 10720
rect 346 11328 369 11368
rect 346 10690 369 10720
rect 277 10638 297 10690
rect 349 10638 369 10690
rect 277 10504 300 10638
rect 346 10504 369 10638
rect 277 10452 297 10504
rect 349 10452 369 10504
rect 277 10412 300 10452
rect 346 10412 369 10452
rect 300 9891 346 9904
rect 570 12513 605 12600
rect 723 12599 815 12600
rect 723 12560 748 12599
rect 794 12560 815 12599
rect 723 12508 743 12560
rect 795 12508 815 12560
rect 937 12599 1053 12769
rect 1653 12612 1725 13049
rect 2318 13007 2366 13053
rect 2412 13007 2478 13053
rect 2318 12890 2478 13007
rect 2318 12844 2366 12890
rect 2412 12844 2478 12890
rect 2318 12726 2478 12844
rect 2318 12680 2366 12726
rect 2412 12680 2478 12726
rect 2073 12622 2165 12652
rect 2073 12614 2093 12622
rect 1196 12600 1242 12612
rect 1420 12603 1466 12612
rect 1644 12603 1725 12612
rect 937 12553 972 12599
rect 1018 12553 1053 12599
rect 937 12513 1053 12553
rect 1173 12599 1265 12600
rect 1173 12560 1196 12599
rect 1242 12560 1265 12599
rect 723 12495 815 12508
rect 723 12449 748 12495
rect 794 12449 815 12495
rect 723 12391 815 12449
rect 723 12374 748 12391
rect 794 12374 815 12391
rect 723 12322 743 12374
rect 795 12322 815 12374
rect 723 12287 815 12322
rect 723 12281 748 12287
rect 794 12281 815 12287
rect 972 12495 1018 12513
rect 972 12391 1018 12449
rect 972 12287 1018 12345
rect 748 12183 794 12241
rect 748 12079 794 12137
rect 748 11975 794 12033
rect 748 11871 794 11929
rect 748 11767 794 11825
rect 748 11663 794 11721
rect 748 11558 794 11617
rect 748 11453 794 11512
rect 748 11348 794 11407
rect 748 11243 794 11302
rect 748 11138 794 11197
rect 748 11033 794 11092
rect 748 10928 794 10987
rect 748 10823 794 10882
rect 748 10718 794 10777
rect 748 10613 794 10672
rect 748 10508 794 10567
rect 748 10403 794 10462
rect 748 10344 794 10357
rect 1173 12508 1193 12560
rect 1245 12508 1265 12560
rect 1173 12495 1265 12508
rect 1173 12449 1196 12495
rect 1242 12449 1265 12495
rect 1385 12599 1725 12603
rect 1385 12553 1420 12599
rect 1466 12553 1644 12599
rect 1690 12553 1725 12599
rect 1385 12495 1725 12553
rect 1385 12483 1420 12495
rect 1173 12391 1265 12449
rect 1173 12374 1196 12391
rect 1242 12374 1265 12391
rect 1173 12322 1193 12374
rect 1245 12322 1265 12374
rect 1173 12287 1265 12322
rect 1173 12281 1196 12287
rect 972 12183 1018 12241
rect 972 12079 1018 12137
rect 972 11975 1018 12033
rect 972 11871 1018 11929
rect 972 11767 1018 11825
rect 972 11663 1018 11721
rect 972 11558 1018 11617
rect 972 11453 1018 11512
rect 972 11348 1018 11407
rect 972 11243 1018 11302
rect 972 11138 1018 11197
rect 972 11033 1018 11092
rect 972 10928 1018 10987
rect 972 10823 1018 10882
rect 972 10718 1018 10777
rect 972 10613 1018 10672
rect 972 10508 1018 10567
rect 972 10403 1018 10462
rect 972 10344 1018 10357
rect 1242 12281 1265 12287
rect 1466 12483 1644 12495
rect 1420 12391 1466 12449
rect 1420 12287 1466 12345
rect 1196 12183 1242 12241
rect 1196 12079 1242 12137
rect 1196 11975 1242 12033
rect 1196 11871 1242 11929
rect 1196 11767 1242 11825
rect 1196 11663 1242 11721
rect 1196 11558 1242 11617
rect 1196 11453 1242 11512
rect 1196 11348 1242 11407
rect 1196 11243 1242 11302
rect 1196 11138 1242 11197
rect 1196 11033 1242 11092
rect 1196 10928 1242 10987
rect 1196 10823 1242 10882
rect 1196 10718 1242 10777
rect 1196 10613 1242 10672
rect 1196 10508 1242 10567
rect 1196 10403 1242 10462
rect 1196 10344 1242 10357
rect 1420 12183 1466 12241
rect 1420 12079 1466 12137
rect 1420 11975 1466 12033
rect 1420 11871 1466 11929
rect 1420 11767 1466 11825
rect 1420 11663 1466 11721
rect 1420 11558 1466 11617
rect 1420 11453 1466 11512
rect 1420 11348 1466 11407
rect 1420 11243 1466 11302
rect 1420 11138 1466 11197
rect 1420 11033 1466 11092
rect 1420 10928 1466 10987
rect 1420 10823 1466 10882
rect 1420 10718 1466 10777
rect 1420 10613 1466 10672
rect 1420 10508 1466 10567
rect 1420 10403 1466 10462
rect 1420 10344 1466 10357
rect 1690 12483 1725 12495
rect 1833 12599 2093 12614
rect 1833 12554 1868 12599
rect 1914 12570 2093 12599
rect 2145 12614 2165 12622
rect 2318 12614 2478 12680
rect 2145 12570 2478 12614
rect 1914 12564 2478 12570
rect 1833 12502 1854 12554
rect 1914 12553 2208 12564
rect 1906 12518 2208 12553
rect 2254 12563 2478 12564
rect 2254 12518 2366 12563
rect 1906 12517 2366 12518
rect 2412 12517 2478 12563
rect 1906 12502 2478 12517
rect 1833 12495 2478 12502
rect 1644 12391 1690 12449
rect 1644 12287 1690 12345
rect 1644 12183 1690 12241
rect 1644 12079 1690 12137
rect 1644 11975 1690 12033
rect 1644 11871 1690 11929
rect 1644 11767 1690 11825
rect 1644 11663 1690 11721
rect 1644 11558 1690 11617
rect 1644 11453 1690 11512
rect 1644 11348 1690 11407
rect 1644 11243 1690 11302
rect 1644 11138 1690 11197
rect 1644 11033 1690 11092
rect 1644 10928 1690 10987
rect 1644 10823 1690 10882
rect 1644 10718 1690 10777
rect 1644 10613 1690 10672
rect 1644 10508 1690 10567
rect 1644 10403 1690 10462
rect 1833 12449 1868 12495
rect 1914 12449 2478 12495
rect 1833 12436 2478 12449
rect 1833 12391 2093 12436
rect 1833 12368 1868 12391
rect 1914 12384 2093 12391
rect 2145 12400 2478 12436
rect 2145 12384 2208 12400
rect 1833 12316 1854 12368
rect 1914 12354 2208 12384
rect 2254 12354 2366 12400
rect 2412 12354 2478 12400
rect 1914 12345 2478 12354
rect 1906 12316 2478 12345
rect 1833 12287 2478 12316
rect 1833 12241 1868 12287
rect 1914 12241 2478 12287
rect 1833 12237 2478 12241
rect 1833 12191 2208 12237
rect 2254 12191 2366 12237
rect 2412 12191 2478 12237
rect 1833 12183 2478 12191
rect 1833 12137 1868 12183
rect 1914 12137 2478 12183
rect 1833 12079 2478 12137
rect 1833 12033 1868 12079
rect 1914 12074 2478 12079
rect 1914 12033 2208 12074
rect 1833 12028 2208 12033
rect 2254 12073 2478 12074
rect 2254 12028 2366 12073
rect 1833 12027 2366 12028
rect 2412 12027 2478 12073
rect 1833 11975 2478 12027
rect 1833 11929 1868 11975
rect 1914 11929 2478 11975
rect 1833 11911 2478 11929
rect 1833 11871 2208 11911
rect 1833 11825 1868 11871
rect 1914 11865 2208 11871
rect 2254 11910 2478 11911
rect 2254 11865 2366 11910
rect 1914 11864 2366 11865
rect 2412 11864 2478 11910
rect 1914 11847 2478 11864
rect 1914 11825 2093 11847
rect 1833 11795 2093 11825
rect 2145 11795 2478 11847
rect 1833 11767 2478 11795
rect 1833 11721 1868 11767
rect 1914 11747 2478 11767
rect 1914 11721 2208 11747
rect 1833 11701 2208 11721
rect 2254 11701 2366 11747
rect 2412 11701 2478 11747
rect 1833 11663 2478 11701
rect 1833 11617 1868 11663
rect 1914 11661 2478 11663
rect 1914 11617 2093 11661
rect 1833 11609 2093 11617
rect 2145 11609 2478 11661
rect 1833 11606 2478 11609
rect 1833 11554 1854 11606
rect 1906 11584 2478 11606
rect 1906 11558 2208 11584
rect 1833 11512 1868 11554
rect 1914 11538 2208 11558
rect 2254 11538 2366 11584
rect 2412 11538 2478 11584
rect 1914 11512 2478 11538
rect 1833 11453 2478 11512
rect 1833 11420 1868 11453
rect 1914 11421 2478 11453
rect 1833 11368 1854 11420
rect 1914 11407 2208 11421
rect 1906 11375 2208 11407
rect 2254 11420 2478 11421
rect 2254 11375 2366 11420
rect 1906 11374 2366 11375
rect 2412 11374 2478 11420
rect 1906 11368 2478 11374
rect 1833 11348 2478 11368
rect 1833 11302 1868 11348
rect 1914 11302 2478 11348
rect 1833 11257 2478 11302
rect 1833 11243 2208 11257
rect 1833 11197 1868 11243
rect 1914 11211 2208 11243
rect 2254 11211 2366 11257
rect 2412 11211 2478 11257
rect 1914 11197 2478 11211
rect 1833 11138 2478 11197
rect 1833 11092 1868 11138
rect 1914 11094 2478 11138
rect 1914 11092 2208 11094
rect 1833 11048 2208 11092
rect 2254 11048 2366 11094
rect 2412 11048 2478 11094
rect 1833 11033 2478 11048
rect 1833 10987 1868 11033
rect 1914 10987 2478 11033
rect 1833 10931 2478 10987
rect 1833 10928 2093 10931
rect 1833 10882 1868 10928
rect 1914 10882 2093 10928
rect 1833 10879 2093 10882
rect 2145 10885 2208 10931
rect 2254 10885 2366 10931
rect 2412 10885 2478 10931
rect 2145 10879 2478 10885
rect 1833 10823 2478 10879
rect 1833 10777 1868 10823
rect 1914 10777 2478 10823
rect 1833 10768 2478 10777
rect 1833 10745 2208 10768
rect 1833 10718 2093 10745
rect 1833 10690 1868 10718
rect 1914 10693 2093 10718
rect 2145 10722 2208 10745
rect 2254 10722 2366 10768
rect 2412 10722 2478 10768
rect 2145 10693 2478 10722
rect 1833 10638 1854 10690
rect 1914 10672 2478 10693
rect 1906 10638 2478 10672
rect 1833 10613 2478 10638
rect 1833 10567 1868 10613
rect 1914 10604 2478 10613
rect 1914 10567 2208 10604
rect 1833 10558 2208 10567
rect 2254 10558 2366 10604
rect 2412 10558 2478 10604
rect 1833 10508 2478 10558
rect 1833 10504 1868 10508
rect 1833 10452 1854 10504
rect 1914 10462 2478 10508
rect 1906 10452 2478 10462
rect 1833 10403 2478 10452
rect 1833 10402 1868 10403
rect 1644 10344 1690 10357
rect 1914 10402 2478 10403
rect 1868 10344 1914 10357
rect 941 10258 1229 10272
rect 941 10212 976 10258
rect 1022 10248 1229 10258
rect 941 10196 978 10212
rect 1030 10196 1229 10248
rect 941 10176 1229 10196
rect 5344 10239 5438 11046
rect 5344 10187 5365 10239
rect 5417 10187 5438 10239
rect 524 9891 570 9904
rect 682 10045 2527 10096
rect 5344 10069 5438 10187
rect 682 9999 1741 10045
rect 1787 9999 2527 10045
rect 682 9977 2527 9999
rect 5345 10053 5437 10069
rect 5345 10001 5365 10053
rect 5417 10001 5437 10053
rect 682 9976 2481 9977
rect 682 9790 798 9976
rect 1629 9891 1675 9904
rect 377 9773 798 9790
rect 377 9727 412 9773
rect 458 9727 798 9773
rect 377 9670 798 9727
rect 898 9838 990 9868
rect 898 9791 918 9838
rect 898 9745 911 9791
rect 970 9786 990 9838
rect 1616 9845 1629 9868
rect 1853 9891 1899 9904
rect 1675 9845 1708 9868
rect 1616 9838 1708 9845
rect 957 9745 990 9786
rect 898 9671 990 9745
rect 898 9625 911 9671
rect 957 9652 990 9671
rect 898 9600 918 9625
rect 970 9600 990 9652
rect 1135 9796 1181 9804
rect 1135 9791 1220 9796
rect 1181 9745 1220 9791
rect 1135 9671 1220 9745
rect 1181 9625 1220 9671
rect 1135 9612 1220 9625
rect 252 9559 394 9570
rect 898 9560 990 9600
rect 252 9519 598 9559
rect 252 9518 300 9519
rect 346 9518 598 9519
rect 252 9466 296 9518
rect 348 9466 508 9518
rect 560 9466 598 9518
rect 252 9425 598 9466
rect 252 9422 394 9425
rect 1148 9413 1220 9612
rect 1616 9786 1636 9838
rect 1688 9786 1708 9838
rect 1616 9771 1708 9786
rect 1616 9725 1629 9771
rect 1675 9725 1708 9771
rect 1853 9771 1899 9845
rect 1616 9652 1708 9725
rect 1616 9600 1636 9652
rect 1688 9600 1708 9652
rect 1616 9560 1708 9600
rect 1817 9725 1853 9749
rect 2481 9849 2527 9931
rect 1899 9725 1933 9749
rect 1629 9420 1675 9433
rect 1018 9339 1503 9413
rect 801 9227 847 9240
rect 801 9117 847 9181
rect 1018 9227 1090 9339
rect 1018 9181 1025 9227
rect 1071 9181 1090 9227
rect 573 9097 881 9117
rect 573 9045 603 9097
rect 655 9045 789 9097
rect 841 9071 881 9097
rect 573 9025 801 9045
rect 847 9025 881 9071
rect 1018 9071 1090 9181
rect 1249 9227 1295 9240
rect 1249 9120 1295 9181
rect 1018 9025 1025 9071
rect 1071 9025 1090 9071
rect 801 9012 847 9025
rect 1018 9022 1090 9025
rect 1221 9080 1313 9120
rect 1221 9028 1241 9080
rect 1293 9071 1313 9080
rect 1221 9025 1249 9028
rect 1295 9025 1313 9071
rect 1025 9012 1071 9022
rect 277 9008 369 9011
rect 265 8981 381 9008
rect 265 8929 297 8981
rect 349 8929 381 8981
rect 265 8925 300 8929
rect 346 8925 381 8929
rect 265 8807 381 8925
rect 265 8795 300 8807
rect 346 8795 381 8807
rect 265 8743 297 8795
rect 349 8743 381 8795
rect 550 8880 956 8899
rect 550 8863 875 8880
rect 550 8811 647 8863
rect 699 8811 833 8863
rect 921 8834 956 8880
rect 885 8811 956 8834
rect 1221 8894 1313 9025
rect 1221 8842 1241 8894
rect 1293 8842 1313 8894
rect 1221 8812 1313 8842
rect 1431 9020 1503 9339
rect 1629 9264 1675 9374
rect 1431 8974 1444 9020
rect 1490 8974 1503 9020
rect 1593 9218 1629 9232
rect 1817 9420 1933 9725
rect 2481 9722 2527 9803
rect 2481 9595 2527 9676
rect 1817 9374 1853 9420
rect 1899 9374 1933 9420
rect 1817 9264 1933 9374
rect 2077 9420 2123 9433
rect 2077 9307 2123 9374
rect 1675 9218 1709 9232
rect 1593 9080 1709 9218
rect 1593 9028 1630 9080
rect 1682 9028 1709 9080
rect 1593 8988 1709 9028
rect 1817 9218 1853 9264
rect 1899 9218 1933 9264
rect 2043 9266 2135 9307
rect 2043 9232 2063 9266
rect 2115 9264 2135 9266
rect 1609 8987 1703 8988
rect 550 8790 956 8811
rect 265 8725 381 8743
rect 1039 8731 1131 8771
rect 276 8724 370 8725
rect 277 8703 369 8724
rect 1039 8679 1059 8731
rect 1111 8679 1131 8731
rect 1039 8636 1131 8679
rect 801 8623 847 8636
rect 461 8523 553 8563
rect 461 8471 481 8523
rect 533 8471 553 8523
rect 461 8364 553 8471
rect 801 8520 847 8577
rect 1025 8623 1131 8636
rect 1071 8577 1131 8623
rect 1025 8545 1131 8577
rect 801 8503 882 8520
rect 847 8457 882 8503
rect 801 8444 882 8457
rect 1025 8503 1059 8545
rect 1111 8493 1131 8545
rect 1071 8463 1131 8493
rect 1249 8623 1347 8636
rect 1295 8577 1347 8623
rect 1249 8503 1347 8577
rect 1025 8444 1071 8457
rect 1295 8457 1347 8503
rect 1249 8444 1347 8457
rect 461 8337 732 8364
rect 461 8285 481 8337
rect 533 8327 732 8337
rect 533 8285 673 8327
rect 461 8281 673 8285
rect 719 8281 732 8327
rect 461 8244 732 8281
rect 810 8341 882 8444
rect 810 8327 1197 8341
rect 810 8281 1117 8327
rect 1163 8281 1197 8327
rect 810 8267 1197 8281
rect 810 8163 882 8267
rect 1275 8163 1347 8444
rect 1431 8252 1503 8974
rect 1610 8894 1702 8987
rect 1610 8842 1630 8894
rect 1682 8842 1702 8894
rect 1610 8812 1702 8842
rect 1817 8908 1933 9218
rect 2041 9214 2063 9232
rect 2123 9232 2135 9264
rect 2481 9245 2527 9549
rect 2705 9977 2751 9990
rect 2751 9933 2864 9963
rect 5345 9960 5437 10001
rect 2751 9931 2792 9933
rect 2705 9881 2792 9931
rect 2844 9881 2864 9933
rect 2705 9849 2864 9881
rect 2751 9803 2864 9849
rect 2705 9747 2864 9803
rect 2705 9722 2792 9747
rect 2751 9695 2792 9722
rect 2844 9695 2864 9747
rect 2751 9676 2864 9695
rect 2705 9655 2864 9676
rect 2705 9654 2788 9655
rect 2705 9595 2751 9654
rect 2705 9536 2751 9549
rect 2123 9218 2157 9232
rect 2115 9214 2157 9218
rect 2041 9080 2157 9214
rect 2041 9028 2063 9080
rect 2115 9028 2157 9080
rect 2041 8988 2157 9028
rect 2481 9138 2527 9199
rect 2481 9031 2527 9092
rect 2481 8924 2527 8985
rect 1817 8788 2157 8908
rect 1431 8206 1444 8252
rect 1490 8206 1503 8252
rect 1431 8195 1503 8206
rect 1629 8705 1675 8718
rect 1629 8585 1675 8659
rect 801 8150 882 8163
rect 322 8124 390 8135
rect 322 7984 333 8124
rect 379 7984 390 8124
rect 322 7894 390 7984
rect 847 8104 882 8150
rect 1025 8150 1071 8163
rect 801 8051 882 8104
rect 1017 8104 1025 8136
rect 1249 8150 1347 8163
rect 1071 8104 1110 8136
rect 1017 8096 1110 8104
rect 801 8030 847 8051
rect 1017 8044 1037 8096
rect 1089 8044 1110 8096
rect 1017 8030 1110 8044
rect 1017 8003 1025 8030
rect 801 7971 847 7984
rect 1023 7984 1025 8003
rect 1071 8004 1110 8030
rect 1295 8104 1347 8150
rect 1249 8030 1347 8104
rect 1071 8003 1106 8004
rect 1071 7984 1095 8003
rect 1023 7894 1095 7984
rect 1295 7984 1347 8030
rect 1249 7971 1347 7984
rect 322 7820 1095 7894
rect 1275 7894 1347 7971
rect 1629 8129 1675 8539
rect 1629 8009 1675 8083
rect 1629 7894 1675 7963
rect 1275 7820 1675 7894
rect 1853 8705 1899 8718
rect 1853 8585 1899 8659
rect 1853 8129 1899 8539
rect 1853 8009 1899 8083
rect 1853 7824 1899 7963
rect 2041 8705 2157 8788
rect 2041 8659 2077 8705
rect 2123 8659 2157 8705
rect 2041 8585 2157 8659
rect 2041 8539 2077 8585
rect 2123 8539 2157 8585
rect 2041 8129 2157 8539
rect 2041 8083 2077 8129
rect 2123 8083 2157 8129
rect 2041 8009 2157 8083
rect 2041 7963 2077 8009
rect 2123 7963 2157 8009
rect 2041 7950 2157 7963
rect 2481 8817 2527 8878
rect 2481 8710 2527 8771
rect 2481 8603 2527 8664
rect 2481 8495 2527 8557
rect 2481 8387 2527 8449
rect 2481 8279 2527 8341
rect 2481 8171 2527 8233
rect 2481 8063 2527 8125
rect 2481 7955 2527 8017
rect 2481 7896 2527 7909
rect 2705 9245 2751 9258
rect 2705 9138 2751 9199
rect 2705 9040 2751 9092
rect 2705 9031 2864 9040
rect 2751 9010 2864 9031
rect 2751 8985 2792 9010
rect 2705 8958 2792 8985
rect 2844 8958 2864 9010
rect 2705 8924 2864 8958
rect 2751 8878 2864 8924
rect 2705 8824 2864 8878
rect 2705 8817 2792 8824
rect 2751 8772 2792 8817
rect 2844 8772 2864 8824
rect 2751 8771 2864 8772
rect 2705 8732 2864 8771
rect 2705 8710 2751 8732
rect 2705 8603 2751 8664
rect 2705 8495 2751 8557
rect 2705 8387 2751 8449
rect 2705 8279 2751 8341
rect 2705 8171 2751 8233
rect 2705 8063 2751 8125
rect 2705 7955 2751 8017
rect 2705 7896 2751 7909
rect 1853 7813 2650 7824
rect 1853 7767 2593 7813
rect 2639 7767 2650 7813
rect 1853 7750 2650 7767
rect 3416 7513 3620 7821
rect 1485 6634 1577 6675
rect 1485 6582 1505 6634
rect 1557 6582 1577 6634
rect 1485 6448 1577 6582
rect 1485 6396 1505 6448
rect 1557 6396 1577 6448
rect 1485 6356 1577 6396
rect 4639 5591 4715 5603
rect 4639 5435 4651 5591
rect 4703 5435 4715 5591
rect 4639 5423 4715 5435
rect 5125 5591 5201 5603
rect 5125 5435 5137 5591
rect 5189 5435 5201 5591
rect 5125 5423 5201 5435
rect 2257 3604 2349 3644
rect 2257 3552 2277 3604
rect 2329 3552 2349 3604
rect 2257 3418 2349 3552
rect 2257 3366 2277 3418
rect 2329 3366 2349 3418
rect 2257 3325 2349 3366
rect 1813 1020 1929 1178
rect 2397 907 2480 1027
rect 2621 979 2677 1001
rect 2621 907 2698 979
rect 3346 907 3413 1001
rect 2621 370 2741 559
rect 3366 370 3466 559
rect 866 -101 1046 -89
rect 866 -153 878 -101
rect 1034 -153 1046 -101
rect 866 -165 1046 -153
rect 3000 -2266 3076 -2254
rect 3000 -2422 3012 -2266
rect 3064 -2422 3076 -2266
rect 3000 -2434 3076 -2422
<< via1 >>
rect 918 28918 970 28956
rect 1532 28918 1584 28956
rect 2157 28918 2209 28956
rect 2771 28918 2823 28956
rect 3395 28918 3447 28956
rect 4009 28918 4061 28956
rect 4634 28918 4686 28956
rect 5248 28918 5300 28956
rect 918 28904 964 28918
rect 964 28904 970 28918
rect 1532 28904 1538 28918
rect 1538 28904 1584 28918
rect 2157 28904 2203 28918
rect 2203 28904 2209 28918
rect 2771 28904 2777 28918
rect 2777 28904 2823 28918
rect 3395 28904 3441 28918
rect 3441 28904 3447 28918
rect 4009 28904 4015 28918
rect 4015 28904 4061 28918
rect 4634 28904 4680 28918
rect 4680 28904 4686 28918
rect 5248 28904 5254 28918
rect 5254 28904 5300 28918
rect 918 28718 970 28770
rect 1532 28718 1584 28770
rect 2157 28718 2209 28770
rect 2771 28718 2823 28770
rect 3395 28718 3447 28770
rect 4009 28718 4061 28770
rect 4634 28718 4686 28770
rect 5248 28718 5300 28770
rect 914 28353 918 28386
rect 918 28353 964 28386
rect 964 28353 966 28386
rect 914 28230 966 28353
rect 914 27578 918 27611
rect 918 27578 964 27611
rect 964 27578 966 27611
rect 914 27455 966 27578
rect 1536 28353 1538 28386
rect 1538 28353 1584 28386
rect 1584 28353 1588 28386
rect 1536 28230 1588 28353
rect 1536 27578 1538 27611
rect 1538 27578 1584 27611
rect 1584 27578 1588 27611
rect 1536 27455 1588 27578
rect 2153 28353 2157 28386
rect 2157 28353 2203 28386
rect 2203 28353 2205 28386
rect 2153 28230 2205 28353
rect 2153 27578 2157 27611
rect 2157 27578 2203 27611
rect 2203 27578 2205 27611
rect 2153 27455 2205 27578
rect 2775 28353 2777 28386
rect 2777 28353 2823 28386
rect 2823 28353 2827 28386
rect 2775 28230 2827 28353
rect 2775 27578 2777 27611
rect 2777 27578 2823 27611
rect 2823 27578 2827 27611
rect 2775 27455 2827 27578
rect 3391 28353 3395 28386
rect 3395 28353 3441 28386
rect 3441 28353 3443 28386
rect 3391 28230 3443 28353
rect 3391 27578 3395 27611
rect 3395 27578 3441 27611
rect 3441 27578 3443 27611
rect 3391 27455 3443 27578
rect 4013 28353 4015 28386
rect 4015 28353 4061 28386
rect 4061 28353 4065 28386
rect 4013 28230 4065 28353
rect 4013 27578 4015 27611
rect 4015 27578 4061 27611
rect 4061 27578 4065 27611
rect 4013 27455 4065 27578
rect 4630 28353 4634 28386
rect 4634 28353 4680 28386
rect 4680 28353 4682 28386
rect 4630 28230 4682 28353
rect 4630 27578 4634 27611
rect 4634 27578 4680 27611
rect 4680 27578 4682 27611
rect 4630 27455 4682 27578
rect 5226 28353 5265 28386
rect 5265 28353 5278 28386
rect 5226 28334 5278 28353
rect 5226 28172 5265 28200
rect 5265 28172 5278 28200
rect 5226 28148 5278 28172
rect 5216 27578 5219 27611
rect 5219 27578 5265 27611
rect 5265 27578 5268 27611
rect 5216 27455 5268 27578
rect 448 27045 500 27097
rect 699 26235 751 26391
rect 1129 26235 1181 26391
rect 1321 26235 1373 26391
rect 1751 26235 1803 26391
rect 1938 26235 1990 26391
rect 2368 26235 2420 26391
rect 2560 26235 2612 26391
rect 2990 26235 3042 26391
rect 3176 26235 3228 26391
rect 3606 26235 3658 26391
rect 3798 26235 3850 26391
rect 4228 26235 4280 26391
rect 4415 26235 4467 26391
rect 4845 26235 4897 26391
rect 5041 26235 5093 26391
rect 5459 26235 5511 26391
rect 1117 25195 1169 25351
rect 1333 25195 1385 25351
rect 1225 24650 1277 24677
rect 1225 24417 1228 24650
rect 1228 24417 1274 24650
rect 1274 24417 1277 24650
rect 909 23917 961 23919
rect 909 23871 912 23917
rect 912 23871 958 23917
rect 958 23871 961 23917
rect 909 23763 961 23871
rect 1541 23917 1593 23919
rect 1541 23871 1544 23917
rect 1544 23871 1590 23917
rect 1590 23871 1593 23917
rect 1541 23763 1593 23871
rect 2356 25195 2408 25351
rect 2572 25195 2624 25351
rect 2464 24650 2516 24677
rect 2464 24417 2467 24650
rect 2467 24417 2513 24650
rect 2513 24417 2516 24650
rect 2148 23917 2200 23919
rect 2148 23871 2151 23917
rect 2151 23871 2197 23917
rect 2197 23871 2200 23917
rect 2148 23763 2200 23871
rect 1124 22166 1176 22218
rect 1326 22166 1378 22218
rect 2780 23917 2832 23919
rect 2780 23871 2783 23917
rect 2783 23871 2829 23917
rect 2829 23871 2832 23917
rect 2780 23763 2832 23871
rect 3594 25195 3646 25351
rect 3810 25195 3862 25351
rect 3702 24650 3754 24677
rect 3702 24417 3705 24650
rect 3705 24417 3751 24650
rect 3751 24417 3754 24650
rect 3386 23917 3438 23919
rect 3386 23871 3389 23917
rect 3389 23871 3435 23917
rect 3435 23871 3438 23917
rect 3386 23763 3438 23871
rect 2363 22166 2415 22218
rect 2565 22166 2617 22218
rect 4018 23917 4070 23919
rect 4018 23871 4021 23917
rect 4021 23871 4067 23917
rect 4067 23871 4070 23917
rect 4018 23763 4070 23871
rect 4833 25195 4885 25351
rect 5053 25195 5105 25351
rect 4941 24650 4993 24677
rect 4941 24417 4944 24650
rect 4944 24417 4990 24650
rect 4990 24417 4993 24650
rect 4625 23917 4677 23919
rect 4625 23871 4628 23917
rect 4628 23871 4674 23917
rect 4674 23871 4677 23917
rect 4625 23763 4677 23871
rect 3601 22166 3653 22218
rect 3803 22166 3855 22218
rect 5257 23917 5309 23919
rect 5257 23871 5260 23917
rect 5260 23871 5306 23917
rect 5306 23871 5309 23917
rect 5257 23763 5309 23871
rect 4840 22166 4892 22218
rect 5042 22166 5094 22218
rect 831 21968 883 22020
rect 1619 21968 1671 22020
rect 2070 21968 2122 22020
rect 2858 21968 2910 22020
rect 3308 21968 3360 22020
rect 4096 21968 4148 22020
rect 4547 21968 4599 22020
rect 5327 21975 5379 22027
rect 699 21760 751 21812
rect 913 20176 918 20212
rect 918 20176 964 20212
rect 964 20176 965 20212
rect 913 20160 965 20176
rect 915 19945 967 19948
rect 915 19899 918 19945
rect 918 19899 964 19945
rect 964 19899 967 19945
rect 915 19896 967 19899
rect 1751 21760 1803 21812
rect 1938 21760 1990 21812
rect 1537 20176 1538 20212
rect 1538 20176 1584 20212
rect 1584 20176 1589 20212
rect 1537 20160 1589 20176
rect 1535 19945 1587 19948
rect 1535 19899 1538 19945
rect 1538 19899 1584 19945
rect 1584 19899 1587 19945
rect 1535 19896 1587 19899
rect 734 18328 786 18380
rect 2152 20176 2157 20212
rect 2157 20176 2203 20212
rect 2203 20176 2204 20212
rect 2152 20160 2204 20176
rect 2154 19945 2206 19948
rect 2154 19899 2157 19945
rect 2157 19899 2203 19945
rect 2203 19899 2206 19945
rect 2154 19896 2206 19899
rect 2990 21760 3042 21812
rect 3176 21760 3228 21812
rect 2776 20176 2777 20212
rect 2777 20176 2823 20212
rect 2823 20176 2828 20212
rect 2776 20160 2828 20176
rect 2774 19945 2826 19948
rect 2774 19899 2777 19945
rect 2777 19899 2823 19945
rect 2823 19899 2826 19945
rect 2774 19896 2826 19899
rect 1747 18328 1799 18380
rect 1933 18328 1985 18380
rect 3390 20176 3395 20212
rect 3395 20176 3441 20212
rect 3441 20176 3442 20212
rect 3390 20160 3442 20176
rect 3392 19945 3444 19948
rect 3392 19899 3395 19945
rect 3395 19899 3441 19945
rect 3441 19899 3444 19945
rect 3392 19896 3444 19899
rect 4228 21760 4280 21812
rect 4415 21760 4467 21812
rect 4014 20176 4015 20212
rect 4015 20176 4061 20212
rect 4061 20176 4066 20212
rect 4014 20160 4066 20176
rect 4012 19945 4064 19948
rect 4012 19899 4015 19945
rect 4015 19899 4061 19945
rect 4061 19899 4064 19945
rect 4012 19896 4064 19899
rect 2985 18328 3037 18380
rect 3171 18328 3223 18380
rect 4629 20176 4634 20212
rect 4634 20176 4680 20212
rect 4680 20176 4681 20212
rect 4629 20160 4681 20176
rect 4631 19945 4683 19948
rect 4631 19899 4634 19945
rect 4634 19899 4680 19945
rect 4680 19899 4683 19945
rect 4631 19896 4683 19899
rect 5459 21759 5511 21811
rect 5253 20176 5254 20212
rect 5254 20176 5300 20212
rect 5300 20176 5305 20212
rect 5253 20160 5305 20176
rect 5251 19945 5303 19949
rect 5251 19899 5254 19945
rect 5254 19899 5300 19945
rect 5300 19899 5303 19945
rect 5251 19897 5303 19899
rect 4224 18328 4276 18380
rect 4410 18328 4462 18380
rect 5429 18328 5481 18380
rect 1699 18168 1751 18171
rect 1699 18122 1702 18168
rect 1702 18122 1748 18168
rect 1748 18122 1751 18168
rect 1699 18119 1751 18122
rect 1990 18168 2042 18171
rect 2938 18168 2990 18171
rect 1990 18122 1993 18168
rect 1993 18122 2039 18168
rect 2039 18122 2042 18168
rect 2938 18122 2941 18168
rect 2941 18122 2987 18168
rect 2987 18122 2990 18168
rect 1990 18119 2042 18122
rect 2938 18119 2990 18122
rect 3229 18168 3281 18171
rect 4176 18168 4228 18171
rect 3229 18122 3231 18168
rect 3231 18122 3277 18168
rect 3277 18122 3281 18168
rect 4176 18122 4179 18168
rect 4179 18122 4225 18168
rect 4225 18122 4228 18168
rect 3229 18119 3281 18122
rect 4176 18119 4228 18122
rect 4467 18168 4519 18171
rect 4467 18122 4470 18168
rect 4470 18122 4516 18168
rect 4516 18122 4519 18168
rect 4467 18119 4519 18122
rect 913 17928 965 17980
rect 973 17713 1025 17817
rect 973 17667 975 17713
rect 975 17667 1021 17713
rect 1021 17667 1025 17713
rect 973 17661 1025 17667
rect 1537 17928 1589 17980
rect 2152 17928 2204 17980
rect 1477 17713 1529 17817
rect 1477 17667 1481 17713
rect 1481 17667 1527 17713
rect 1527 17667 1529 17713
rect 1477 17661 1529 17667
rect 2212 17713 2264 17817
rect 2212 17667 2214 17713
rect 2214 17667 2260 17713
rect 2260 17667 2264 17713
rect 2212 17661 2264 17667
rect 2776 17928 2828 17980
rect 3390 17928 3442 17980
rect 2716 17713 2768 17817
rect 2716 17667 2720 17713
rect 2720 17667 2766 17713
rect 2766 17667 2768 17713
rect 2716 17661 2768 17667
rect 3450 17713 3502 17817
rect 3450 17667 3452 17713
rect 3452 17667 3498 17713
rect 3498 17667 3502 17713
rect 3450 17661 3502 17667
rect 4014 17928 4066 17980
rect 4629 17928 4681 17980
rect 3954 17713 4006 17817
rect 3954 17667 3958 17713
rect 3958 17667 4004 17713
rect 4004 17667 4006 17713
rect 3954 17661 4006 17667
rect 4689 17713 4741 17817
rect 4689 17667 4691 17713
rect 4691 17667 4737 17713
rect 4737 17667 4741 17713
rect 4689 17661 4741 17667
rect 5254 17929 5306 17981
rect 5174 17713 5226 17817
rect 5174 17667 5197 17713
rect 5197 17667 5226 17713
rect 5174 17661 5226 17667
rect 915 16881 967 16933
rect 1535 16881 1587 16933
rect 2154 16881 2206 16933
rect 2774 16881 2826 16933
rect 3392 16881 3444 16933
rect 4012 16881 4064 16933
rect 4631 16881 4683 16933
rect 5251 16881 5303 16933
rect 728 16564 780 16616
rect 914 16564 966 16616
rect 1745 16564 1797 16616
rect 1931 16564 1983 16616
rect 1108 16356 1160 16408
rect 1294 16356 1346 16408
rect 2346 16356 2398 16408
rect 2532 16356 2584 16408
rect 4854 16356 4906 16408
rect 5040 16356 5092 16408
rect 967 16131 1019 16183
rect 1806 16128 1858 16180
rect 2017 16128 2069 16180
rect 2227 16128 2279 16180
rect 2438 16128 2490 16180
rect 2650 16128 2702 16180
rect 2861 16128 2913 16180
rect 3071 16128 3123 16180
rect 3282 16128 3334 16180
rect 3758 16128 3810 16180
rect 3969 16128 4021 16180
rect 4181 16128 4233 16180
rect 4392 16128 4444 16180
rect 536 15894 588 15946
rect 2278 15877 2330 15929
rect 297 15553 300 15605
rect 300 15553 346 15605
rect 346 15553 349 15605
rect 297 15367 300 15419
rect 300 15367 346 15419
rect 346 15367 349 15419
rect 297 14954 300 15006
rect 300 14954 346 15006
rect 346 14954 349 15006
rect 297 14768 300 14820
rect 300 14768 346 14820
rect 346 14768 349 14820
rect 297 13497 300 13549
rect 300 13497 346 13549
rect 346 13497 349 13549
rect 297 13311 300 13363
rect 300 13311 346 13363
rect 346 13311 349 13363
rect 1419 15682 1471 15734
rect 2278 15691 2330 15743
rect 967 15315 990 15358
rect 990 15315 1019 15358
rect 967 15306 1019 15315
rect 1419 15496 1471 15548
rect 1657 15555 1709 15558
rect 1843 15555 1895 15558
rect 1657 15509 1665 15555
rect 1665 15509 1709 15555
rect 1843 15509 1895 15555
rect 1657 15506 1709 15509
rect 1843 15506 1895 15509
rect 1377 15088 1429 15140
rect 1377 14902 1429 14954
rect 1867 14992 1919 15040
rect 1867 14988 1868 14992
rect 1868 14988 1914 14992
rect 1914 14988 1919 14992
rect 1867 14842 1868 14854
rect 1868 14842 1914 14854
rect 1914 14842 1919 14854
rect 1867 14802 1919 14842
rect 740 14299 792 14351
rect 740 14138 748 14165
rect 748 14138 792 14165
rect 740 14113 792 14138
rect 1193 14299 1245 14351
rect 1193 14138 1196 14165
rect 1196 14138 1242 14165
rect 1242 14138 1245 14165
rect 1193 14113 1245 14138
rect 1867 13528 1919 13549
rect 1867 13497 1868 13528
rect 1868 13497 1914 13528
rect 1914 13497 1919 13528
rect 1867 13318 1919 13363
rect 1867 13311 1868 13318
rect 1868 13311 1914 13318
rect 1914 13311 1919 13318
rect 297 12502 300 12554
rect 300 12502 346 12554
rect 346 12502 349 12554
rect 297 12316 300 12368
rect 300 12316 346 12368
rect 346 12316 349 12368
rect 297 11554 300 11606
rect 300 11554 346 11606
rect 346 11554 349 11606
rect 297 11368 300 11420
rect 300 11368 346 11420
rect 346 11368 349 11420
rect 297 10638 300 10690
rect 300 10638 346 10690
rect 346 10638 349 10690
rect 297 10452 300 10504
rect 300 10452 346 10504
rect 346 10452 349 10504
rect 743 12553 748 12560
rect 748 12553 794 12560
rect 794 12553 795 12560
rect 743 12508 795 12553
rect 743 12345 748 12374
rect 748 12345 794 12374
rect 794 12345 795 12374
rect 743 12322 795 12345
rect 1193 12553 1196 12560
rect 1196 12553 1242 12560
rect 1242 12553 1245 12560
rect 1193 12508 1245 12553
rect 1193 12345 1196 12374
rect 1196 12345 1242 12374
rect 1242 12345 1245 12374
rect 1193 12322 1245 12345
rect 2093 12570 2145 12622
rect 1854 12553 1868 12554
rect 1868 12553 1906 12554
rect 1854 12502 1906 12553
rect 2093 12384 2145 12436
rect 1854 12345 1868 12368
rect 1868 12345 1906 12368
rect 1854 12316 1906 12345
rect 2093 11795 2145 11847
rect 2093 11609 2145 11661
rect 1854 11558 1906 11606
rect 1854 11554 1868 11558
rect 1868 11554 1906 11558
rect 1854 11407 1868 11420
rect 1868 11407 1906 11420
rect 1854 11368 1906 11407
rect 2093 10879 2145 10931
rect 2093 10693 2145 10745
rect 1854 10672 1868 10690
rect 1868 10672 1906 10690
rect 1854 10638 1906 10672
rect 1854 10462 1868 10504
rect 1868 10462 1906 10504
rect 1854 10452 1906 10462
rect 978 10212 1022 10248
rect 1022 10212 1030 10248
rect 978 10196 1030 10212
rect 5365 10187 5417 10239
rect 5365 10001 5417 10053
rect 918 9791 970 9838
rect 918 9786 957 9791
rect 957 9786 970 9791
rect 918 9625 957 9652
rect 957 9625 970 9652
rect 918 9600 970 9625
rect 296 9473 300 9518
rect 300 9473 346 9518
rect 346 9473 348 9518
rect 296 9466 348 9473
rect 508 9466 560 9518
rect 1636 9786 1688 9838
rect 1636 9600 1688 9652
rect 603 9045 655 9097
rect 789 9071 841 9097
rect 789 9045 801 9071
rect 801 9045 841 9071
rect 1241 9071 1293 9080
rect 1241 9028 1249 9071
rect 1249 9028 1293 9071
rect 297 8971 349 8981
rect 297 8929 300 8971
rect 300 8929 346 8971
rect 346 8929 349 8971
rect 297 8761 300 8795
rect 300 8761 346 8795
rect 346 8761 349 8795
rect 297 8743 349 8761
rect 647 8811 699 8863
rect 833 8834 875 8863
rect 875 8834 885 8863
rect 833 8811 885 8834
rect 1241 8842 1293 8894
rect 1630 9028 1682 9080
rect 2063 9264 2115 9266
rect 1059 8679 1111 8731
rect 481 8471 533 8523
rect 1059 8503 1111 8545
rect 1059 8493 1071 8503
rect 1071 8493 1111 8503
rect 481 8285 533 8337
rect 1630 8842 1682 8894
rect 2063 9218 2077 9264
rect 2077 9218 2115 9264
rect 2792 9881 2844 9933
rect 2792 9695 2844 9747
rect 2063 9214 2115 9218
rect 2063 9028 2115 9080
rect 1037 8044 1089 8096
rect 2792 8958 2844 9010
rect 2792 8772 2844 8824
rect 1505 6582 1557 6634
rect 1505 6396 1557 6448
rect 4651 5435 4703 5591
rect 5137 5435 5189 5591
rect 2277 3552 2329 3604
rect 2277 3366 2329 3418
rect 878 -153 1034 -101
rect 3012 -2422 3064 -2266
<< metal2 >>
rect 697 27561 753 28978
rect 877 28958 1005 28980
rect 877 28902 916 28958
rect 972 28902 1005 28958
rect 877 28772 1005 28902
rect 877 28716 916 28772
rect 972 28716 1005 28772
rect 877 28697 1005 28716
rect 902 28386 978 28398
rect 902 28230 914 28386
rect 966 28337 978 28386
rect 1127 28337 1183 28978
rect 966 28281 1183 28337
rect 966 28230 978 28281
rect 902 28218 978 28230
rect 902 27611 978 27623
rect 902 27561 914 27611
rect 697 27505 914 27561
rect 271 27118 478 27121
rect 271 27097 540 27118
rect 271 27045 448 27097
rect 500 27045 540 27097
rect 271 27025 540 27045
rect 271 27024 478 27025
rect 80 22626 174 26890
rect 80 22570 99 22626
rect 155 22570 174 22626
rect 80 22440 174 22570
rect 80 22384 99 22440
rect 155 22384 174 22440
rect 80 16131 174 22384
rect 271 15970 366 27024
rect 473 22626 568 26890
rect 697 26403 753 27505
rect 902 27455 914 27505
rect 966 27455 978 27611
rect 902 27443 978 27455
rect 1127 26403 1183 28281
rect 1319 28337 1375 28978
rect 1497 28958 1625 28980
rect 1497 28902 1530 28958
rect 1586 28902 1625 28958
rect 1497 28772 1625 28902
rect 1497 28716 1530 28772
rect 1586 28716 1625 28772
rect 1497 28697 1625 28716
rect 1524 28386 1600 28398
rect 1524 28337 1536 28386
rect 1319 28281 1536 28337
rect 1319 26403 1375 28281
rect 1524 28230 1536 28281
rect 1588 28230 1600 28386
rect 1524 28218 1600 28230
rect 1524 27611 1600 27623
rect 1524 27455 1536 27611
rect 1588 27561 1600 27611
rect 1749 27561 1805 28978
rect 1588 27505 1805 27561
rect 1588 27455 1600 27505
rect 1524 27443 1600 27455
rect 1749 26403 1805 27505
rect 1936 27561 1992 28978
rect 2116 28958 2244 28980
rect 2116 28902 2155 28958
rect 2211 28902 2244 28958
rect 2116 28772 2244 28902
rect 2116 28716 2155 28772
rect 2211 28716 2244 28772
rect 2116 28697 2244 28716
rect 2141 28386 2217 28398
rect 2141 28230 2153 28386
rect 2205 28337 2217 28386
rect 2366 28337 2422 28978
rect 2205 28281 2422 28337
rect 2205 28230 2217 28281
rect 2141 28218 2217 28230
rect 2141 27611 2217 27623
rect 2141 27561 2153 27611
rect 1936 27505 2153 27561
rect 1936 26403 1992 27505
rect 2141 27455 2153 27505
rect 2205 27455 2217 27611
rect 2141 27443 2217 27455
rect 2366 26403 2422 28281
rect 2558 28337 2614 28978
rect 2736 28958 2864 28980
rect 2736 28902 2769 28958
rect 2825 28902 2864 28958
rect 2736 28772 2864 28902
rect 2736 28716 2769 28772
rect 2825 28716 2864 28772
rect 2736 28697 2864 28716
rect 2763 28386 2839 28398
rect 2763 28337 2775 28386
rect 2558 28281 2775 28337
rect 2558 26403 2614 28281
rect 2763 28230 2775 28281
rect 2827 28230 2839 28386
rect 2763 28218 2839 28230
rect 2763 27611 2839 27623
rect 2763 27455 2775 27611
rect 2827 27561 2839 27611
rect 2988 27561 3044 28978
rect 2827 27505 3044 27561
rect 2827 27455 2839 27505
rect 2763 27443 2839 27455
rect 2988 26403 3044 27505
rect 3174 27561 3230 28978
rect 3354 28958 3482 28980
rect 3354 28902 3393 28958
rect 3449 28902 3482 28958
rect 3354 28772 3482 28902
rect 3354 28716 3393 28772
rect 3449 28716 3482 28772
rect 3354 28697 3482 28716
rect 3379 28386 3455 28398
rect 3379 28230 3391 28386
rect 3443 28337 3455 28386
rect 3604 28337 3660 28978
rect 3443 28281 3660 28337
rect 3443 28230 3455 28281
rect 3379 28218 3455 28230
rect 3379 27611 3455 27623
rect 3379 27561 3391 27611
rect 3174 27505 3391 27561
rect 3174 26403 3230 27505
rect 3379 27455 3391 27505
rect 3443 27455 3455 27611
rect 3379 27443 3455 27455
rect 3604 26403 3660 28281
rect 3796 28337 3852 28978
rect 3974 28958 4102 28980
rect 3974 28902 4007 28958
rect 4063 28902 4102 28958
rect 3974 28772 4102 28902
rect 3974 28716 4007 28772
rect 4063 28716 4102 28772
rect 3974 28697 4102 28716
rect 4001 28386 4077 28398
rect 4001 28337 4013 28386
rect 3796 28281 4013 28337
rect 3796 26403 3852 28281
rect 4001 28230 4013 28281
rect 4065 28230 4077 28386
rect 4001 28218 4077 28230
rect 4001 27611 4077 27623
rect 4001 27455 4013 27611
rect 4065 27561 4077 27611
rect 4226 27561 4282 28978
rect 4065 27505 4282 27561
rect 4065 27455 4077 27505
rect 4001 27443 4077 27455
rect 4226 26403 4282 27505
rect 4413 27561 4469 28978
rect 4593 28958 4721 28980
rect 4593 28902 4632 28958
rect 4688 28902 4721 28958
rect 4593 28772 4721 28902
rect 4593 28716 4632 28772
rect 4688 28716 4721 28772
rect 4593 28697 4721 28716
rect 4618 28386 4694 28398
rect 4618 28230 4630 28386
rect 4682 28337 4694 28386
rect 4843 28337 4899 28978
rect 4682 28281 4899 28337
rect 4682 28230 4694 28281
rect 4618 28218 4694 28230
rect 4618 27611 4694 27623
rect 4618 27561 4630 27611
rect 4413 27505 4630 27561
rect 4413 26403 4469 27505
rect 4618 27455 4630 27505
rect 4682 27455 4694 27611
rect 4618 27443 4694 27455
rect 4843 26403 4899 28281
rect 5039 28337 5095 29028
rect 5212 28958 5341 28980
rect 5212 28902 5246 28958
rect 5302 28902 5341 28958
rect 5212 28772 5341 28902
rect 5212 28716 5246 28772
rect 5302 28716 5341 28772
rect 5212 28697 5341 28716
rect 5206 28386 5298 28426
rect 5206 28337 5226 28386
rect 5039 28334 5226 28337
rect 5278 28334 5298 28386
rect 5039 28281 5298 28334
rect 5039 26403 5095 28281
rect 5206 28200 5298 28281
rect 5206 28148 5226 28200
rect 5278 28148 5298 28200
rect 5206 28108 5298 28148
rect 5204 27611 5280 27623
rect 5204 27455 5216 27611
rect 5268 27561 5280 27611
rect 5457 27561 5513 29028
rect 5268 27505 5513 27561
rect 5268 27455 5280 27505
rect 5204 27443 5280 27455
rect 5457 26403 5513 27505
rect 687 26391 763 26403
rect 687 26235 699 26391
rect 751 26235 763 26391
rect 687 26223 763 26235
rect 1117 26391 1193 26403
rect 1117 26235 1129 26391
rect 1181 26235 1193 26391
rect 1117 26223 1193 26235
rect 1309 26391 1385 26403
rect 1309 26235 1321 26391
rect 1373 26235 1385 26391
rect 1309 26223 1385 26235
rect 1739 26391 1815 26403
rect 1739 26235 1751 26391
rect 1803 26235 1815 26391
rect 1739 26223 1815 26235
rect 1926 26391 2002 26403
rect 1926 26235 1938 26391
rect 1990 26235 2002 26391
rect 1926 26223 2002 26235
rect 2356 26391 2432 26403
rect 2356 26235 2368 26391
rect 2420 26235 2432 26391
rect 2356 26223 2432 26235
rect 2548 26391 2624 26403
rect 2548 26235 2560 26391
rect 2612 26235 2624 26391
rect 2548 26223 2624 26235
rect 2978 26391 3054 26403
rect 2978 26235 2990 26391
rect 3042 26235 3054 26391
rect 2978 26223 3054 26235
rect 3164 26391 3240 26403
rect 3164 26235 3176 26391
rect 3228 26235 3240 26391
rect 3164 26223 3240 26235
rect 3594 26391 3670 26403
rect 3594 26235 3606 26391
rect 3658 26235 3670 26391
rect 3594 26223 3670 26235
rect 3786 26391 3862 26403
rect 3786 26235 3798 26391
rect 3850 26235 3862 26391
rect 3786 26223 3862 26235
rect 4216 26391 4292 26403
rect 4216 26235 4228 26391
rect 4280 26235 4292 26391
rect 4216 26223 4292 26235
rect 4403 26391 4479 26403
rect 4403 26235 4415 26391
rect 4467 26235 4479 26391
rect 4403 26223 4479 26235
rect 4833 26391 4909 26403
rect 4833 26235 4845 26391
rect 4897 26235 4909 26391
rect 4833 26223 4909 26235
rect 5029 26391 5105 26403
rect 5029 26235 5041 26391
rect 5093 26235 5105 26391
rect 5029 26223 5105 26235
rect 5447 26391 5523 26403
rect 5447 26235 5459 26391
rect 5511 26235 5523 26391
rect 5447 26223 5523 26235
rect 473 22570 492 22626
rect 548 22570 568 22626
rect 473 22440 568 22570
rect 473 22384 492 22440
rect 548 22384 568 22440
rect 473 16131 568 22384
rect 697 21824 753 26223
rect 1127 25363 1183 26223
rect 1105 25351 1183 25363
rect 1105 25195 1117 25351
rect 1169 25195 1183 25351
rect 1105 25183 1183 25195
rect 1319 25363 1375 26223
rect 1319 25351 1397 25363
rect 1319 25195 1333 25351
rect 1385 25195 1397 25351
rect 1319 25183 1397 25195
rect 1213 24679 1289 24689
rect 1213 24415 1223 24679
rect 1279 24415 1289 24679
rect 1213 24405 1289 24415
rect 897 23919 973 23931
rect 897 23763 909 23919
rect 961 23763 973 23919
rect 897 23751 973 23763
rect 1529 23919 1605 23931
rect 1529 23763 1541 23919
rect 1593 23763 1605 23919
rect 1529 23751 1605 23763
rect 907 22150 963 23751
rect 1112 22218 1390 22230
rect 1112 22166 1124 22218
rect 1176 22166 1326 22218
rect 1378 22166 1390 22218
rect 1112 22154 1390 22166
rect 907 22094 1030 22150
rect 819 22020 895 22032
rect 819 22009 831 22020
rect 883 22009 895 22020
rect 819 21849 829 22009
rect 885 21849 895 22009
rect 819 21839 895 21849
rect 687 21812 763 21824
rect 687 21760 699 21812
rect 751 21760 763 21812
rect 687 21748 763 21760
rect 678 20236 770 21270
rect 974 20408 1030 22094
rect 974 20352 1138 20408
rect 678 20212 1001 20236
rect 678 20160 913 20212
rect 965 20160 1001 20212
rect 678 20139 1001 20160
rect 678 18642 770 20139
rect 903 19950 979 19960
rect 1082 19950 1138 20352
rect 903 19948 1138 19950
rect 903 19896 915 19948
rect 967 19896 1138 19948
rect 903 19894 1138 19896
rect 903 19884 979 19894
rect 678 18606 772 18642
rect 678 18604 977 18606
rect 678 18548 697 18604
rect 753 18548 977 18604
rect 678 18509 977 18548
rect 699 18400 826 18401
rect 697 18380 826 18400
rect 697 18328 734 18380
rect 786 18328 826 18380
rect 697 18308 826 18328
rect 697 16641 787 18308
rect 901 17980 977 18509
rect 901 17928 913 17980
rect 965 17928 977 17980
rect 901 17908 977 17928
rect 1082 17829 1138 19894
rect 961 17817 1138 17829
rect 961 17661 973 17817
rect 1025 17661 1138 17817
rect 961 17649 1138 17661
rect 877 16935 1005 17031
rect 877 16879 913 16935
rect 969 16879 1005 16935
rect 877 16802 1005 16879
rect 1223 16754 1279 22154
rect 1539 22150 1595 23751
rect 1472 22094 1595 22150
rect 1472 20408 1528 22094
rect 1607 22020 1683 22032
rect 1607 22009 1619 22020
rect 1671 22009 1683 22020
rect 1607 21849 1617 22009
rect 1673 21849 1683 22009
rect 1607 21839 1683 21849
rect 1749 21824 1805 26223
rect 1936 21824 1992 26223
rect 2366 25363 2422 26223
rect 2344 25351 2422 25363
rect 2344 25195 2356 25351
rect 2408 25195 2422 25351
rect 2344 25183 2422 25195
rect 2558 25363 2614 26223
rect 2558 25351 2636 25363
rect 2558 25195 2572 25351
rect 2624 25195 2636 25351
rect 2558 25183 2636 25195
rect 2452 24679 2528 24689
rect 2452 24415 2462 24679
rect 2518 24415 2528 24679
rect 2452 24405 2528 24415
rect 2136 23919 2212 23931
rect 2136 23763 2148 23919
rect 2200 23763 2212 23919
rect 2136 23751 2212 23763
rect 2768 23919 2844 23931
rect 2768 23763 2780 23919
rect 2832 23763 2844 23919
rect 2768 23751 2844 23763
rect 2146 22150 2202 23751
rect 2351 22218 2629 22230
rect 2351 22166 2363 22218
rect 2415 22166 2565 22218
rect 2617 22166 2629 22218
rect 2351 22154 2629 22166
rect 2146 22094 2269 22150
rect 2058 22020 2134 22032
rect 2058 22009 2070 22020
rect 2122 22009 2134 22020
rect 2058 21849 2068 22009
rect 2124 21849 2134 22009
rect 2058 21839 2134 21849
rect 1739 21812 1815 21824
rect 1739 21760 1751 21812
rect 1803 21760 1815 21812
rect 1739 21748 1815 21760
rect 1926 21812 2002 21824
rect 1926 21760 1938 21812
rect 1990 21760 2002 21812
rect 1926 21748 2002 21760
rect 1364 20352 1528 20408
rect 1364 19950 1420 20352
rect 1732 20236 1824 21270
rect 1501 20212 1824 20236
rect 1501 20160 1537 20212
rect 1589 20160 1824 20212
rect 1501 20139 1824 20160
rect 1523 19950 1599 19960
rect 1364 19948 1599 19950
rect 1364 19896 1535 19948
rect 1587 19896 1599 19948
rect 1364 19894 1599 19896
rect 1364 17829 1420 19894
rect 1523 19884 1599 19894
rect 1732 18957 1824 20139
rect 1917 20236 2009 21270
rect 2213 20408 2269 22094
rect 2213 20352 2377 20408
rect 1917 20212 2240 20236
rect 1917 20160 2152 20212
rect 2204 20160 2240 20212
rect 1917 20139 2240 20160
rect 1917 19284 2009 20139
rect 2142 19950 2218 19960
rect 2321 19950 2377 20352
rect 2142 19948 2377 19950
rect 2142 19896 2154 19948
rect 2206 19896 2377 19948
rect 2142 19894 2377 19896
rect 2142 19884 2218 19894
rect 1916 19246 2010 19284
rect 1916 19190 1935 19246
rect 1991 19190 2010 19246
rect 1916 19151 2010 19190
rect 1732 18919 1826 18957
rect 1732 18863 1751 18919
rect 1807 18863 1826 18919
rect 1732 18824 1826 18863
rect 1732 18606 1824 18824
rect 1525 18509 1824 18606
rect 1917 18606 2009 19151
rect 1917 18509 2216 18606
rect 1525 17980 1601 18509
rect 1717 18380 2025 18400
rect 1717 18328 1747 18380
rect 1799 18328 1933 18380
rect 1985 18328 2025 18380
rect 1717 18308 2025 18328
rect 1525 17928 1537 17980
rect 1589 17928 1601 17980
rect 1525 17908 1601 17928
rect 1687 18173 1763 18195
rect 1687 18013 1697 18173
rect 1753 18013 1763 18173
rect 1687 17913 1763 18013
rect 1364 17817 1541 17829
rect 1364 17661 1477 17817
rect 1529 17661 1541 17817
rect 1364 17649 1541 17661
rect 1497 16935 1625 17031
rect 1497 16879 1533 16935
rect 1589 16879 1625 16935
rect 1497 16802 1625 16879
rect 697 16636 814 16641
rect 697 16616 1006 16636
rect 697 16564 728 16616
rect 780 16564 914 16616
rect 966 16564 1006 16616
rect 697 16544 1006 16564
rect 271 15946 628 15970
rect 271 15894 536 15946
rect 588 15894 628 15946
rect 271 15873 628 15894
rect 277 15607 369 15635
rect 277 15551 295 15607
rect 351 15551 369 15607
rect 277 15421 369 15551
rect 277 15365 295 15421
rect 351 15365 369 15421
rect 277 15327 369 15365
rect 277 15008 369 15036
rect 277 14952 295 15008
rect 351 14952 369 15008
rect 277 14822 369 14952
rect 277 14766 295 14822
rect 351 14766 369 14822
rect 277 14728 369 14766
rect 719 14351 814 16544
rect 1207 16432 1297 16754
rect 1172 16428 1297 16432
rect 1078 16408 1386 16428
rect 1078 16356 1108 16408
rect 1160 16356 1294 16408
rect 1346 16356 1386 16408
rect 1078 16336 1386 16356
rect 1172 16335 1297 16336
rect 928 16185 1058 16224
rect 928 16129 965 16185
rect 1021 16129 1058 16185
rect 928 16090 1058 16129
rect 719 14299 740 14351
rect 792 14299 814 14351
rect 719 14165 814 14299
rect 719 14113 740 14165
rect 792 14113 814 14165
rect 277 13551 369 13579
rect 277 13495 295 13551
rect 351 13495 369 13551
rect 277 13365 369 13495
rect 277 13309 295 13365
rect 351 13309 369 13365
rect 277 13271 369 13309
rect 719 12600 814 14113
rect 946 15358 1040 16090
rect 946 15306 967 15358
rect 1019 15306 1040 15358
rect 277 12556 369 12584
rect 277 12500 295 12556
rect 351 12500 369 12556
rect 277 12370 369 12500
rect 277 12314 295 12370
rect 351 12314 369 12370
rect 277 12276 369 12314
rect 719 12560 815 12600
rect 719 12508 743 12560
rect 795 12508 815 12560
rect 719 12374 815 12508
rect 719 12322 743 12374
rect 795 12322 815 12374
rect 719 12282 815 12322
rect 277 11608 369 11636
rect 277 11552 295 11608
rect 351 11552 369 11608
rect 277 11422 369 11552
rect 277 11366 295 11422
rect 351 11366 369 11422
rect 277 11328 369 11366
rect 277 10692 369 10720
rect 277 10636 295 10692
rect 351 10636 369 10692
rect 277 10506 369 10636
rect 277 10450 295 10506
rect 351 10450 369 10506
rect 277 10412 369 10450
rect 946 10269 1040 15306
rect 1172 14351 1266 16335
rect 1514 15775 1608 16802
rect 1826 16636 1916 18308
rect 1978 18173 2054 18195
rect 1978 18013 1988 18173
rect 2044 18013 2054 18173
rect 1978 17913 2054 18013
rect 2140 17980 2216 18509
rect 2140 17928 2152 17980
rect 2204 17928 2216 17980
rect 2140 17908 2216 17928
rect 2321 17829 2377 19894
rect 2200 17817 2377 17829
rect 2200 17661 2212 17817
rect 2264 17661 2377 17817
rect 2200 17649 2377 17661
rect 2116 16935 2244 17031
rect 2116 16879 2152 16935
rect 2208 16879 2244 16935
rect 2116 16802 2244 16879
rect 2462 16754 2518 22154
rect 2778 22150 2834 23751
rect 2711 22094 2834 22150
rect 2711 20408 2767 22094
rect 2846 22020 2922 22032
rect 2846 22009 2858 22020
rect 2910 22009 2922 22020
rect 2846 21849 2856 22009
rect 2912 21849 2922 22009
rect 2846 21839 2922 21849
rect 2988 21824 3044 26223
rect 3174 21824 3230 26223
rect 3604 25363 3660 26223
rect 3582 25351 3660 25363
rect 3582 25195 3594 25351
rect 3646 25195 3660 25351
rect 3582 25183 3660 25195
rect 3796 25363 3852 26223
rect 3796 25351 3874 25363
rect 3796 25195 3810 25351
rect 3862 25195 3874 25351
rect 3796 25183 3874 25195
rect 3690 24679 3766 24689
rect 3690 24415 3700 24679
rect 3756 24415 3766 24679
rect 3690 24405 3766 24415
rect 3374 23919 3450 23931
rect 3374 23763 3386 23919
rect 3438 23763 3450 23919
rect 3374 23751 3450 23763
rect 4006 23919 4082 23931
rect 4006 23763 4018 23919
rect 4070 23763 4082 23919
rect 4006 23751 4082 23763
rect 3384 22150 3440 23751
rect 3589 22218 3867 22230
rect 3589 22166 3601 22218
rect 3653 22166 3803 22218
rect 3855 22166 3867 22218
rect 3589 22154 3867 22166
rect 3384 22094 3507 22150
rect 3296 22020 3372 22032
rect 3296 22009 3308 22020
rect 3360 22009 3372 22020
rect 3296 21849 3306 22009
rect 3362 21849 3372 22009
rect 3296 21839 3372 21849
rect 2978 21812 3054 21824
rect 2978 21760 2990 21812
rect 3042 21760 3054 21812
rect 2978 21748 3054 21760
rect 3164 21812 3240 21824
rect 3164 21760 3176 21812
rect 3228 21760 3240 21812
rect 3164 21748 3240 21760
rect 2603 20352 2767 20408
rect 2603 19950 2659 20352
rect 2971 20236 3063 21270
rect 2740 20212 3063 20236
rect 2740 20160 2776 20212
rect 2828 20160 3063 20212
rect 2740 20139 3063 20160
rect 2762 19950 2838 19960
rect 2603 19948 2838 19950
rect 2603 19896 2774 19948
rect 2826 19896 2838 19948
rect 2603 19894 2838 19896
rect 2603 17829 2659 19894
rect 2762 19884 2838 19894
rect 2971 19596 3063 20139
rect 3155 20256 3247 21270
rect 3451 20408 3507 22094
rect 3451 20352 3615 20408
rect 3155 20236 3249 20256
rect 3155 20218 3478 20236
rect 3155 20162 3174 20218
rect 3230 20212 3478 20218
rect 3230 20162 3390 20212
rect 3155 20160 3390 20162
rect 3442 20160 3478 20212
rect 3155 20139 3478 20160
rect 3155 20123 3249 20139
rect 2970 19558 3064 19596
rect 2970 19502 2989 19558
rect 3045 19502 3064 19558
rect 2970 19463 3064 19502
rect 2971 18606 3063 19463
rect 2764 18509 3063 18606
rect 3155 18606 3247 20123
rect 3380 19950 3456 19960
rect 3559 19950 3615 20352
rect 3380 19948 3615 19950
rect 3380 19896 3392 19948
rect 3444 19896 3615 19948
rect 3380 19894 3615 19896
rect 3380 19884 3456 19894
rect 3155 18509 3454 18606
rect 2764 17980 2840 18509
rect 2955 18380 3263 18400
rect 2955 18328 2985 18380
rect 3037 18328 3171 18380
rect 3223 18328 3263 18380
rect 2955 18308 3263 18328
rect 2764 17928 2776 17980
rect 2828 17928 2840 17980
rect 2764 17908 2840 17928
rect 2926 18173 3002 18195
rect 2926 18013 2936 18173
rect 2992 18013 3002 18173
rect 2926 17913 3002 18013
rect 2603 17817 2780 17829
rect 2603 17661 2716 17817
rect 2768 17661 2780 17817
rect 2603 17649 2780 17661
rect 2736 16935 2864 17031
rect 2736 16879 2772 16935
rect 2828 16879 2864 16935
rect 2736 16802 2864 16879
rect 1715 16616 2023 16636
rect 1715 16564 1745 16616
rect 1797 16564 1931 16616
rect 1983 16564 2023 16616
rect 1715 16544 2023 16564
rect 2446 16428 2535 16754
rect 3065 16639 3154 18308
rect 3217 18173 3293 18195
rect 3217 18013 3227 18173
rect 3283 18013 3293 18173
rect 3217 17913 3293 18013
rect 3378 17980 3454 18509
rect 3378 17928 3390 17980
rect 3442 17928 3454 17980
rect 3378 17908 3454 17928
rect 3559 17829 3615 19894
rect 3438 17817 3615 17829
rect 3438 17661 3450 17817
rect 3502 17661 3615 17817
rect 3438 17649 3615 17661
rect 3354 16935 3482 17031
rect 3354 16879 3390 16935
rect 3446 16879 3482 16935
rect 3354 16802 3482 16879
rect 3700 16752 3756 22154
rect 4016 22150 4072 23751
rect 3949 22094 4072 22150
rect 3949 20408 4005 22094
rect 4084 22020 4160 22032
rect 4084 22009 4096 22020
rect 4148 22009 4160 22020
rect 4084 21849 4094 22009
rect 4150 21849 4160 22009
rect 4084 21839 4160 21849
rect 4226 21824 4282 26223
rect 4413 21824 4469 26223
rect 4843 25363 4899 26223
rect 4821 25351 4899 25363
rect 4821 25195 4833 25351
rect 4885 25195 4899 25351
rect 4821 25183 4899 25195
rect 5039 25363 5095 26223
rect 5039 25351 5117 25363
rect 5039 25195 5053 25351
rect 5105 25195 5117 25351
rect 5039 25183 5117 25195
rect 4929 24679 5005 24689
rect 4929 24415 4939 24679
rect 4995 24415 5005 24679
rect 4929 24405 5005 24415
rect 4613 23919 4689 23931
rect 4613 23763 4625 23919
rect 4677 23763 4689 23919
rect 4613 23751 4689 23763
rect 5245 23919 5321 23931
rect 5245 23763 5257 23919
rect 5309 23763 5321 23919
rect 5245 23751 5321 23763
rect 4623 22150 4679 23751
rect 4828 22218 5106 22230
rect 4828 22166 4840 22218
rect 4892 22166 5042 22218
rect 5094 22166 5106 22218
rect 4828 22154 5106 22166
rect 5255 22157 5311 23751
rect 4623 22094 4746 22150
rect 4535 22020 4611 22032
rect 4535 22009 4547 22020
rect 4599 22009 4611 22020
rect 4535 21849 4545 22009
rect 4601 21849 4611 22009
rect 4535 21839 4611 21849
rect 4216 21812 4292 21824
rect 4216 21760 4228 21812
rect 4280 21760 4292 21812
rect 4216 21748 4292 21760
rect 4403 21812 4479 21824
rect 4403 21760 4415 21812
rect 4467 21760 4479 21812
rect 4403 21748 4479 21760
rect 3841 20352 4005 20408
rect 4209 20569 4301 21270
rect 4394 20898 4486 21270
rect 4393 20860 4487 20898
rect 4393 20804 4412 20860
rect 4468 20804 4487 20860
rect 4393 20765 4487 20804
rect 4209 20531 4303 20569
rect 4209 20475 4228 20531
rect 4284 20475 4303 20531
rect 4209 20436 4303 20475
rect 3841 19950 3897 20352
rect 4209 20236 4301 20436
rect 3978 20212 4301 20236
rect 3978 20160 4014 20212
rect 4066 20160 4301 20212
rect 3978 20139 4301 20160
rect 4000 19950 4076 19960
rect 3841 19948 4076 19950
rect 3841 19896 4012 19948
rect 4064 19896 4076 19948
rect 3841 19894 4076 19896
rect 3841 17829 3897 19894
rect 4000 19884 4076 19894
rect 4209 18606 4301 20139
rect 4002 18509 4301 18606
rect 4394 20236 4486 20765
rect 4690 20408 4746 22094
rect 4690 20352 4854 20408
rect 4394 20212 4717 20236
rect 4394 20160 4629 20212
rect 4681 20160 4717 20212
rect 4394 20139 4717 20160
rect 4394 18606 4486 20139
rect 4619 19950 4695 19960
rect 4798 19950 4854 20352
rect 4619 19948 4854 19950
rect 4619 19896 4631 19948
rect 4683 19896 4854 19948
rect 4619 19894 4854 19896
rect 4619 19884 4695 19894
rect 4394 18509 4693 18606
rect 4002 17980 4078 18509
rect 4194 18380 4502 18400
rect 4194 18328 4224 18380
rect 4276 18328 4410 18380
rect 4462 18328 4502 18380
rect 4194 18308 4502 18328
rect 4002 17928 4014 17980
rect 4066 17928 4078 17980
rect 4002 17908 4078 17928
rect 4164 18173 4240 18195
rect 4164 18013 4174 18173
rect 4230 18013 4240 18173
rect 4164 17913 4240 18013
rect 3841 17817 4018 17829
rect 3841 17661 3954 17817
rect 4006 17661 4018 17817
rect 3841 17649 4018 17661
rect 3974 16935 4102 17031
rect 3974 16879 4010 16935
rect 4066 16879 4102 16935
rect 3974 16802 4102 16879
rect 4303 16639 4393 18308
rect 4455 18173 4531 18195
rect 4455 18013 4465 18173
rect 4521 18013 4531 18173
rect 4455 17913 4531 18013
rect 4617 17980 4693 18509
rect 4617 17928 4629 17980
rect 4681 17928 4693 17980
rect 4617 17908 4693 17928
rect 4798 17829 4854 19894
rect 4677 17817 4854 17829
rect 4677 17661 4689 17817
rect 4741 17661 4854 17817
rect 4677 17649 4854 17661
rect 4593 16935 4721 17031
rect 4593 16879 4629 16935
rect 4685 16879 4721 16935
rect 4593 16802 4721 16879
rect 4939 16752 4995 22154
rect 5179 22101 5311 22157
rect 5179 20408 5235 22101
rect 5315 22027 5391 22039
rect 5315 22016 5327 22027
rect 5379 22016 5391 22027
rect 5315 21856 5325 22016
rect 5381 21856 5391 22016
rect 5315 21846 5391 21856
rect 5457 21823 5513 26223
rect 5447 21811 5523 21823
rect 5447 21759 5459 21811
rect 5511 21759 5523 21811
rect 5447 21747 5523 21759
rect 5080 20352 5235 20408
rect 5447 21217 5541 21270
rect 5447 21179 5542 21217
rect 5447 21123 5467 21179
rect 5523 21123 5542 21179
rect 5447 21084 5542 21123
rect 5080 19950 5136 20352
rect 5447 20236 5541 21084
rect 5217 20212 5541 20236
rect 5217 20160 5253 20212
rect 5305 20160 5541 20212
rect 5217 20139 5541 20160
rect 5239 19950 5315 19961
rect 5080 19949 5315 19950
rect 5080 19897 5251 19949
rect 5303 19897 5315 19949
rect 5080 19894 5315 19897
rect 5080 17829 5136 19894
rect 5239 19885 5315 19894
rect 5447 18606 5541 20139
rect 5242 18509 5541 18606
rect 5242 17981 5318 18509
rect 5389 18380 5522 18401
rect 5389 18328 5429 18380
rect 5481 18328 5522 18380
rect 5389 18308 5522 18328
rect 5242 17929 5254 17981
rect 5306 17929 5318 17981
rect 5242 17908 5318 17929
rect 5080 17817 5238 17829
rect 5080 17661 5174 17817
rect 5226 17661 5238 17817
rect 5080 17649 5238 17661
rect 5212 16935 5341 17031
rect 5212 16879 5249 16935
rect 5305 16879 5341 16935
rect 5212 16802 5341 16879
rect 5432 16432 5522 18308
rect 5045 16428 5522 16432
rect 2316 16408 2624 16428
rect 2316 16356 2346 16408
rect 2398 16356 2532 16408
rect 2584 16356 2624 16408
rect 2316 16336 2624 16356
rect 4824 16408 5522 16428
rect 4824 16356 4854 16408
rect 4906 16356 5040 16408
rect 5092 16356 5522 16408
rect 4824 16336 5522 16356
rect 2446 16335 2535 16336
rect 5045 16335 5522 16336
rect 1768 16182 3373 16220
rect 1768 16126 1804 16182
rect 1860 16126 2015 16182
rect 2071 16126 2225 16182
rect 2281 16126 2436 16182
rect 2492 16126 2648 16182
rect 2704 16126 2859 16182
rect 2915 16126 3069 16182
rect 3125 16126 3280 16182
rect 3336 16126 3373 16182
rect 1768 16087 3373 16126
rect 3720 16182 4482 16220
rect 3720 16126 3756 16182
rect 3812 16126 3967 16182
rect 4023 16126 4179 16182
rect 4235 16126 4390 16182
rect 4446 16126 4482 16182
rect 3720 16087 4482 16126
rect 1398 15734 1608 15775
rect 1398 15682 1419 15734
rect 1471 15682 1608 15734
rect 1398 15678 1608 15682
rect 1398 15548 1492 15678
rect 1398 15496 1419 15548
rect 1471 15496 1492 15548
rect 1398 15455 1492 15496
rect 1627 15560 1935 15578
rect 1627 15504 1655 15560
rect 1711 15504 1841 15560
rect 1897 15504 1935 15560
rect 1627 15486 1935 15504
rect 1357 15142 1449 15170
rect 1357 15086 1375 15142
rect 1431 15086 1449 15142
rect 1357 14956 1449 15086
rect 1357 14900 1375 14956
rect 1431 14900 1449 14956
rect 1357 14862 1449 14900
rect 1847 15042 1939 15070
rect 1847 14986 1865 15042
rect 1921 14986 1939 15042
rect 1847 14856 1939 14986
rect 1847 14800 1865 14856
rect 1921 14800 1939 14856
rect 1847 14762 1939 14800
rect 1172 14299 1193 14351
rect 1245 14299 1266 14351
rect 1172 14165 1266 14299
rect 1172 14113 1193 14165
rect 1245 14113 1266 14165
rect 1172 12560 1266 14113
rect 1847 13551 1939 13579
rect 1847 13495 1865 13551
rect 1921 13495 1939 13551
rect 1847 13365 1939 13495
rect 1847 13309 1865 13365
rect 1921 13309 1939 13365
rect 1847 13271 1939 13309
rect 2072 12624 2166 15972
rect 1172 12508 1193 12560
rect 1245 12508 1266 12560
rect 1172 12374 1266 12508
rect 1172 12322 1193 12374
rect 1245 12322 1266 12374
rect 1172 12282 1266 12322
rect 1834 12556 1926 12584
rect 1834 12500 1852 12556
rect 1908 12500 1926 12556
rect 1834 12370 1926 12500
rect 1834 12314 1852 12370
rect 1908 12314 1926 12370
rect 1834 12276 1926 12314
rect 2072 12568 2091 12624
rect 2147 12568 2166 12624
rect 2072 12438 2166 12568
rect 2072 12382 2091 12438
rect 2147 12382 2166 12438
rect 2072 11849 2166 12382
rect 2072 11793 2091 11849
rect 2147 11793 2166 11849
rect 2072 11663 2166 11793
rect 1834 11608 1926 11636
rect 1834 11552 1852 11608
rect 1908 11552 1926 11608
rect 1834 11422 1926 11552
rect 1834 11366 1852 11422
rect 1908 11366 1926 11422
rect 1834 11328 1926 11366
rect 2072 11607 2091 11663
rect 2147 11607 2166 11663
rect 2072 10933 2166 11607
rect 2072 10877 2091 10933
rect 2147 10877 2166 10933
rect 2072 10747 2166 10877
rect 1834 10692 1926 10720
rect 1834 10636 1852 10692
rect 1908 10636 1926 10692
rect 1834 10506 1926 10636
rect 1834 10450 1852 10506
rect 1908 10450 1926 10506
rect 1834 10412 1926 10450
rect 2072 10691 2091 10747
rect 2147 10691 2166 10747
rect 943 10248 1070 10269
rect 2072 10257 2166 10691
rect 2256 15929 2351 15970
rect 2256 15877 2278 15929
rect 2330 15877 2351 15929
rect 2256 15743 2351 15877
rect 2256 15691 2278 15743
rect 2330 15691 2351 15743
rect 943 10196 978 10248
rect 1030 10196 1913 10248
rect 943 10192 1913 10196
rect 943 10176 1070 10192
rect 898 9840 990 9868
rect 898 9784 916 9840
rect 972 9784 990 9840
rect 898 9654 990 9784
rect 1616 9840 1708 9868
rect 1616 9784 1634 9840
rect 1690 9784 1708 9840
rect 898 9598 916 9654
rect 972 9598 990 9654
rect 898 9560 990 9598
rect 1420 9695 1514 9733
rect 1420 9639 1439 9695
rect 1495 9639 1514 9695
rect 258 9520 598 9559
rect 258 9464 294 9520
rect 350 9464 506 9520
rect 562 9464 598 9520
rect 258 9425 598 9464
rect 1420 9509 1514 9639
rect 1616 9654 1708 9784
rect 1616 9598 1634 9654
rect 1690 9598 1708 9654
rect 1616 9560 1708 9598
rect 1420 9453 1439 9509
rect 1495 9453 1514 9509
rect 573 9099 881 9117
rect 573 9043 601 9099
rect 657 9043 787 9099
rect 843 9043 881 9099
rect 573 9025 881 9043
rect 1221 9082 1313 9120
rect 1221 9026 1239 9082
rect 1295 9026 1313 9082
rect 277 8983 369 9011
rect 277 8927 295 8983
rect 351 8927 369 8983
rect 277 8797 369 8927
rect 1221 8896 1313 9026
rect 277 8741 295 8797
rect 351 8741 369 8797
rect 617 8863 926 8883
rect 617 8811 647 8863
rect 699 8811 833 8863
rect 885 8811 926 8863
rect 1221 8840 1239 8896
rect 1295 8840 1313 8896
rect 1221 8812 1313 8840
rect 617 8791 926 8811
rect 277 8703 369 8741
rect 461 8523 553 8563
rect 461 8471 481 8523
rect 533 8471 553 8523
rect 461 8427 553 8471
rect 460 8337 554 8427
rect 460 8285 481 8337
rect 533 8285 554 8337
rect 460 -1 554 8285
rect 831 7768 926 8791
rect 1039 8733 1131 8771
rect 1039 8677 1057 8733
rect 1113 8677 1131 8733
rect 1039 8547 1131 8677
rect 1039 8491 1057 8547
rect 1113 8491 1131 8547
rect 1039 8463 1131 8491
rect 1017 8121 1110 8136
rect 1420 8121 1514 9453
rect 1610 9082 1702 9120
rect 1610 9026 1628 9082
rect 1684 9026 1702 9082
rect 1610 8896 1702 9026
rect 1610 8840 1628 8896
rect 1684 8840 1702 8896
rect 1610 8812 1702 8840
rect 1016 8096 1514 8121
rect 1016 8044 1037 8096
rect 1089 8044 1514 8096
rect 1016 8024 1514 8044
rect 1017 8004 1110 8024
rect 831 7634 1158 7768
rect 1063 5917 1158 7634
rect 1857 7689 1913 10192
rect 2043 9266 2135 9306
rect 2043 9214 2063 9266
rect 2115 9214 2135 9266
rect 2043 9121 2135 9214
rect 2042 9082 2135 9121
rect 2042 9026 2061 9082
rect 2117 9026 2135 9082
rect 2042 8896 2135 9026
rect 2042 8840 2061 8896
rect 2117 8840 2135 8896
rect 2042 8802 2135 8840
rect 2256 7803 2351 15691
rect 2441 12624 2535 15972
rect 2441 12568 2460 12624
rect 2516 12568 2535 12624
rect 2441 12438 2535 12568
rect 2441 12382 2460 12438
rect 2516 12382 2535 12438
rect 2441 11849 2535 12382
rect 2441 11793 2460 11849
rect 2516 11793 2535 11849
rect 2441 11663 2535 11793
rect 2441 11607 2460 11663
rect 2516 11607 2535 11663
rect 2441 10933 2535 11607
rect 2441 10877 2460 10933
rect 2516 10877 2535 10933
rect 2441 10747 2535 10877
rect 2441 10691 2460 10747
rect 2516 10691 2535 10747
rect 2441 10257 2535 10691
rect 5345 10239 5437 10279
rect 5345 10187 5365 10239
rect 5417 10187 5437 10239
rect 5345 10100 5437 10187
rect 5344 10053 5438 10100
rect 5344 10001 5365 10053
rect 5417 10001 5438 10053
rect 2772 9935 2864 9963
rect 2772 9879 2790 9935
rect 2846 9879 2864 9935
rect 2772 9749 2864 9879
rect 2772 9693 2790 9749
rect 2846 9693 2864 9749
rect 2772 9655 2864 9693
rect 2772 9012 2864 9040
rect 2772 8956 2790 9012
rect 2846 8956 2864 9012
rect 2772 8826 2864 8956
rect 2772 8770 2790 8826
rect 2846 8770 2864 8826
rect 2772 8732 2864 8770
rect 4233 8339 4327 8518
rect 4692 8470 4786 8518
rect 4692 8373 5050 8470
rect 4233 8242 4435 8339
rect 4956 8158 5050 8373
rect 1857 7633 2004 7689
rect 2256 7687 2863 7803
rect 1497 6674 1591 6675
rect 1485 6634 1591 6674
rect 1485 6582 1505 6634
rect 1557 6582 1591 6634
rect 1485 6448 1591 6582
rect 1485 6396 1505 6448
rect 1557 6396 1591 6448
rect 1485 6356 1591 6396
rect 845 5811 1158 5917
rect 845 1505 940 5811
rect 1497 5738 1591 6356
rect 1948 6076 2004 7633
rect 1308 5625 1591 5738
rect 1877 6020 2004 6076
rect 911 -89 1006 1366
rect 1308 1 1402 5625
rect 1877 1853 1933 6020
rect 2298 4999 2354 5859
rect 2768 5039 2863 7687
rect 5344 6043 5438 10001
rect 4370 5909 4715 6043
rect 4639 5591 4715 5909
rect 4639 5435 4651 5591
rect 4703 5435 4715 5591
rect 4639 5423 4715 5435
rect 5125 5909 5438 6043
rect 5125 5591 5201 5909
rect 5125 5435 5137 5591
rect 5189 5435 5201 5591
rect 5125 5423 5201 5435
rect 2131 4989 2354 4999
rect 2131 4933 2141 4989
rect 2301 4933 2354 4989
rect 2466 4948 2863 5039
rect 2131 4923 2311 4933
rect 2466 4680 2577 4948
rect 2256 4594 2577 4680
rect 2256 3604 2351 4594
rect 2256 3552 2277 3604
rect 2329 3552 2351 3604
rect 2256 3418 2351 3552
rect 2256 3366 2277 3418
rect 2329 3366 2351 3418
rect 2256 3325 2351 3366
rect 1877 1797 1984 1853
rect 1928 986 1984 1797
rect 1928 910 2054 986
rect 866 -101 1046 -89
rect 866 -153 878 -101
rect 1034 -153 1046 -101
rect 866 -165 1046 -153
rect 1998 -1907 2054 910
rect 1998 -1963 3066 -1907
rect 3010 -2254 3066 -1963
rect 3000 -2266 3076 -2254
rect 3000 -2422 3012 -2266
rect 3064 -2422 3076 -2266
rect 3000 -2434 3076 -2422
<< via2 >>
rect 916 28956 972 28958
rect 916 28904 918 28956
rect 918 28904 970 28956
rect 970 28904 972 28956
rect 916 28902 972 28904
rect 916 28770 972 28772
rect 916 28718 918 28770
rect 918 28718 970 28770
rect 970 28718 972 28770
rect 916 28716 972 28718
rect 99 22570 155 22626
rect 99 22384 155 22440
rect 1530 28956 1586 28958
rect 1530 28904 1532 28956
rect 1532 28904 1584 28956
rect 1584 28904 1586 28956
rect 1530 28902 1586 28904
rect 1530 28770 1586 28772
rect 1530 28718 1532 28770
rect 1532 28718 1584 28770
rect 1584 28718 1586 28770
rect 1530 28716 1586 28718
rect 2155 28956 2211 28958
rect 2155 28904 2157 28956
rect 2157 28904 2209 28956
rect 2209 28904 2211 28956
rect 2155 28902 2211 28904
rect 2155 28770 2211 28772
rect 2155 28718 2157 28770
rect 2157 28718 2209 28770
rect 2209 28718 2211 28770
rect 2155 28716 2211 28718
rect 2769 28956 2825 28958
rect 2769 28904 2771 28956
rect 2771 28904 2823 28956
rect 2823 28904 2825 28956
rect 2769 28902 2825 28904
rect 2769 28770 2825 28772
rect 2769 28718 2771 28770
rect 2771 28718 2823 28770
rect 2823 28718 2825 28770
rect 2769 28716 2825 28718
rect 3393 28956 3449 28958
rect 3393 28904 3395 28956
rect 3395 28904 3447 28956
rect 3447 28904 3449 28956
rect 3393 28902 3449 28904
rect 3393 28770 3449 28772
rect 3393 28718 3395 28770
rect 3395 28718 3447 28770
rect 3447 28718 3449 28770
rect 3393 28716 3449 28718
rect 4007 28956 4063 28958
rect 4007 28904 4009 28956
rect 4009 28904 4061 28956
rect 4061 28904 4063 28956
rect 4007 28902 4063 28904
rect 4007 28770 4063 28772
rect 4007 28718 4009 28770
rect 4009 28718 4061 28770
rect 4061 28718 4063 28770
rect 4007 28716 4063 28718
rect 4632 28956 4688 28958
rect 4632 28904 4634 28956
rect 4634 28904 4686 28956
rect 4686 28904 4688 28956
rect 4632 28902 4688 28904
rect 4632 28770 4688 28772
rect 4632 28718 4634 28770
rect 4634 28718 4686 28770
rect 4686 28718 4688 28770
rect 4632 28716 4688 28718
rect 5246 28956 5302 28958
rect 5246 28904 5248 28956
rect 5248 28904 5300 28956
rect 5300 28904 5302 28956
rect 5246 28902 5302 28904
rect 5246 28770 5302 28772
rect 5246 28718 5248 28770
rect 5248 28718 5300 28770
rect 5300 28718 5302 28770
rect 5246 28716 5302 28718
rect 492 22570 548 22626
rect 492 22384 548 22440
rect 1223 24677 1279 24679
rect 1223 24417 1225 24677
rect 1225 24417 1277 24677
rect 1277 24417 1279 24677
rect 1223 24415 1279 24417
rect 829 21968 831 22009
rect 831 21968 883 22009
rect 883 21968 885 22009
rect 829 21849 885 21968
rect 697 18548 753 18604
rect 913 16933 969 16935
rect 913 16881 915 16933
rect 915 16881 967 16933
rect 967 16881 969 16933
rect 913 16879 969 16881
rect 1617 21968 1619 22009
rect 1619 21968 1671 22009
rect 1671 21968 1673 22009
rect 1617 21849 1673 21968
rect 2462 24677 2518 24679
rect 2462 24417 2464 24677
rect 2464 24417 2516 24677
rect 2516 24417 2518 24677
rect 2462 24415 2518 24417
rect 2068 21968 2070 22009
rect 2070 21968 2122 22009
rect 2122 21968 2124 22009
rect 2068 21849 2124 21968
rect 1935 19190 1991 19246
rect 1751 18863 1807 18919
rect 1697 18171 1753 18173
rect 1697 18119 1699 18171
rect 1699 18119 1751 18171
rect 1751 18119 1753 18171
rect 1697 18013 1753 18119
rect 1533 16933 1589 16935
rect 1533 16881 1535 16933
rect 1535 16881 1587 16933
rect 1587 16881 1589 16933
rect 1533 16879 1589 16881
rect 295 15605 351 15607
rect 295 15553 297 15605
rect 297 15553 349 15605
rect 349 15553 351 15605
rect 295 15551 351 15553
rect 295 15419 351 15421
rect 295 15367 297 15419
rect 297 15367 349 15419
rect 349 15367 351 15419
rect 295 15365 351 15367
rect 295 15006 351 15008
rect 295 14954 297 15006
rect 297 14954 349 15006
rect 349 14954 351 15006
rect 295 14952 351 14954
rect 295 14820 351 14822
rect 295 14768 297 14820
rect 297 14768 349 14820
rect 349 14768 351 14820
rect 295 14766 351 14768
rect 965 16183 1021 16185
rect 965 16131 967 16183
rect 967 16131 1019 16183
rect 1019 16131 1021 16183
rect 965 16129 1021 16131
rect 295 13549 351 13551
rect 295 13497 297 13549
rect 297 13497 349 13549
rect 349 13497 351 13549
rect 295 13495 351 13497
rect 295 13363 351 13365
rect 295 13311 297 13363
rect 297 13311 349 13363
rect 349 13311 351 13363
rect 295 13309 351 13311
rect 295 12554 351 12556
rect 295 12502 297 12554
rect 297 12502 349 12554
rect 349 12502 351 12554
rect 295 12500 351 12502
rect 295 12368 351 12370
rect 295 12316 297 12368
rect 297 12316 349 12368
rect 349 12316 351 12368
rect 295 12314 351 12316
rect 295 11606 351 11608
rect 295 11554 297 11606
rect 297 11554 349 11606
rect 349 11554 351 11606
rect 295 11552 351 11554
rect 295 11420 351 11422
rect 295 11368 297 11420
rect 297 11368 349 11420
rect 349 11368 351 11420
rect 295 11366 351 11368
rect 295 10690 351 10692
rect 295 10638 297 10690
rect 297 10638 349 10690
rect 349 10638 351 10690
rect 295 10636 351 10638
rect 295 10504 351 10506
rect 295 10452 297 10504
rect 297 10452 349 10504
rect 349 10452 351 10504
rect 295 10450 351 10452
rect 1988 18171 2044 18173
rect 1988 18119 1990 18171
rect 1990 18119 2042 18171
rect 2042 18119 2044 18171
rect 1988 18013 2044 18119
rect 2152 16933 2208 16935
rect 2152 16881 2154 16933
rect 2154 16881 2206 16933
rect 2206 16881 2208 16933
rect 2152 16879 2208 16881
rect 2856 21968 2858 22009
rect 2858 21968 2910 22009
rect 2910 21968 2912 22009
rect 2856 21849 2912 21968
rect 3700 24677 3756 24679
rect 3700 24417 3702 24677
rect 3702 24417 3754 24677
rect 3754 24417 3756 24677
rect 3700 24415 3756 24417
rect 3306 21968 3308 22009
rect 3308 21968 3360 22009
rect 3360 21968 3362 22009
rect 3306 21849 3362 21968
rect 3174 20162 3230 20218
rect 2989 19502 3045 19558
rect 2936 18171 2992 18173
rect 2936 18119 2938 18171
rect 2938 18119 2990 18171
rect 2990 18119 2992 18171
rect 2936 18013 2992 18119
rect 2772 16933 2828 16935
rect 2772 16881 2774 16933
rect 2774 16881 2826 16933
rect 2826 16881 2828 16933
rect 2772 16879 2828 16881
rect 3227 18171 3283 18173
rect 3227 18119 3229 18171
rect 3229 18119 3281 18171
rect 3281 18119 3283 18171
rect 3227 18013 3283 18119
rect 3390 16933 3446 16935
rect 3390 16881 3392 16933
rect 3392 16881 3444 16933
rect 3444 16881 3446 16933
rect 3390 16879 3446 16881
rect 4094 21968 4096 22009
rect 4096 21968 4148 22009
rect 4148 21968 4150 22009
rect 4094 21849 4150 21968
rect 4939 24677 4995 24679
rect 4939 24417 4941 24677
rect 4941 24417 4993 24677
rect 4993 24417 4995 24677
rect 4939 24415 4995 24417
rect 4545 21968 4547 22009
rect 4547 21968 4599 22009
rect 4599 21968 4601 22009
rect 4545 21849 4601 21968
rect 4412 20804 4468 20860
rect 4228 20475 4284 20531
rect 4174 18171 4230 18173
rect 4174 18119 4176 18171
rect 4176 18119 4228 18171
rect 4228 18119 4230 18171
rect 4174 18013 4230 18119
rect 4010 16933 4066 16935
rect 4010 16881 4012 16933
rect 4012 16881 4064 16933
rect 4064 16881 4066 16933
rect 4010 16879 4066 16881
rect 4465 18171 4521 18173
rect 4465 18119 4467 18171
rect 4467 18119 4519 18171
rect 4519 18119 4521 18171
rect 4465 18013 4521 18119
rect 4629 16933 4685 16935
rect 4629 16881 4631 16933
rect 4631 16881 4683 16933
rect 4683 16881 4685 16933
rect 4629 16879 4685 16881
rect 5325 21975 5327 22016
rect 5327 21975 5379 22016
rect 5379 21975 5381 22016
rect 5325 21856 5381 21975
rect 5467 21123 5523 21179
rect 5249 16933 5305 16935
rect 5249 16881 5251 16933
rect 5251 16881 5303 16933
rect 5303 16881 5305 16933
rect 5249 16879 5305 16881
rect 1804 16180 1860 16182
rect 1804 16128 1806 16180
rect 1806 16128 1858 16180
rect 1858 16128 1860 16180
rect 1804 16126 1860 16128
rect 2015 16180 2071 16182
rect 2015 16128 2017 16180
rect 2017 16128 2069 16180
rect 2069 16128 2071 16180
rect 2015 16126 2071 16128
rect 2225 16180 2281 16182
rect 2225 16128 2227 16180
rect 2227 16128 2279 16180
rect 2279 16128 2281 16180
rect 2225 16126 2281 16128
rect 2436 16180 2492 16182
rect 2436 16128 2438 16180
rect 2438 16128 2490 16180
rect 2490 16128 2492 16180
rect 2436 16126 2492 16128
rect 2648 16180 2704 16182
rect 2648 16128 2650 16180
rect 2650 16128 2702 16180
rect 2702 16128 2704 16180
rect 2648 16126 2704 16128
rect 2859 16180 2915 16182
rect 2859 16128 2861 16180
rect 2861 16128 2913 16180
rect 2913 16128 2915 16180
rect 2859 16126 2915 16128
rect 3069 16180 3125 16182
rect 3069 16128 3071 16180
rect 3071 16128 3123 16180
rect 3123 16128 3125 16180
rect 3069 16126 3125 16128
rect 3280 16180 3336 16182
rect 3280 16128 3282 16180
rect 3282 16128 3334 16180
rect 3334 16128 3336 16180
rect 3280 16126 3336 16128
rect 3756 16180 3812 16182
rect 3756 16128 3758 16180
rect 3758 16128 3810 16180
rect 3810 16128 3812 16180
rect 3756 16126 3812 16128
rect 3967 16180 4023 16182
rect 3967 16128 3969 16180
rect 3969 16128 4021 16180
rect 4021 16128 4023 16180
rect 3967 16126 4023 16128
rect 4179 16180 4235 16182
rect 4179 16128 4181 16180
rect 4181 16128 4233 16180
rect 4233 16128 4235 16180
rect 4179 16126 4235 16128
rect 4390 16180 4446 16182
rect 4390 16128 4392 16180
rect 4392 16128 4444 16180
rect 4444 16128 4446 16180
rect 4390 16126 4446 16128
rect 1655 15558 1711 15560
rect 1655 15506 1657 15558
rect 1657 15506 1709 15558
rect 1709 15506 1711 15558
rect 1655 15504 1711 15506
rect 1841 15558 1897 15560
rect 1841 15506 1843 15558
rect 1843 15506 1895 15558
rect 1895 15506 1897 15558
rect 1841 15504 1897 15506
rect 1375 15140 1431 15142
rect 1375 15088 1377 15140
rect 1377 15088 1429 15140
rect 1429 15088 1431 15140
rect 1375 15086 1431 15088
rect 1375 14954 1431 14956
rect 1375 14902 1377 14954
rect 1377 14902 1429 14954
rect 1429 14902 1431 14954
rect 1375 14900 1431 14902
rect 1865 15040 1921 15042
rect 1865 14988 1867 15040
rect 1867 14988 1919 15040
rect 1919 14988 1921 15040
rect 1865 14986 1921 14988
rect 1865 14854 1921 14856
rect 1865 14802 1867 14854
rect 1867 14802 1919 14854
rect 1919 14802 1921 14854
rect 1865 14800 1921 14802
rect 1865 13549 1921 13551
rect 1865 13497 1867 13549
rect 1867 13497 1919 13549
rect 1919 13497 1921 13549
rect 1865 13495 1921 13497
rect 1865 13363 1921 13365
rect 1865 13311 1867 13363
rect 1867 13311 1919 13363
rect 1919 13311 1921 13363
rect 1865 13309 1921 13311
rect 1852 12554 1908 12556
rect 1852 12502 1854 12554
rect 1854 12502 1906 12554
rect 1906 12502 1908 12554
rect 1852 12500 1908 12502
rect 1852 12368 1908 12370
rect 1852 12316 1854 12368
rect 1854 12316 1906 12368
rect 1906 12316 1908 12368
rect 1852 12314 1908 12316
rect 2091 12622 2147 12624
rect 2091 12570 2093 12622
rect 2093 12570 2145 12622
rect 2145 12570 2147 12622
rect 2091 12568 2147 12570
rect 2091 12436 2147 12438
rect 2091 12384 2093 12436
rect 2093 12384 2145 12436
rect 2145 12384 2147 12436
rect 2091 12382 2147 12384
rect 2091 11847 2147 11849
rect 2091 11795 2093 11847
rect 2093 11795 2145 11847
rect 2145 11795 2147 11847
rect 2091 11793 2147 11795
rect 1852 11606 1908 11608
rect 1852 11554 1854 11606
rect 1854 11554 1906 11606
rect 1906 11554 1908 11606
rect 1852 11552 1908 11554
rect 1852 11420 1908 11422
rect 1852 11368 1854 11420
rect 1854 11368 1906 11420
rect 1906 11368 1908 11420
rect 1852 11366 1908 11368
rect 2091 11661 2147 11663
rect 2091 11609 2093 11661
rect 2093 11609 2145 11661
rect 2145 11609 2147 11661
rect 2091 11607 2147 11609
rect 2091 10931 2147 10933
rect 2091 10879 2093 10931
rect 2093 10879 2145 10931
rect 2145 10879 2147 10931
rect 2091 10877 2147 10879
rect 1852 10690 1908 10692
rect 1852 10638 1854 10690
rect 1854 10638 1906 10690
rect 1906 10638 1908 10690
rect 1852 10636 1908 10638
rect 1852 10504 1908 10506
rect 1852 10452 1854 10504
rect 1854 10452 1906 10504
rect 1906 10452 1908 10504
rect 1852 10450 1908 10452
rect 2091 10745 2147 10747
rect 2091 10693 2093 10745
rect 2093 10693 2145 10745
rect 2145 10693 2147 10745
rect 2091 10691 2147 10693
rect 916 9838 972 9840
rect 916 9786 918 9838
rect 918 9786 970 9838
rect 970 9786 972 9838
rect 916 9784 972 9786
rect 1634 9838 1690 9840
rect 1634 9786 1636 9838
rect 1636 9786 1688 9838
rect 1688 9786 1690 9838
rect 1634 9784 1690 9786
rect 916 9652 972 9654
rect 916 9600 918 9652
rect 918 9600 970 9652
rect 970 9600 972 9652
rect 916 9598 972 9600
rect 1439 9639 1495 9695
rect 294 9518 350 9520
rect 294 9466 296 9518
rect 296 9466 348 9518
rect 348 9466 350 9518
rect 294 9464 350 9466
rect 506 9518 562 9520
rect 506 9466 508 9518
rect 508 9466 560 9518
rect 560 9466 562 9518
rect 506 9464 562 9466
rect 1634 9652 1690 9654
rect 1634 9600 1636 9652
rect 1636 9600 1688 9652
rect 1688 9600 1690 9652
rect 1634 9598 1690 9600
rect 1439 9453 1495 9509
rect 601 9097 657 9099
rect 601 9045 603 9097
rect 603 9045 655 9097
rect 655 9045 657 9097
rect 601 9043 657 9045
rect 787 9097 843 9099
rect 787 9045 789 9097
rect 789 9045 841 9097
rect 841 9045 843 9097
rect 787 9043 843 9045
rect 1239 9080 1295 9082
rect 1239 9028 1241 9080
rect 1241 9028 1293 9080
rect 1293 9028 1295 9080
rect 1239 9026 1295 9028
rect 295 8981 351 8983
rect 295 8929 297 8981
rect 297 8929 349 8981
rect 349 8929 351 8981
rect 295 8927 351 8929
rect 295 8795 351 8797
rect 295 8743 297 8795
rect 297 8743 349 8795
rect 349 8743 351 8795
rect 295 8741 351 8743
rect 1239 8894 1295 8896
rect 1239 8842 1241 8894
rect 1241 8842 1293 8894
rect 1293 8842 1295 8894
rect 1239 8840 1295 8842
rect 1057 8731 1113 8733
rect 1057 8679 1059 8731
rect 1059 8679 1111 8731
rect 1111 8679 1113 8731
rect 1057 8677 1113 8679
rect 1057 8545 1113 8547
rect 1057 8493 1059 8545
rect 1059 8493 1111 8545
rect 1111 8493 1113 8545
rect 1057 8491 1113 8493
rect 1628 9080 1684 9082
rect 1628 9028 1630 9080
rect 1630 9028 1682 9080
rect 1682 9028 1684 9080
rect 1628 9026 1684 9028
rect 1628 8894 1684 8896
rect 1628 8842 1630 8894
rect 1630 8842 1682 8894
rect 1682 8842 1684 8894
rect 1628 8840 1684 8842
rect 2061 9080 2117 9082
rect 2061 9028 2063 9080
rect 2063 9028 2115 9080
rect 2115 9028 2117 9080
rect 2061 9026 2117 9028
rect 2061 8840 2117 8896
rect 2460 12568 2516 12624
rect 2460 12382 2516 12438
rect 2460 11793 2516 11849
rect 2460 11607 2516 11663
rect 2460 10877 2516 10933
rect 2460 10691 2516 10747
rect 2790 9933 2846 9935
rect 2790 9881 2792 9933
rect 2792 9881 2844 9933
rect 2844 9881 2846 9933
rect 2790 9879 2846 9881
rect 2790 9747 2846 9749
rect 2790 9695 2792 9747
rect 2792 9695 2844 9747
rect 2844 9695 2846 9747
rect 2790 9693 2846 9695
rect 2790 9010 2846 9012
rect 2790 8958 2792 9010
rect 2792 8958 2844 9010
rect 2844 8958 2846 9010
rect 2790 8956 2846 8958
rect 2790 8824 2846 8826
rect 2790 8772 2792 8824
rect 2792 8772 2844 8824
rect 2844 8772 2846 8824
rect 2790 8770 2846 8772
rect 2141 4933 2301 4989
<< metal3 >>
rect 322 28958 5618 29100
rect 322 28902 916 28958
rect 972 28902 1530 28958
rect 1586 28902 2155 28958
rect 2211 28902 2769 28958
rect 2825 28902 3393 28958
rect 3449 28902 4007 28958
rect 4063 28902 4632 28958
rect 4688 28902 5246 28958
rect 5302 28902 5618 28958
rect 322 28772 5618 28902
rect 322 28716 916 28772
rect 972 28716 1530 28772
rect 1586 28716 2155 28772
rect 2211 28716 2769 28772
rect 2825 28716 3393 28772
rect 3449 28716 4007 28772
rect 4063 28716 4632 28772
rect 4688 28716 5246 28772
rect 5302 28716 5618 28772
rect 322 27291 5618 28716
rect -269 24679 7633 24689
rect -269 24415 1223 24679
rect 1279 24415 2462 24679
rect 2518 24415 3700 24679
rect 3756 24415 4939 24679
rect 4995 24415 7633 24679
rect -269 24405 7633 24415
rect -1 22626 5603 23409
rect -1 22570 99 22626
rect 155 22570 492 22626
rect 548 22570 5603 22626
rect -1 22440 5603 22570
rect -1 22384 99 22440
rect 155 22384 492 22440
rect 548 22384 5603 22440
rect -1 22016 5603 22384
rect -1 22009 5325 22016
rect -1 21849 829 22009
rect 885 21849 1617 22009
rect 1673 21849 2068 22009
rect 2124 21849 2856 22009
rect 2912 21849 3306 22009
rect 3362 21849 4094 22009
rect 4150 21849 4545 22009
rect 4601 21856 5325 22009
rect 5381 21856 5603 22016
rect 4601 21849 5603 21856
rect -1 21410 5603 21849
rect 322 21179 5603 21299
rect 322 21123 5467 21179
rect 5523 21123 5603 21179
rect 322 21084 5603 21123
rect 322 20860 5603 20977
rect 322 20804 4412 20860
rect 4468 20804 5603 20860
rect 322 20762 5603 20804
rect 322 20531 5603 20656
rect 322 20475 4228 20531
rect 4284 20475 5603 20531
rect 322 20441 5603 20475
rect 4209 20436 4303 20441
rect 322 20218 5603 20334
rect 322 20162 3174 20218
rect 3230 20162 5603 20218
rect 322 20119 5603 20162
rect 322 19558 5603 19642
rect 322 19502 2989 19558
rect 3045 19502 5603 19558
rect 322 19427 5603 19502
rect 322 19246 5603 19320
rect 322 19190 1935 19246
rect 1991 19190 5603 19246
rect 322 19105 5603 19190
rect 322 18919 5603 18998
rect 322 18863 1751 18919
rect 1807 18863 5603 18919
rect 322 18783 5603 18863
rect 322 18604 5603 18676
rect 322 18548 697 18604
rect 753 18548 5603 18604
rect 322 18461 5603 18548
rect 322 18173 5603 18355
rect 322 18013 1697 18173
rect 1753 18013 1988 18173
rect 2044 18013 2936 18173
rect 2992 18013 3227 18173
rect 3283 18013 4174 18173
rect 4230 18013 4465 18173
rect 4521 18013 5603 18173
rect 322 17913 5603 18013
rect 322 16935 5603 17257
rect 322 16879 913 16935
rect 969 16879 1533 16935
rect 1589 16879 2152 16935
rect 2208 16879 2772 16935
rect 2828 16879 3390 16935
rect 3446 16879 4010 16935
rect 4066 16879 4629 16935
rect 4685 16879 5249 16935
rect 5305 16879 5603 16935
rect 322 16802 5603 16879
rect 368 16185 5517 16228
rect 368 16129 965 16185
rect 1021 16182 5517 16185
rect 1021 16129 1804 16182
rect 368 16126 1804 16129
rect 1860 16126 2015 16182
rect 2071 16126 2225 16182
rect 2281 16126 2436 16182
rect 2492 16126 2648 16182
rect 2704 16126 2859 16182
rect 2915 16126 3069 16182
rect 3125 16126 3280 16182
rect 3336 16126 3756 16182
rect 3812 16126 3967 16182
rect 4023 16126 4179 16182
rect 4235 16126 4390 16182
rect 4446 16126 5517 16182
rect 368 16000 5517 16126
rect 276 15607 2779 15713
rect 276 15551 295 15607
rect 351 15560 2779 15607
rect 351 15551 1655 15560
rect 276 15504 1655 15551
rect 1711 15504 1841 15560
rect 1897 15504 2779 15560
rect 276 15421 2779 15504
rect 276 15365 295 15421
rect 351 15365 2779 15421
rect 276 15142 2779 15365
rect 276 15086 1375 15142
rect 1431 15086 2779 15142
rect 276 15042 2779 15086
rect 276 15008 1865 15042
rect 276 14952 295 15008
rect 351 14986 1865 15008
rect 1921 14986 2779 15042
rect 351 14956 2779 14986
rect 351 14952 1375 14956
rect 276 14900 1375 14952
rect 1431 14900 2779 14956
rect 276 14856 2779 14900
rect 276 14822 1865 14856
rect 276 14766 295 14822
rect 351 14800 1865 14822
rect 1921 14800 2779 14856
rect 351 14766 2779 14800
rect 276 13551 2779 14766
rect 276 13495 295 13551
rect 351 13495 1865 13551
rect 1921 13495 2779 13551
rect 276 13365 2779 13495
rect 276 13309 295 13365
rect 351 13309 1865 13365
rect 1921 13309 2779 13365
rect 276 12991 2779 13309
rect 5493 12991 5794 15714
rect 276 12624 2779 12705
rect 276 12568 2091 12624
rect 2147 12568 2460 12624
rect 2516 12568 2779 12624
rect 276 12556 2779 12568
rect 276 12500 295 12556
rect 351 12500 1852 12556
rect 1908 12500 2779 12556
rect 276 12438 2779 12500
rect 276 12382 2091 12438
rect 2147 12382 2460 12438
rect 2516 12382 2779 12438
rect 276 12370 2779 12382
rect 276 12314 295 12370
rect 351 12314 1852 12370
rect 1908 12314 2779 12370
rect 276 11849 2779 12314
rect 276 11793 2091 11849
rect 2147 11793 2460 11849
rect 2516 11793 2779 11849
rect 276 11663 2779 11793
rect 276 11608 2091 11663
rect 276 11552 295 11608
rect 351 11552 1852 11608
rect 1908 11607 2091 11608
rect 2147 11607 2460 11663
rect 2516 11607 2779 11663
rect 1908 11552 2779 11607
rect 276 11422 2779 11552
rect 276 11366 295 11422
rect 351 11366 1852 11422
rect 1908 11366 2779 11422
rect 276 10933 2779 11366
rect 276 10877 2091 10933
rect 2147 10877 2460 10933
rect 2516 10877 2779 10933
rect 276 10747 2779 10877
rect 276 10692 2091 10747
rect 276 10636 295 10692
rect 351 10636 1852 10692
rect 1908 10691 2091 10692
rect 2147 10691 2460 10747
rect 2516 10691 2779 10747
rect 1908 10636 2779 10691
rect 276 10506 2779 10636
rect 276 10450 295 10506
rect 351 10450 1852 10506
rect 1908 10450 2779 10506
rect 276 9963 2779 10450
rect 276 9935 2865 9963
rect 276 9879 2790 9935
rect 2846 9879 2865 9935
rect 276 9840 2865 9879
rect 276 9784 916 9840
rect 972 9784 1634 9840
rect 1690 9784 2865 9840
rect 276 9749 2865 9784
rect 276 9695 2790 9749
rect 276 9654 1439 9695
rect 276 9598 916 9654
rect 972 9639 1439 9654
rect 1495 9693 2790 9695
rect 2846 9693 2865 9749
rect 1495 9654 2865 9693
rect 1495 9639 1634 9654
rect 972 9598 1634 9639
rect 1690 9598 2779 9654
rect 276 9559 2779 9598
rect 258 9520 2779 9559
rect 258 9464 294 9520
rect 350 9464 506 9520
rect 562 9509 2779 9520
rect 562 9464 1439 9509
rect 258 9453 1439 9464
rect 1495 9453 2779 9509
rect 258 9425 2779 9453
rect 276 9303 2779 9425
rect 276 9099 2779 9153
rect 276 9043 601 9099
rect 657 9043 787 9099
rect 843 9082 2779 9099
rect 843 9043 1239 9082
rect 276 9026 1239 9043
rect 1295 9026 1628 9082
rect 1684 9026 2061 9082
rect 2117 9040 2779 9082
rect 2117 9026 2865 9040
rect 276 9012 2865 9026
rect 276 8983 2790 9012
rect 276 8927 295 8983
rect 351 8956 2790 8983
rect 2846 8956 2865 9012
rect 351 8927 2865 8956
rect 276 8896 2865 8927
rect 276 8840 1239 8896
rect 1295 8840 1628 8896
rect 1684 8840 2061 8896
rect 2117 8840 2865 8896
rect 276 8826 2865 8840
rect 276 8797 2790 8826
rect 276 8741 295 8797
rect 351 8770 2790 8797
rect 2846 8770 2865 8826
rect 351 8741 2865 8770
rect 276 8733 2865 8741
rect 276 8677 1057 8733
rect 1113 8731 2865 8733
rect 1113 8677 2779 8731
rect 276 8547 2779 8677
rect 276 8491 1057 8547
rect 1113 8491 2779 8547
rect 276 8436 2779 8491
rect 318 4989 2311 5005
rect 318 4933 2141 4989
rect 2301 4933 2311 4989
rect 318 4917 2311 4933
rect 5627 3128 5794 4490
rect 5636 149 5794 604
use din_256x8m81  din_256x8m81_0
timestamp 1749760379
transform 1 0 323 0 1 7805
box -46 -15 2450 8740
use M2_M1$$45012012_256x8m81  M2_M1$$45012012_256x8m81_0
timestamp 1749760379
transform 1 0 2570 0 1 16154
box 0 0 1 1
use M2_M1$$45013036_256x8m81  M2_M1$$45013036_256x8m81_0
timestamp 1749760379
transform 1 0 4101 0 1 16154
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_0
timestamp 1749760379
transform 0 -1 5163 1 0 5513
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_1
timestamp 1749760379
transform 0 -1 4677 1 0 5513
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_2
timestamp 1749760379
transform 1 0 956 0 1 -127
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_0
timestamp 1749760379
transform 1 0 3038 0 1 -2344
box 0 0 1 1
use m2_saout01_256x8m81  m2_saout01_256x8m81_0
timestamp 1749760379
transform 1 0 686 0 1 28980
box -89 -63 4849 2153
use M3_M2$$43370540_256x8m81  M3_M2$$43370540_256x8m81_0
timestamp 1749760379
transform 1 0 4101 0 1 16154
box 0 0 1 1
use M3_M2$$44741676_256x8m81  M3_M2$$44741676_256x8m81_0
timestamp 1749760379
transform 1 0 2570 0 1 16154
box 0 0 1 1
use M3_M2431059087814_256x8m81  M3_M2431059087814_256x8m81_0
timestamp 1749760379
transform 1 0 2221 0 1 4961
box 0 0 1 1
use mux821_256x8m81  mux821_256x8m81_0
timestamp 1749760379
transform 1 0 553 0 1 16662
box -9 164 5035 12234
use outbuf_oe_256x8m81  outbuf_oe_256x8m81_0
timestamp 1749760379
transform 1 0 632 0 1 5509
box -532 -359 5177 3324
use sa_256x8m81  sa_256x8m81_0
timestamp 1749760379
transform 1 0 632 0 1 8608
box -357 -196 5034 8146
use sacntl_2_256x8m81  sacntl_2_256x8m81_0
timestamp 1749760379
transform 1 0 632 0 1 23
box -530 -24 5176 5655
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_0
timestamp 1749760379
transform 1 0 2073 0 1 12344
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_1
timestamp 1749760379
transform 1 0 2073 0 1 11569
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_2
timestamp 1749760379
transform 1 0 2073 0 1 10653
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_0
timestamp 1749760379
transform 0 1 5389 1 0 18308
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_1
timestamp 1749760379
transform 0 -1 628 1 0 15874
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_2
timestamp 1749760379
transform 0 -1 540 1 0 27025
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_3
timestamp 1749760379
transform 0 -1 826 1 0 18308
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_0
timestamp 1749760379
transform -1 0 2350 0 -1 15969
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_1
timestamp 1749760379
transform -1 0 1577 0 -1 6674
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_2
timestamp 1749760379
transform 1 0 2257 0 1 3326
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_3
timestamp 1749760379
transform 1 0 5345 0 1 9961
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_4
timestamp 1749760379
transform 1 0 461 0 1 8245
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_0
timestamp 1749760379
transform 0 -1 5132 1 0 16336
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_1
timestamp 1749760379
transform 0 -1 2025 1 0 18308
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_2
timestamp 1749760379
transform 0 -1 3263 1 0 18308
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_3
timestamp 1749760379
transform 0 -1 4502 1 0 18308
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_4
timestamp 1749760379
transform 0 -1 925 1 0 8791
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_0
timestamp 1749760379
transform -1 0 771 0 1 18510
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_1
timestamp 1749760379
transform -1 0 1825 0 1 18825
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_2
timestamp 1749760379
transform -1 0 2009 0 1 19152
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_3
timestamp 1749760379
transform -1 0 4302 0 1 20437
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_4
timestamp 1749760379
transform -1 0 4486 0 1 20766
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_5
timestamp 1749760379
transform -1 0 5541 0 1 21085
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_6
timestamp 1749760379
transform 1 0 2971 0 1 19464
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_7
timestamp 1749760379
transform 1 0 3156 0 1 20124
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_0
timestamp 1749760379
transform 1 0 474 0 1 22346
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_1
timestamp 1749760379
transform 1 0 81 0 1 22346
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_2
timestamp 1749760379
transform 1 0 2442 0 1 12344
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_3
timestamp 1749760379
transform 1 0 2442 0 1 11569
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_4
timestamp 1749760379
transform 1 0 2442 0 1 10653
box 0 0 1 1
use wen_wm1_256x8m81  wen_wm1_256x8m81_0
timestamp 1749760379
transform 1 0 322 0 1 -3376
box -156 -24 4946 3287
<< labels >>
rlabel metal1 s 993 27075 993 27075 4 pcb
port 1 nsew
rlabel metal1 s 698 8313 698 8313 4 datain
port 2 nsew
rlabel metal1 s 993 27073 993 27073 4 pcb
port 1 nsew
rlabel metal1 s 933 18156 933 18156 4 vdd
port 3 nsew
flabel metal1 s 709 -3344 709 -3344 0 FreeSans 600 0 0 0 WEN
port 4 nsew
rlabel metal3 s 810 18907 810 18907 4 ypass[1]
port 5 nsew
rlabel metal3 s 810 19224 810 19224 4 ypass[2]
port 6 nsew
rlabel metal3 s 810 19542 810 19542 4 ypass[3]
port 7 nsew
rlabel metal3 s 810 20197 810 20197 4 ypass[4]
port 8 nsew
rlabel metal3 s 810 20521 810 20521 4 ypass[5]
port 9 nsew
rlabel metal3 s 810 20838 810 20838 4 ypass[6]
port 10 nsew
rlabel metal3 s 810 21156 810 21156 4 ypass[7]
port 11 nsew
rlabel metal3 s 881 1460 881 1460 4 men
port 12 nsew
rlabel metal3 s 373 1086 373 1086 4 vss
port 13 nsew
rlabel metal3 s 440 2179 440 2179 4 vss
port 13 nsew
rlabel metal3 s 810 20197 810 20197 4 ypass[4]
port 8 nsew
rlabel metal3 s 545 3843 545 3843 4 vdd
port 3 nsew
rlabel metal3 s 393 399 393 399 4 vdd
port 3 nsew
rlabel metal3 s 454 6155 454 6155 4 vss
port 13 nsew
rlabel metal3 s 439 11029 439 11029 4 vss
port 13 nsew
rlabel metal3 s 810 21156 810 21156 4 ypass[7]
port 11 nsew
rlabel metal3 s 810 20838 810 20838 4 ypass[6]
port 10 nsew
rlabel metal3 s 810 20521 810 20521 4 ypass[5]
port 9 nsew
rlabel metal3 s 810 19542 810 19542 4 ypass[3]
port 7 nsew
rlabel metal3 s 810 19224 810 19224 4 ypass[2]
port 6 nsew
rlabel metal3 s 810 18907 810 18907 4 ypass[1]
port 5 nsew
rlabel metal3 s 810 18585 810 18585 4 ypass[0]
port 14 nsew
rlabel metal3 s 398 1458 398 1458 4 men
port 12 nsew
rlabel metal3 s 933 28895 933 28895 4 vdd
port 3 nsew
rlabel metal3 s 949 22008 949 22008 4 vss
port 13 nsew
rlabel metal3 s 477 17166 477 17166 4 vss
port 13 nsew
rlabel metal3 s 466 13763 466 13763 4 vdd
port 3 nsew
rlabel metal3 s 401 8726 401 8726 4 vdd
port 3 nsew
rlabel metal3 s 335 7368 335 7368 4 vdd
port 3 nsew
rlabel metal3 s 810 18585 810 18585 4 ypass[0]
port 14 nsew
flabel metal3 s 644 4959 644 4959 0 FreeSans 600 0 0 0 GWE
port 15 nsew
rlabel metal3 s 393 -592 393 -592 4 vdd
port 3 nsew
rlabel metal3 s 373 -1762 373 -1762 4 vss
port 13 nsew
rlabel metal3 s 373 -2331 373 -2331 4 vss
port 13 nsew
rlabel metal3 s 393 -2997 393 -2997 4 vdd
port 3 nsew
rlabel metal3 s 373 -1375 373 -1375 4 vss
port 13 nsew
flabel metal3 s 705 -2005 705 -2005 0 FreeSans 600 0 0 0 GWEN
port 16 nsew
rlabel metal2 s 501 1625 501 1625 4 datain
port 2 nsew
rlabel metal2 s 5501 28725 5501 28725 4 b[7]
port 17 nsew
rlabel metal2 s 4464 28725 4464 28725 4 b[6]
port 18 nsew
rlabel metal2 s 4256 28725 4256 28725 4 b[5]
port 19 nsew
rlabel metal2 s 3228 28725 3228 28725 4 b[4]
port 20 nsew
rlabel metal2 s 3024 28725 3024 28725 4 b[3]
port 21 nsew
rlabel metal2 s 1983 28725 1983 28725 4 b[2]
port 22 nsew
rlabel metal2 s 1781 28725 1781 28725 4 b[1]
port 23 nsew
rlabel metal2 s 736 28727 736 28727 4 b[0]
port 24 nsew
rlabel metal2 s 4880 28727 4880 28727 4 bb[6]
port 25 nsew
rlabel metal2 s 5082 28734 5082 28734 4 bb[7]
port 26 nsew
rlabel metal2 s 3841 28727 3841 28727 4 bb[5]
port 27 nsew
rlabel metal2 s 1351 1158 1351 1158 4 q
port 28 nsew
rlabel metal2 s 3641 28727 3641 28727 4 bb[4]
port 29 nsew
rlabel metal2 s 2604 28734 2604 28734 4 bb[3]
port 30 nsew
rlabel metal2 s 2405 28730 2405 28730 4 bb[2]
port 31 nsew
rlabel metal2 s 1162 28725 1162 28725 4 bb[0]
port 32 nsew
rlabel metal2 s 1368 28725 1368 28725 4 bb[1]
port 33 nsew
rlabel metal2 s 1351 1124 1351 1124 4 q
port 28 nsew
<< properties >>
string GDS_END 819092
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 810738
string path 10.130 4.930 10.130 -9.675 15.190 -9.675 15.190 -12.125 
<< end >>
