magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 453 3894 1094
<< pwell >>
rect -86 -86 3894 453
<< metal1 >>
rect 0 918 3808 1098
rect 49 710 95 918
rect 273 664 319 872
rect 477 710 523 918
rect 701 664 747 872
rect 925 710 971 918
rect 1149 664 1195 872
rect 1373 710 1419 918
rect 1597 664 1643 872
rect 1821 710 1867 918
rect 2045 664 2091 872
rect 2269 710 2315 918
rect 2493 664 2539 872
rect 2717 710 2763 918
rect 2941 664 2987 872
rect 3165 710 3211 918
rect 3389 664 3435 872
rect 3613 710 3659 918
rect 273 618 3435 664
rect 126 454 1604 530
rect 1653 349 1813 618
rect 1859 454 3337 530
rect 273 303 3455 349
rect 49 90 95 257
rect 273 189 325 303
rect 497 90 543 257
rect 721 189 767 303
rect 945 90 991 257
rect 1169 189 1215 303
rect 1393 90 1439 257
rect 1617 189 1663 303
rect 1841 90 1887 257
rect 2065 189 2111 303
rect 2289 90 2335 257
rect 2513 189 2559 303
rect 2737 90 2783 257
rect 2961 189 3007 303
rect 3185 90 3231 257
rect 3409 189 3455 303
rect 3633 90 3679 257
rect 0 -90 3808 90
<< labels >>
rlabel metal1 s 1859 454 3337 530 6 I
port 1 nsew default input
rlabel metal1 s 126 454 1604 530 6 I
port 1 nsew default input
rlabel metal1 s 3409 189 3455 303 6 ZN
port 2 nsew default output
rlabel metal1 s 2961 189 3007 303 6 ZN
port 2 nsew default output
rlabel metal1 s 2513 189 2559 303 6 ZN
port 2 nsew default output
rlabel metal1 s 2065 189 2111 303 6 ZN
port 2 nsew default output
rlabel metal1 s 1617 189 1663 303 6 ZN
port 2 nsew default output
rlabel metal1 s 1169 189 1215 303 6 ZN
port 2 nsew default output
rlabel metal1 s 721 189 767 303 6 ZN
port 2 nsew default output
rlabel metal1 s 273 189 325 303 6 ZN
port 2 nsew default output
rlabel metal1 s 273 303 3455 349 6 ZN
port 2 nsew default output
rlabel metal1 s 1653 349 1813 618 6 ZN
port 2 nsew default output
rlabel metal1 s 273 618 3435 664 6 ZN
port 2 nsew default output
rlabel metal1 s 3389 664 3435 872 6 ZN
port 2 nsew default output
rlabel metal1 s 2941 664 2987 872 6 ZN
port 2 nsew default output
rlabel metal1 s 2493 664 2539 872 6 ZN
port 2 nsew default output
rlabel metal1 s 2045 664 2091 872 6 ZN
port 2 nsew default output
rlabel metal1 s 1597 664 1643 872 6 ZN
port 2 nsew default output
rlabel metal1 s 1149 664 1195 872 6 ZN
port 2 nsew default output
rlabel metal1 s 701 664 747 872 6 ZN
port 2 nsew default output
rlabel metal1 s 273 664 319 872 6 ZN
port 2 nsew default output
rlabel metal1 s 3613 710 3659 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 710 3211 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 710 2763 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 710 2315 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 710 1867 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 710 1419 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 710 971 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 710 523 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 918 3808 1098 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 453 3894 1094 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 3894 453 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -90 3808 90 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3633 90 3679 257 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3185 90 3231 257 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2737 90 2783 257 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2289 90 2335 257 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1841 90 1887 257 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1393 90 1439 257 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 257 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 257 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 257 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1474654
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1465608
<< end >>
