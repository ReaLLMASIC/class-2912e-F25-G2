magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 352 2774 870
<< pwell >>
rect -86 -86 2774 352
<< mvnmos >>
rect 124 79 244 172
rect 384 93 504 172
rect 552 93 672 172
rect 720 93 840 172
rect 944 93 1064 172
rect 1112 93 1232 172
rect 1280 93 1400 172
rect 1540 93 1660 186
rect 1760 93 1880 186
rect 2132 139 2252 232
rect 2392 68 2512 232
<< mvpmos >>
rect 124 531 224 716
rect 476 590 576 716
rect 680 590 780 716
rect 828 590 928 716
rect 1032 590 1132 716
rect 1192 590 1292 716
rect 1540 590 1640 716
rect 1780 531 1880 716
rect 2132 531 2232 716
rect 2412 472 2512 716
<< mvndiff >>
rect 2044 204 2132 232
rect 1460 172 1540 186
rect 36 152 124 172
rect 36 106 49 152
rect 95 106 124 152
rect 36 79 124 106
rect 244 152 384 172
rect 244 106 273 152
rect 319 106 384 152
rect 244 93 384 106
rect 504 93 552 172
rect 672 93 720 172
rect 840 152 944 172
rect 840 106 869 152
rect 915 106 944 152
rect 840 93 944 106
rect 1064 93 1112 172
rect 1232 93 1280 172
rect 1400 158 1540 172
rect 1400 112 1465 158
rect 1511 112 1540 158
rect 1400 93 1540 112
rect 1660 93 1760 186
rect 1880 167 1968 186
rect 1880 121 1909 167
rect 1955 121 1968 167
rect 2044 158 2057 204
rect 2103 158 2132 204
rect 2044 139 2132 158
rect 2252 204 2392 232
rect 2252 158 2281 204
rect 2327 158 2392 204
rect 2252 139 2392 158
rect 1880 93 1968 121
rect 244 79 324 93
rect 2312 68 2392 139
rect 2512 204 2600 232
rect 2512 158 2541 204
rect 2587 158 2600 204
rect 2512 68 2600 158
<< mvpdiff >>
rect 36 651 124 716
rect 36 605 49 651
rect 95 605 124 651
rect 36 531 124 605
rect 224 703 312 716
rect 224 563 253 703
rect 299 563 312 703
rect 388 667 476 716
rect 388 621 401 667
rect 447 621 476 667
rect 388 590 476 621
rect 576 703 680 716
rect 576 657 605 703
rect 651 657 680 703
rect 576 590 680 657
rect 780 590 828 716
rect 928 667 1032 716
rect 928 621 957 667
rect 1003 621 1032 667
rect 928 590 1032 621
rect 1132 590 1192 716
rect 1292 703 1540 716
rect 1292 657 1403 703
rect 1449 657 1540 703
rect 1292 590 1540 657
rect 1640 667 1780 716
rect 1640 621 1705 667
rect 1751 621 1780 667
rect 1640 590 1780 621
rect 224 531 312 563
rect 1700 531 1780 590
rect 1880 703 1968 716
rect 1880 563 1909 703
rect 1955 563 1968 703
rect 1880 531 1968 563
rect 2044 639 2132 716
rect 2044 593 2057 639
rect 2103 593 2132 639
rect 2044 531 2132 593
rect 2232 703 2412 716
rect 2232 563 2337 703
rect 2383 563 2412 703
rect 2232 531 2412 563
rect 2312 472 2412 531
rect 2512 665 2600 716
rect 2512 525 2541 665
rect 2587 525 2600 665
rect 2512 472 2600 525
<< mvndiffc >>
rect 49 106 95 152
rect 273 106 319 152
rect 869 106 915 152
rect 1465 112 1511 158
rect 1909 121 1955 167
rect 2057 158 2103 204
rect 2281 158 2327 204
rect 2541 158 2587 204
<< mvpdiffc >>
rect 49 605 95 651
rect 253 563 299 703
rect 401 621 447 667
rect 605 657 651 703
rect 957 621 1003 667
rect 1403 657 1449 703
rect 1705 621 1751 667
rect 1909 563 1955 703
rect 2057 593 2103 639
rect 2337 563 2383 703
rect 2541 525 2587 665
<< polysilicon >>
rect 124 716 224 760
rect 476 716 576 760
rect 680 716 780 760
rect 828 716 928 760
rect 1032 716 1132 760
rect 1192 716 1292 760
rect 1540 716 1640 760
rect 1780 716 1880 760
rect 2132 716 2232 760
rect 2412 716 2512 760
rect 124 340 224 531
rect 476 519 576 590
rect 476 504 503 519
rect 384 473 503 504
rect 549 473 576 519
rect 384 454 576 473
rect 124 255 244 340
rect 124 209 163 255
rect 209 209 244 255
rect 124 172 244 209
rect 384 172 504 454
rect 680 406 780 590
rect 552 366 780 406
rect 828 427 928 590
rect 828 381 855 427
rect 901 423 928 427
rect 901 381 984 423
rect 828 368 984 381
rect 552 312 672 366
rect 552 266 592 312
rect 638 266 672 312
rect 552 172 672 266
rect 720 253 840 266
rect 720 207 755 253
rect 801 207 840 253
rect 720 172 840 207
rect 944 260 984 368
rect 1032 408 1132 590
rect 1032 362 1045 408
rect 1091 362 1132 408
rect 1032 349 1132 362
rect 1192 496 1292 590
rect 1192 450 1233 496
rect 1279 450 1292 496
rect 1192 437 1292 450
rect 1540 496 1640 590
rect 1540 450 1566 496
rect 1612 450 1640 496
rect 1540 440 1640 450
rect 1780 440 1880 531
rect 1192 260 1232 437
rect 944 172 1064 260
rect 1112 172 1232 260
rect 1280 359 1400 372
rect 1280 313 1317 359
rect 1363 313 1400 359
rect 1280 172 1400 313
rect 1540 267 1660 440
rect 1540 221 1566 267
rect 1612 221 1660 267
rect 1540 186 1660 221
rect 1760 404 1880 440
rect 1760 358 1815 404
rect 1861 358 1880 404
rect 1760 186 1880 358
rect 2132 435 2232 531
rect 2132 404 2252 435
rect 2132 358 2168 404
rect 2214 358 2252 404
rect 2412 404 2512 472
rect 2412 394 2429 404
rect 2132 232 2252 358
rect 2392 358 2429 394
rect 2475 358 2512 404
rect 2392 232 2512 358
rect 124 24 244 79
rect 384 24 504 93
rect 552 24 672 93
rect 720 24 840 93
rect 944 24 1064 93
rect 1112 24 1232 93
rect 1280 24 1400 93
rect 1540 24 1660 93
rect 1760 24 1880 93
rect 2132 24 2252 139
rect 2392 24 2512 68
<< polycontact >>
rect 503 473 549 519
rect 163 209 209 255
rect 855 381 901 427
rect 592 266 638 312
rect 755 207 801 253
rect 1045 362 1091 408
rect 1233 450 1279 496
rect 1566 450 1612 496
rect 1317 313 1363 359
rect 1566 221 1612 267
rect 1815 358 1861 404
rect 2168 358 2214 404
rect 2429 358 2475 404
<< metal1 >>
rect 0 724 2688 844
rect 253 703 299 724
rect 38 651 95 662
rect 38 605 49 651
rect 38 427 95 605
rect 594 703 662 724
rect 401 667 447 678
rect 594 657 605 703
rect 651 657 662 703
rect 1392 703 1460 724
rect 401 611 447 621
rect 712 621 957 667
rect 1003 621 1289 667
rect 1392 657 1403 703
rect 1449 657 1460 703
rect 1909 703 1955 724
rect 1705 667 1751 678
rect 712 611 758 621
rect 401 565 758 611
rect 1239 611 1289 621
rect 1239 565 1623 611
rect 253 531 299 563
rect 800 519 1187 536
rect 476 473 503 519
rect 549 473 1187 519
rect 38 381 855 427
rect 901 381 928 427
rect 1032 408 1095 427
rect 38 152 106 381
rect 1032 362 1045 408
rect 1091 362 1095 408
rect 457 312 662 326
rect 457 266 592 312
rect 638 266 662 312
rect 152 209 163 255
rect 209 209 411 255
rect 457 248 662 266
rect 1032 253 1095 362
rect 1141 359 1187 473
rect 1233 496 1509 507
rect 1279 450 1509 496
rect 1555 496 1623 565
rect 1555 450 1566 496
rect 1612 450 1623 496
rect 1233 439 1509 450
rect 1463 404 1509 439
rect 1705 404 1751 621
rect 2326 703 2394 724
rect 1909 531 1955 563
rect 2057 639 2103 650
rect 2057 514 2103 593
rect 2326 563 2337 703
rect 2383 563 2394 703
rect 2530 665 2662 676
rect 2530 525 2541 665
rect 2587 525 2662 665
rect 1141 313 1317 359
rect 1363 313 1400 359
rect 1463 358 1751 404
rect 365 200 411 209
rect 735 207 755 253
rect 801 207 1095 253
rect 1373 221 1566 267
rect 1612 221 1623 267
rect 735 200 781 207
rect 38 106 49 152
rect 95 106 106 152
rect 273 152 319 163
rect 365 136 781 200
rect 1373 152 1419 221
rect 858 106 869 152
rect 915 106 1419 152
rect 1465 158 1511 175
rect 1705 167 1751 358
rect 1802 404 1880 471
rect 2057 468 2339 514
rect 2530 506 2662 525
rect 2293 404 2339 468
rect 1802 358 1815 404
rect 1861 358 1880 404
rect 1802 217 1880 358
rect 1952 358 2168 404
rect 2214 358 2225 404
rect 2293 358 2429 404
rect 2475 358 2486 404
rect 1952 167 1998 358
rect 2293 307 2339 358
rect 1705 121 1909 167
rect 1955 121 1998 167
rect 2057 261 2339 307
rect 2057 204 2103 261
rect 2600 224 2662 506
rect 2057 147 2103 158
rect 2281 204 2327 215
rect 273 60 319 106
rect 1465 60 1511 112
rect 2281 60 2327 158
rect 2486 204 2662 224
rect 2486 158 2541 204
rect 2587 158 2662 204
rect 2486 120 2662 158
rect 0 -60 2688 60
<< labels >>
flabel metal1 s 1802 217 1880 471 0 FreeSans 400 0 0 0 SETN
port 4 nsew default input
flabel metal1 s 2530 506 2662 676 0 FreeSans 400 0 0 0 Q
port 5 nsew default output
flabel metal1 s 800 519 1187 536 0 FreeSans 400 0 0 0 RN
port 3 nsew default input
flabel metal1 s 2281 175 2327 215 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 1032 255 1095 427 0 FreeSans 400 0 0 0 E
port 2 nsew clock input
flabel metal1 s 0 724 2688 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 457 248 662 326 0 FreeSans 400 0 0 0 D
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 1032 253 1095 255 1 E
port 2 nsew clock input
rlabel metal1 s 152 253 411 255 1 E
port 2 nsew clock input
rlabel metal1 s 735 209 1095 253 1 E
port 2 nsew clock input
rlabel metal1 s 152 209 411 253 1 E
port 2 nsew clock input
rlabel metal1 s 735 207 1095 209 1 E
port 2 nsew clock input
rlabel metal1 s 365 207 411 209 1 E
port 2 nsew clock input
rlabel metal1 s 735 200 781 207 1 E
port 2 nsew clock input
rlabel metal1 s 365 200 411 207 1 E
port 2 nsew clock input
rlabel metal1 s 365 136 781 200 1 E
port 2 nsew clock input
rlabel metal1 s 476 473 1187 519 1 RN
port 3 nsew default input
rlabel metal1 s 1141 359 1187 473 1 RN
port 3 nsew default input
rlabel metal1 s 1141 313 1400 359 1 RN
port 3 nsew default input
rlabel metal1 s 2600 224 2662 506 1 Q
port 5 nsew default output
rlabel metal1 s 2486 120 2662 224 1 Q
port 5 nsew default output
rlabel metal1 s 2326 657 2394 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1909 657 1955 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1392 657 1460 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 594 657 662 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 657 299 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2326 563 2394 657 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1909 563 1955 657 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 563 299 657 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1909 531 1955 563 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 531 299 563 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2281 163 2327 175 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1465 163 1511 175 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2281 60 2327 163 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1465 60 1511 163 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 163 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2688 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2688 784
string GDS_END 625276
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 618684
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
