magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< metal1 >>
rect 742 2131 1686 2143
rect 742 2079 754 2131
rect 806 2079 878 2131
rect 930 2079 1002 2131
rect 1054 2079 1126 2131
rect 1178 2079 1250 2131
rect 1302 2079 1374 2131
rect 1426 2079 1498 2131
rect 1550 2079 1622 2131
rect 1674 2079 1686 2131
rect 742 2007 1686 2079
rect 742 1955 754 2007
rect 806 1955 878 2007
rect 930 1955 1002 2007
rect 1054 1955 1126 2007
rect 1178 1955 1250 2007
rect 1302 1955 1374 2007
rect 1426 1955 1498 2007
rect 1550 1955 1622 2007
rect 1674 1955 1686 2007
rect 742 1883 1686 1955
rect 742 1831 754 1883
rect 806 1831 878 1883
rect 930 1831 1002 1883
rect 1054 1831 1126 1883
rect 1178 1831 1250 1883
rect 1302 1831 1374 1883
rect 1426 1831 1498 1883
rect 1550 1831 1622 1883
rect 1674 1831 1686 1883
rect 742 1819 1686 1831
rect 148 75 312 1728
<< via1 >>
rect 754 2079 806 2131
rect 878 2079 930 2131
rect 1002 2079 1054 2131
rect 1126 2079 1178 2131
rect 1250 2079 1302 2131
rect 1374 2079 1426 2131
rect 1498 2079 1550 2131
rect 1622 2079 1674 2131
rect 754 1955 806 2007
rect 878 1955 930 2007
rect 1002 1955 1054 2007
rect 1126 1955 1178 2007
rect 1250 1955 1302 2007
rect 1374 1955 1426 2007
rect 1498 1955 1550 2007
rect 1622 1955 1674 2007
rect 754 1831 806 1883
rect 878 1831 930 1883
rect 1002 1831 1054 1883
rect 1126 1831 1178 1883
rect 1250 1831 1302 1883
rect 1374 1831 1426 1883
rect 1498 1831 1550 1883
rect 1622 1831 1674 1883
<< metal2 >>
rect 742 2133 1686 2143
rect 742 2077 752 2133
rect 808 2077 876 2133
rect 932 2077 1000 2133
rect 1056 2077 1124 2133
rect 1180 2077 1248 2133
rect 1304 2077 1372 2133
rect 1428 2077 1496 2133
rect 1552 2077 1620 2133
rect 1676 2077 1686 2133
rect 742 2009 1686 2077
rect 742 1953 752 2009
rect 808 1953 876 2009
rect 932 1953 1000 2009
rect 1056 1953 1124 2009
rect 1180 1953 1248 2009
rect 1304 1953 1372 2009
rect 1428 1953 1496 2009
rect 1552 1953 1620 2009
rect 1676 1953 1686 2009
rect 742 1885 1686 1953
rect 742 1829 752 1885
rect 808 1829 876 1885
rect 932 1829 1000 1885
rect 1056 1829 1124 1885
rect 1180 1829 1248 1885
rect 1304 1829 1372 1885
rect 1428 1829 1496 1885
rect 1552 1829 1620 1885
rect 1676 1829 1686 1885
rect 742 1819 1686 1829
rect -484 1588 460 1598
rect -484 1532 -474 1588
rect -418 1532 -350 1588
rect -294 1532 -226 1588
rect -170 1532 -102 1588
rect -46 1532 22 1588
rect 78 1532 146 1588
rect 202 1532 270 1588
rect 326 1532 394 1588
rect 450 1532 460 1588
rect -484 1464 460 1532
rect -484 1408 -474 1464
rect -418 1408 -350 1464
rect -294 1408 -226 1464
rect -170 1408 -102 1464
rect -46 1408 22 1464
rect 78 1408 146 1464
rect 202 1408 270 1464
rect 326 1408 394 1464
rect 450 1408 460 1464
rect -484 1340 460 1408
rect -484 1284 -474 1340
rect -418 1284 -350 1340
rect -294 1284 -226 1340
rect -170 1284 -102 1340
rect -46 1284 22 1340
rect 78 1284 146 1340
rect 202 1284 270 1340
rect 326 1284 394 1340
rect 450 1284 460 1340
rect -484 1216 460 1284
rect -484 1160 -474 1216
rect -418 1160 -350 1216
rect -294 1160 -226 1216
rect -170 1160 -102 1216
rect -46 1160 22 1216
rect 78 1160 146 1216
rect 202 1160 270 1216
rect 326 1160 394 1216
rect 450 1160 460 1216
rect -484 1092 460 1160
rect -484 1036 -474 1092
rect -418 1036 -350 1092
rect -294 1036 -226 1092
rect -170 1036 -102 1092
rect -46 1036 22 1092
rect 78 1036 146 1092
rect 202 1036 270 1092
rect 326 1036 394 1092
rect 450 1036 460 1092
rect -484 968 460 1036
rect -484 912 -474 968
rect -418 912 -350 968
rect -294 912 -226 968
rect -170 912 -102 968
rect -46 912 22 968
rect 78 912 146 968
rect 202 912 270 968
rect 326 912 394 968
rect 450 912 460 968
rect -484 844 460 912
rect -484 788 -474 844
rect -418 788 -350 844
rect -294 788 -226 844
rect -170 788 -102 844
rect -46 788 22 844
rect 78 788 146 844
rect 202 788 270 844
rect 326 788 394 844
rect 450 788 460 844
rect -484 720 460 788
rect -484 664 -474 720
rect -418 664 -350 720
rect -294 664 -226 720
rect -170 664 -102 720
rect -46 664 22 720
rect 78 664 146 720
rect 202 664 270 720
rect 326 664 394 720
rect 450 664 460 720
rect -484 654 460 664
rect 360 0 460 654
<< via2 >>
rect 752 2131 808 2133
rect 752 2079 754 2131
rect 754 2079 806 2131
rect 806 2079 808 2131
rect 752 2077 808 2079
rect 876 2131 932 2133
rect 876 2079 878 2131
rect 878 2079 930 2131
rect 930 2079 932 2131
rect 876 2077 932 2079
rect 1000 2131 1056 2133
rect 1000 2079 1002 2131
rect 1002 2079 1054 2131
rect 1054 2079 1056 2131
rect 1000 2077 1056 2079
rect 1124 2131 1180 2133
rect 1124 2079 1126 2131
rect 1126 2079 1178 2131
rect 1178 2079 1180 2131
rect 1124 2077 1180 2079
rect 1248 2131 1304 2133
rect 1248 2079 1250 2131
rect 1250 2079 1302 2131
rect 1302 2079 1304 2131
rect 1248 2077 1304 2079
rect 1372 2131 1428 2133
rect 1372 2079 1374 2131
rect 1374 2079 1426 2131
rect 1426 2079 1428 2131
rect 1372 2077 1428 2079
rect 1496 2131 1552 2133
rect 1496 2079 1498 2131
rect 1498 2079 1550 2131
rect 1550 2079 1552 2131
rect 1496 2077 1552 2079
rect 1620 2131 1676 2133
rect 1620 2079 1622 2131
rect 1622 2079 1674 2131
rect 1674 2079 1676 2131
rect 1620 2077 1676 2079
rect 752 2007 808 2009
rect 752 1955 754 2007
rect 754 1955 806 2007
rect 806 1955 808 2007
rect 752 1953 808 1955
rect 876 2007 932 2009
rect 876 1955 878 2007
rect 878 1955 930 2007
rect 930 1955 932 2007
rect 876 1953 932 1955
rect 1000 2007 1056 2009
rect 1000 1955 1002 2007
rect 1002 1955 1054 2007
rect 1054 1955 1056 2007
rect 1000 1953 1056 1955
rect 1124 2007 1180 2009
rect 1124 1955 1126 2007
rect 1126 1955 1178 2007
rect 1178 1955 1180 2007
rect 1124 1953 1180 1955
rect 1248 2007 1304 2009
rect 1248 1955 1250 2007
rect 1250 1955 1302 2007
rect 1302 1955 1304 2007
rect 1248 1953 1304 1955
rect 1372 2007 1428 2009
rect 1372 1955 1374 2007
rect 1374 1955 1426 2007
rect 1426 1955 1428 2007
rect 1372 1953 1428 1955
rect 1496 2007 1552 2009
rect 1496 1955 1498 2007
rect 1498 1955 1550 2007
rect 1550 1955 1552 2007
rect 1496 1953 1552 1955
rect 1620 2007 1676 2009
rect 1620 1955 1622 2007
rect 1622 1955 1674 2007
rect 1674 1955 1676 2007
rect 1620 1953 1676 1955
rect 752 1883 808 1885
rect 752 1831 754 1883
rect 754 1831 806 1883
rect 806 1831 808 1883
rect 752 1829 808 1831
rect 876 1883 932 1885
rect 876 1831 878 1883
rect 878 1831 930 1883
rect 930 1831 932 1883
rect 876 1829 932 1831
rect 1000 1883 1056 1885
rect 1000 1831 1002 1883
rect 1002 1831 1054 1883
rect 1054 1831 1056 1883
rect 1000 1829 1056 1831
rect 1124 1883 1180 1885
rect 1124 1831 1126 1883
rect 1126 1831 1178 1883
rect 1178 1831 1180 1883
rect 1124 1829 1180 1831
rect 1248 1883 1304 1885
rect 1248 1831 1250 1883
rect 1250 1831 1302 1883
rect 1302 1831 1304 1883
rect 1248 1829 1304 1831
rect 1372 1883 1428 1885
rect 1372 1831 1374 1883
rect 1374 1831 1426 1883
rect 1426 1831 1428 1883
rect 1372 1829 1428 1831
rect 1496 1883 1552 1885
rect 1496 1831 1498 1883
rect 1498 1831 1550 1883
rect 1550 1831 1552 1883
rect 1496 1829 1552 1831
rect 1620 1883 1676 1885
rect 1620 1831 1622 1883
rect 1622 1831 1674 1883
rect 1674 1831 1676 1883
rect 1620 1829 1676 1831
rect -474 1532 -418 1588
rect -350 1532 -294 1588
rect -226 1532 -170 1588
rect -102 1532 -46 1588
rect 22 1532 78 1588
rect 146 1532 202 1588
rect 270 1532 326 1588
rect 394 1532 450 1588
rect -474 1408 -418 1464
rect -350 1408 -294 1464
rect -226 1408 -170 1464
rect -102 1408 -46 1464
rect 22 1408 78 1464
rect 146 1408 202 1464
rect 270 1408 326 1464
rect 394 1408 450 1464
rect -474 1284 -418 1340
rect -350 1284 -294 1340
rect -226 1284 -170 1340
rect -102 1284 -46 1340
rect 22 1284 78 1340
rect 146 1284 202 1340
rect 270 1284 326 1340
rect 394 1284 450 1340
rect -474 1160 -418 1216
rect -350 1160 -294 1216
rect -226 1160 -170 1216
rect -102 1160 -46 1216
rect 22 1160 78 1216
rect 146 1160 202 1216
rect 270 1160 326 1216
rect 394 1160 450 1216
rect -474 1036 -418 1092
rect -350 1036 -294 1092
rect -226 1036 -170 1092
rect -102 1036 -46 1092
rect 22 1036 78 1092
rect 146 1036 202 1092
rect 270 1036 326 1092
rect 394 1036 450 1092
rect -474 912 -418 968
rect -350 912 -294 968
rect -226 912 -170 968
rect -102 912 -46 968
rect 22 912 78 968
rect 146 912 202 968
rect 270 912 326 968
rect 394 912 450 968
rect -474 788 -418 844
rect -350 788 -294 844
rect -226 788 -170 844
rect -102 788 -46 844
rect 22 788 78 844
rect 146 788 202 844
rect 270 788 326 844
rect 394 788 450 844
rect -474 664 -418 720
rect -350 664 -294 720
rect -226 664 -170 720
rect -102 664 -46 720
rect 22 664 78 720
rect 146 664 202 720
rect 270 664 326 720
rect 394 664 450 720
<< metal3 >>
rect -511 1588 489 2425
rect 714 2133 1714 2425
rect 714 2077 752 2133
rect 808 2077 876 2133
rect 932 2077 1000 2133
rect 1056 2077 1124 2133
rect 1180 2077 1248 2133
rect 1304 2077 1372 2133
rect 1428 2077 1496 2133
rect 1552 2077 1620 2133
rect 1676 2077 1714 2133
rect 714 2009 1714 2077
rect 714 1953 752 2009
rect 808 1953 876 2009
rect 932 1953 1000 2009
rect 1056 1953 1124 2009
rect 1180 1953 1248 2009
rect 1304 1953 1372 2009
rect 1428 1953 1496 2009
rect 1552 1953 1620 2009
rect 1676 1953 1714 2009
rect 714 1885 1714 1953
rect 714 1829 752 1885
rect 808 1829 876 1885
rect 932 1829 1000 1885
rect 1056 1829 1124 1885
rect 1180 1829 1248 1885
rect 1304 1829 1372 1885
rect 1428 1829 1496 1885
rect 1552 1829 1620 1885
rect 1676 1829 1714 1885
rect 714 1817 1714 1829
rect -511 1532 -474 1588
rect -418 1532 -350 1588
rect -294 1532 -226 1588
rect -170 1532 -102 1588
rect -46 1532 22 1588
rect 78 1532 146 1588
rect 202 1532 270 1588
rect 326 1532 394 1588
rect 450 1532 489 1588
rect -511 1464 489 1532
rect -511 1408 -474 1464
rect -418 1408 -350 1464
rect -294 1408 -226 1464
rect -170 1408 -102 1464
rect -46 1408 22 1464
rect 78 1408 146 1464
rect 202 1408 270 1464
rect 326 1408 394 1464
rect 450 1408 489 1464
rect -511 1340 489 1408
rect -511 1284 -474 1340
rect -418 1284 -350 1340
rect -294 1284 -226 1340
rect -170 1284 -102 1340
rect -46 1284 22 1340
rect 78 1284 146 1340
rect 202 1284 270 1340
rect 326 1284 394 1340
rect 450 1284 489 1340
rect -511 1216 489 1284
rect -511 1160 -474 1216
rect -418 1160 -350 1216
rect -294 1160 -226 1216
rect -170 1160 -102 1216
rect -46 1160 22 1216
rect 78 1160 146 1216
rect 202 1160 270 1216
rect 326 1160 394 1216
rect 450 1160 489 1216
rect -511 1092 489 1160
rect -511 1036 -474 1092
rect -418 1036 -350 1092
rect -294 1036 -226 1092
rect -170 1036 -102 1092
rect -46 1036 22 1092
rect 78 1036 146 1092
rect 202 1036 270 1092
rect 326 1036 394 1092
rect 450 1036 489 1092
rect -511 968 489 1036
rect -511 912 -474 968
rect -418 912 -350 968
rect -294 912 -226 968
rect -170 912 -102 968
rect -46 912 22 968
rect 78 912 146 968
rect 202 912 270 968
rect 326 912 394 968
rect 450 912 489 968
rect -511 844 489 912
rect -511 788 -474 844
rect -418 788 -350 844
rect -294 788 -226 844
rect -170 788 -102 844
rect -46 788 22 844
rect 78 788 146 844
rect 202 788 270 844
rect 326 788 394 844
rect 450 788 489 844
rect -511 720 489 788
rect -511 664 -474 720
rect -418 664 -350 720
rect -294 664 -226 720
rect -170 664 -102 720
rect -46 664 22 720
rect 78 664 146 720
rect 202 664 270 720
rect 326 664 394 720
rect 450 664 489 720
rect -511 625 489 664
use M2_M14310590878179_256x8m81  M2_M14310590878179_256x8m81_0
timestamp 1749760379
transform 1 0 1214 0 1 1981
box 0 0 1 1
use M3_M24310590878178_256x8m81  M3_M24310590878178_256x8m81_0
timestamp 1749760379
transform 1 0 1214 0 1 1981
box 0 0 1 1
use M3_M24310590878180_256x8m81  M3_M24310590878180_256x8m81_0
timestamp 1749760379
transform 1 0 -12 0 1 1126
box 0 0 1 1
<< properties >>
string GDS_END 1878186
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1877800
string path -0.055 12.125 -0.055 3.125 
<< end >>
