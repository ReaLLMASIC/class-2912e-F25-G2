magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< isosubstrate >>
rect 1479 -83 2795 2911
<< nwell >>
rect -83 1213 1139 2911
rect 1479 1213 2795 2911
rect 669 -711 1197 -183
rect 1547 -711 2075 -183
<< mvnmos >>
rect 354 270 494 870
rect 598 270 738 870
rect 1999 270 2139 870
rect 2243 270 2383 870
<< mvpmos >>
rect 354 1958 494 2558
rect 598 1958 738 2558
rect 1999 1358 2139 2558
rect 2243 1358 2383 2558
<< mvndiff >>
rect 266 857 354 870
rect 266 811 279 857
rect 325 811 354 857
rect 266 752 354 811
rect 266 706 279 752
rect 325 706 354 752
rect 266 647 354 706
rect 266 601 279 647
rect 325 601 354 647
rect 266 541 354 601
rect 266 495 279 541
rect 325 495 354 541
rect 266 435 354 495
rect 266 389 279 435
rect 325 389 354 435
rect 266 329 354 389
rect 266 283 279 329
rect 325 283 354 329
rect 266 270 354 283
rect 494 857 598 870
rect 494 811 523 857
rect 569 811 598 857
rect 494 752 598 811
rect 494 706 523 752
rect 569 706 598 752
rect 494 647 598 706
rect 494 601 523 647
rect 569 601 598 647
rect 494 541 598 601
rect 494 495 523 541
rect 569 495 598 541
rect 494 435 598 495
rect 494 389 523 435
rect 569 389 598 435
rect 494 329 598 389
rect 494 283 523 329
rect 569 283 598 329
rect 494 270 598 283
rect 738 857 826 870
rect 738 811 767 857
rect 813 811 826 857
rect 738 752 826 811
rect 738 706 767 752
rect 813 706 826 752
rect 738 647 826 706
rect 738 601 767 647
rect 813 601 826 647
rect 738 541 826 601
rect 738 495 767 541
rect 813 495 826 541
rect 738 435 826 495
rect 738 389 767 435
rect 813 389 826 435
rect 738 329 826 389
rect 738 283 767 329
rect 813 283 826 329
rect 738 270 826 283
rect 1911 857 1999 870
rect 1911 811 1924 857
rect 1970 811 1999 857
rect 1911 752 1999 811
rect 1911 706 1924 752
rect 1970 706 1999 752
rect 1911 647 1999 706
rect 1911 601 1924 647
rect 1970 601 1999 647
rect 1911 541 1999 601
rect 1911 495 1924 541
rect 1970 495 1999 541
rect 1911 435 1999 495
rect 1911 389 1924 435
rect 1970 389 1999 435
rect 1911 329 1999 389
rect 1911 283 1924 329
rect 1970 283 1999 329
rect 1911 270 1999 283
rect 2139 857 2243 870
rect 2139 811 2168 857
rect 2214 811 2243 857
rect 2139 752 2243 811
rect 2139 706 2168 752
rect 2214 706 2243 752
rect 2139 647 2243 706
rect 2139 601 2168 647
rect 2214 601 2243 647
rect 2139 541 2243 601
rect 2139 495 2168 541
rect 2214 495 2243 541
rect 2139 435 2243 495
rect 2139 389 2168 435
rect 2214 389 2243 435
rect 2139 329 2243 389
rect 2139 283 2168 329
rect 2214 283 2243 329
rect 2139 270 2243 283
rect 2383 857 2471 870
rect 2383 811 2412 857
rect 2458 811 2471 857
rect 2383 752 2471 811
rect 2383 706 2412 752
rect 2458 706 2471 752
rect 2383 647 2471 706
rect 2383 601 2412 647
rect 2458 601 2471 647
rect 2383 541 2471 601
rect 2383 495 2412 541
rect 2458 495 2471 541
rect 2383 435 2471 495
rect 2383 389 2412 435
rect 2458 389 2471 435
rect 2383 329 2471 389
rect 2383 283 2412 329
rect 2458 283 2471 329
rect 2383 270 2471 283
<< mvpdiff >>
rect 266 2545 354 2558
rect 266 2499 279 2545
rect 325 2499 354 2545
rect 266 2440 354 2499
rect 266 2394 279 2440
rect 325 2394 354 2440
rect 266 2335 354 2394
rect 266 2289 279 2335
rect 325 2289 354 2335
rect 266 2229 354 2289
rect 266 2183 279 2229
rect 325 2183 354 2229
rect 266 2123 354 2183
rect 266 2077 279 2123
rect 325 2077 354 2123
rect 266 2017 354 2077
rect 266 1971 279 2017
rect 325 1971 354 2017
rect 266 1958 354 1971
rect 494 2545 598 2558
rect 494 2499 523 2545
rect 569 2499 598 2545
rect 494 2440 598 2499
rect 494 2394 523 2440
rect 569 2394 598 2440
rect 494 2335 598 2394
rect 494 2289 523 2335
rect 569 2289 598 2335
rect 494 2229 598 2289
rect 494 2183 523 2229
rect 569 2183 598 2229
rect 494 2123 598 2183
rect 494 2077 523 2123
rect 569 2077 598 2123
rect 494 2017 598 2077
rect 494 1971 523 2017
rect 569 1971 598 2017
rect 494 1958 598 1971
rect 738 2545 826 2558
rect 738 2499 767 2545
rect 813 2499 826 2545
rect 738 2440 826 2499
rect 738 2394 767 2440
rect 813 2394 826 2440
rect 738 2335 826 2394
rect 738 2289 767 2335
rect 813 2289 826 2335
rect 738 2229 826 2289
rect 738 2183 767 2229
rect 813 2183 826 2229
rect 738 2123 826 2183
rect 738 2077 767 2123
rect 813 2077 826 2123
rect 738 2017 826 2077
rect 738 1971 767 2017
rect 813 1971 826 2017
rect 738 1958 826 1971
rect 1911 2545 1999 2558
rect 1911 1989 1924 2545
rect 1970 1989 1999 2545
rect 1911 1932 1999 1989
rect 1911 1886 1924 1932
rect 1970 1886 1999 1932
rect 1911 1829 1999 1886
rect 1911 1783 1924 1829
rect 1970 1783 1999 1829
rect 1911 1726 1999 1783
rect 1911 1680 1924 1726
rect 1970 1680 1999 1726
rect 1911 1623 1999 1680
rect 1911 1577 1924 1623
rect 1970 1577 1999 1623
rect 1911 1520 1999 1577
rect 1911 1474 1924 1520
rect 1970 1474 1999 1520
rect 1911 1417 1999 1474
rect 1911 1371 1924 1417
rect 1970 1371 1999 1417
rect 1911 1358 1999 1371
rect 2139 2545 2243 2558
rect 2139 1989 2168 2545
rect 2214 1989 2243 2545
rect 2139 1932 2243 1989
rect 2139 1886 2168 1932
rect 2214 1886 2243 1932
rect 2139 1829 2243 1886
rect 2139 1783 2168 1829
rect 2214 1783 2243 1829
rect 2139 1726 2243 1783
rect 2139 1680 2168 1726
rect 2214 1680 2243 1726
rect 2139 1623 2243 1680
rect 2139 1577 2168 1623
rect 2214 1577 2243 1623
rect 2139 1520 2243 1577
rect 2139 1474 2168 1520
rect 2214 1474 2243 1520
rect 2139 1417 2243 1474
rect 2139 1371 2168 1417
rect 2214 1371 2243 1417
rect 2139 1358 2243 1371
rect 2383 2545 2471 2558
rect 2383 1989 2412 2545
rect 2458 1989 2471 2545
rect 2383 1932 2471 1989
rect 2383 1886 2412 1932
rect 2458 1886 2471 1932
rect 2383 1829 2471 1886
rect 2383 1783 2412 1829
rect 2458 1783 2471 1829
rect 2383 1726 2471 1783
rect 2383 1680 2412 1726
rect 2458 1680 2471 1726
rect 2383 1623 2471 1680
rect 2383 1577 2412 1623
rect 2458 1577 2471 1623
rect 2383 1520 2471 1577
rect 2383 1474 2412 1520
rect 2458 1474 2471 1520
rect 2383 1417 2471 1474
rect 2383 1371 2412 1417
rect 2458 1371 2471 1417
rect 2383 1358 2471 1371
<< mvndiffc >>
rect 279 811 325 857
rect 279 706 325 752
rect 279 601 325 647
rect 279 495 325 541
rect 279 389 325 435
rect 279 283 325 329
rect 523 811 569 857
rect 523 706 569 752
rect 523 601 569 647
rect 523 495 569 541
rect 523 389 569 435
rect 523 283 569 329
rect 767 811 813 857
rect 767 706 813 752
rect 767 601 813 647
rect 767 495 813 541
rect 767 389 813 435
rect 767 283 813 329
rect 1924 811 1970 857
rect 1924 706 1970 752
rect 1924 601 1970 647
rect 1924 495 1970 541
rect 1924 389 1970 435
rect 1924 283 1970 329
rect 2168 811 2214 857
rect 2168 706 2214 752
rect 2168 601 2214 647
rect 2168 495 2214 541
rect 2168 389 2214 435
rect 2168 283 2214 329
rect 2412 811 2458 857
rect 2412 706 2458 752
rect 2412 601 2458 647
rect 2412 495 2458 541
rect 2412 389 2458 435
rect 2412 283 2458 329
<< mvpdiffc >>
rect 279 2499 325 2545
rect 279 2394 325 2440
rect 279 2289 325 2335
rect 279 2183 325 2229
rect 279 2077 325 2123
rect 279 1971 325 2017
rect 523 2499 569 2545
rect 523 2394 569 2440
rect 523 2289 569 2335
rect 523 2183 569 2229
rect 523 2077 569 2123
rect 523 1971 569 2017
rect 767 2499 813 2545
rect 767 2394 813 2440
rect 767 2289 813 2335
rect 767 2183 813 2229
rect 767 2077 813 2123
rect 767 1971 813 2017
rect 1924 1989 1970 2545
rect 1924 1886 1970 1932
rect 1924 1783 1970 1829
rect 1924 1680 1970 1726
rect 1924 1577 1970 1623
rect 1924 1474 1970 1520
rect 1924 1371 1970 1417
rect 2168 1989 2214 2545
rect 2168 1886 2214 1932
rect 2168 1783 2214 1829
rect 2168 1680 2214 1726
rect 2168 1577 2214 1623
rect 2168 1474 2214 1520
rect 2168 1371 2214 1417
rect 2412 1989 2458 2545
rect 2412 1886 2458 1932
rect 2412 1783 2458 1829
rect 2412 1680 2458 1726
rect 2412 1577 2458 1623
rect 2412 1474 2458 1520
rect 2412 1371 2458 1417
<< psubdiff >>
rect 0 1008 90 1030
rect 0 22 22 1008
rect 68 90 90 1008
rect 966 914 1056 936
rect 966 90 988 914
rect 68 68 988 90
rect 68 22 176 68
rect 880 22 988 68
rect 1034 22 1056 914
rect 0 0 1056 22
rect 1562 914 1652 936
rect 1562 22 1584 914
rect 1630 90 1652 914
rect 2622 1008 2712 1030
rect 2622 90 2644 1008
rect 1630 68 2644 90
rect 1630 22 1738 68
rect 2536 22 2644 68
rect 2690 22 2712 1008
rect 1562 0 2712 22
<< nsubdiff >>
rect 0 2806 1056 2828
rect 0 1350 22 2806
rect 68 2760 176 2806
rect 880 2760 988 2806
rect 68 2738 988 2760
rect 68 1350 90 2738
rect 0 1328 90 1350
rect 966 1350 988 2738
rect 1034 1350 1056 2806
rect 966 1328 1056 1350
rect 1562 2806 2712 2828
rect 1562 1350 1584 2806
rect 1630 2760 1738 2806
rect 2536 2760 2644 2806
rect 1630 2738 2644 2760
rect 1630 1350 1652 2738
rect 1562 1328 1652 1350
rect 2622 1350 2644 2738
rect 2690 1350 2712 2806
rect 2622 1328 2712 1350
<< mvnsubdiff >>
rect 717 -244 1149 -231
rect 717 -290 730 -244
rect 776 -290 850 -244
rect 896 -290 970 -244
rect 1016 -290 1090 -244
rect 1136 -290 1149 -244
rect 717 -303 1149 -290
rect 717 -364 789 -303
rect 717 -410 730 -364
rect 776 -410 789 -364
rect 1077 -364 1149 -303
rect 717 -484 789 -410
rect 717 -530 730 -484
rect 776 -530 789 -484
rect 1077 -410 1090 -364
rect 1136 -410 1149 -364
rect 1077 -484 1149 -410
rect 717 -591 789 -530
rect 1077 -530 1090 -484
rect 1136 -530 1149 -484
rect 1077 -591 1149 -530
rect 717 -604 1149 -591
rect 717 -650 730 -604
rect 776 -650 850 -604
rect 896 -650 970 -604
rect 1016 -650 1090 -604
rect 1136 -650 1149 -604
rect 717 -663 1149 -650
rect 1595 -244 2027 -231
rect 1595 -290 1608 -244
rect 1654 -290 1728 -244
rect 1774 -290 1848 -244
rect 1894 -290 1968 -244
rect 2014 -290 2027 -244
rect 1595 -303 2027 -290
rect 1595 -364 1667 -303
rect 1595 -410 1608 -364
rect 1654 -410 1667 -364
rect 1955 -364 2027 -303
rect 1595 -484 1667 -410
rect 1595 -530 1608 -484
rect 1654 -530 1667 -484
rect 1955 -410 1968 -364
rect 2014 -410 2027 -364
rect 1955 -484 2027 -410
rect 1595 -591 1667 -530
rect 1955 -530 1968 -484
rect 2014 -530 2027 -484
rect 1955 -591 2027 -530
rect 1595 -604 2027 -591
rect 1595 -650 1608 -604
rect 1654 -650 1728 -604
rect 1774 -650 1848 -604
rect 1894 -650 1968 -604
rect 2014 -650 2027 -604
rect 1595 -663 2027 -650
<< psubdiffcont >>
rect 22 22 68 1008
rect 176 22 880 68
rect 988 22 1034 914
rect 1584 22 1630 914
rect 1738 22 2536 68
rect 2644 22 2690 1008
<< nsubdiffcont >>
rect 22 1350 68 2806
rect 176 2760 880 2806
rect 988 1350 1034 2806
rect 1584 1350 1630 2806
rect 1738 2760 2536 2806
rect 2644 1350 2690 2806
<< mvnsubdiffcont >>
rect 730 -290 776 -244
rect 850 -290 896 -244
rect 970 -290 1016 -244
rect 1090 -290 1136 -244
rect 730 -410 776 -364
rect 730 -530 776 -484
rect 1090 -410 1136 -364
rect 1090 -530 1136 -484
rect 730 -650 776 -604
rect 850 -650 896 -604
rect 970 -650 1016 -604
rect 1090 -650 1136 -604
rect 1608 -290 1654 -244
rect 1728 -290 1774 -244
rect 1848 -290 1894 -244
rect 1968 -290 2014 -244
rect 1608 -410 1654 -364
rect 1608 -530 1654 -484
rect 1968 -410 2014 -364
rect 1968 -530 2014 -484
rect 1608 -650 1654 -604
rect 1728 -650 1774 -604
rect 1848 -650 1894 -604
rect 1968 -650 2014 -604
<< polysilicon >>
rect 354 2558 494 2602
rect 598 2558 738 2602
rect 354 1537 494 1958
rect 354 1397 401 1537
rect 447 1397 494 1537
rect 354 870 494 1397
rect 598 1537 738 1958
rect 598 1397 645 1537
rect 691 1397 738 1537
rect 598 870 738 1397
rect 1999 2558 2139 2602
rect 2243 2558 2383 2602
rect 1999 1213 2139 1358
rect 1783 1178 2139 1213
rect 1783 1038 1802 1178
rect 1848 1038 2139 1178
rect 1783 1002 2139 1038
rect 354 226 494 270
rect 598 226 738 270
rect 1999 870 2139 1002
rect 2243 1178 2383 1358
rect 2243 1038 2282 1178
rect 2328 1038 2383 1178
rect 2243 870 2383 1038
rect 1999 226 2139 270
rect 2243 226 2383 270
<< polycontact >>
rect 401 1397 447 1537
rect 645 1397 691 1537
rect 1802 1038 1848 1178
rect 2282 1038 2328 1178
<< mvpdiode >>
rect 885 -424 981 -399
rect 885 -470 910 -424
rect 956 -470 981 -424
rect 885 -495 981 -470
rect 1763 -424 1859 -399
rect 1763 -470 1788 -424
rect 1834 -470 1859 -424
rect 1763 -495 1859 -470
<< mvpdiodec >>
rect 910 -470 956 -424
rect 1788 -470 1834 -424
<< metal1 >>
rect 11 2806 1045 2817
rect 11 1350 22 2806
rect 68 2760 176 2806
rect 880 2760 988 2806
rect 68 2749 988 2760
rect 68 1350 79 2749
rect 264 2545 340 2749
rect 264 2499 279 2545
rect 325 2499 340 2545
rect 264 2440 340 2499
rect 264 2394 279 2440
rect 325 2394 340 2440
rect 264 2335 340 2394
rect 264 2289 279 2335
rect 325 2289 340 2335
rect 264 2229 340 2289
rect 264 2183 279 2229
rect 325 2183 340 2229
rect 264 2123 340 2183
rect 264 2077 279 2123
rect 325 2077 340 2123
rect 264 2017 340 2077
rect 264 1971 279 2017
rect 325 1971 340 2017
rect 264 1958 340 1971
rect 508 2545 584 2558
rect 508 2499 523 2545
rect 569 2499 584 2545
rect 508 2440 584 2499
rect 508 2394 523 2440
rect 569 2394 584 2440
rect 508 2335 584 2394
rect 508 2289 523 2335
rect 569 2289 584 2335
rect 508 2229 584 2289
rect 508 2183 523 2229
rect 569 2183 584 2229
rect 508 2123 584 2183
rect 508 2077 523 2123
rect 569 2077 584 2123
rect 508 2017 584 2077
rect 508 1971 523 2017
rect 569 1971 584 2017
rect 508 1794 584 1971
rect 752 2545 828 2749
rect 752 2499 767 2545
rect 813 2499 828 2545
rect 752 2440 828 2499
rect 752 2394 767 2440
rect 813 2394 828 2440
rect 752 2335 828 2394
rect 752 2289 767 2335
rect 813 2289 828 2335
rect 752 2229 828 2289
rect 752 2183 767 2229
rect 813 2183 828 2229
rect 752 2123 828 2183
rect 752 2077 767 2123
rect 813 2077 828 2123
rect 752 2017 828 2077
rect 752 1971 767 2017
rect 813 1971 828 2017
rect 752 1958 828 1971
rect 508 1718 828 1794
rect 386 1544 462 1556
rect 386 1388 398 1544
rect 450 1388 462 1544
rect 386 1376 462 1388
rect 630 1544 706 1556
rect 630 1388 642 1544
rect 694 1388 706 1544
rect 630 1376 706 1388
rect 11 1339 79 1350
rect 752 1197 828 1718
rect 977 1350 988 2749
rect 1034 1350 1045 2806
rect 977 1339 1045 1350
rect 1573 2806 2701 2817
rect 1573 1350 1584 2806
rect 1630 2760 1738 2806
rect 2536 2760 2644 2806
rect 1630 2749 2644 2760
rect 1630 1350 1641 2749
rect 1573 1339 1641 1350
rect 1909 2545 1985 2558
rect 1909 1989 1924 2545
rect 1970 1989 1985 2545
rect 1909 1932 1985 1989
rect 1909 1886 1924 1932
rect 1970 1886 1985 1932
rect 1909 1829 1985 1886
rect 1909 1783 1924 1829
rect 1970 1783 1985 1829
rect 1909 1726 1985 1783
rect 1909 1680 1924 1726
rect 1970 1680 1985 1726
rect 1909 1623 1985 1680
rect 1909 1577 1924 1623
rect 1970 1577 1985 1623
rect 1909 1520 1985 1577
rect 1909 1474 1924 1520
rect 1970 1474 1985 1520
rect 1909 1417 1985 1474
rect 1909 1371 1924 1417
rect 1970 1371 1985 1417
rect 1909 1197 1985 1371
rect 2153 2545 2229 2749
rect 2153 1989 2168 2545
rect 2214 1989 2229 2545
rect 2153 1932 2229 1989
rect 2153 1886 2168 1932
rect 2214 1886 2229 1932
rect 2153 1829 2229 1886
rect 2153 1783 2168 1829
rect 2214 1783 2229 1829
rect 2153 1726 2229 1783
rect 2153 1680 2168 1726
rect 2214 1680 2229 1726
rect 2153 1623 2229 1680
rect 2153 1577 2168 1623
rect 2214 1577 2229 1623
rect 2153 1520 2229 1577
rect 2153 1474 2168 1520
rect 2214 1474 2229 1520
rect 2153 1417 2229 1474
rect 2153 1371 2168 1417
rect 2214 1371 2229 1417
rect 2153 1358 2229 1371
rect 2397 2545 2473 2558
rect 2397 1989 2412 2545
rect 2458 1989 2473 2545
rect 2397 1932 2473 1989
rect 2397 1886 2412 1932
rect 2458 1886 2473 1932
rect 2397 1829 2473 1886
rect 2397 1783 2412 1829
rect 2458 1783 2473 1829
rect 2397 1726 2473 1783
rect 2397 1680 2412 1726
rect 2458 1680 2473 1726
rect 2397 1623 2473 1680
rect 2397 1577 2412 1623
rect 2458 1577 2473 1623
rect 2397 1520 2473 1577
rect 2397 1474 2412 1520
rect 2458 1474 2473 1520
rect 2397 1417 2473 1474
rect 2397 1371 2412 1417
rect 2458 1371 2473 1417
rect 752 1189 1804 1197
rect 752 1178 1859 1189
rect 752 1038 1802 1178
rect 1848 1038 1859 1178
rect 752 1027 1859 1038
rect 1909 1178 2347 1197
rect 1909 1038 2282 1178
rect 2328 1038 2347 1178
rect 752 1019 1804 1027
rect 1909 1019 2347 1038
rect 11 1008 79 1019
rect 11 22 22 1008
rect 68 79 79 1008
rect 264 857 340 870
rect 264 811 279 857
rect 325 811 340 857
rect 264 752 340 811
rect 264 706 279 752
rect 325 706 340 752
rect 264 647 340 706
rect 264 601 279 647
rect 325 601 340 647
rect 264 541 340 601
rect 264 495 279 541
rect 325 495 340 541
rect 264 435 340 495
rect 264 389 279 435
rect 325 389 340 435
rect 264 329 340 389
rect 264 283 279 329
rect 325 283 340 329
rect 264 79 340 283
rect 523 857 569 870
rect 523 752 569 811
rect 523 647 569 706
rect 523 541 569 601
rect 523 435 569 495
rect 523 329 569 389
rect 523 270 569 283
rect 752 857 828 1019
rect 752 811 767 857
rect 813 811 828 857
rect 752 752 828 811
rect 752 706 767 752
rect 813 706 828 752
rect 752 647 828 706
rect 752 601 767 647
rect 813 601 828 647
rect 752 541 828 601
rect 752 495 767 541
rect 813 495 828 541
rect 752 435 828 495
rect 752 389 767 435
rect 813 389 828 435
rect 752 329 828 389
rect 752 283 767 329
rect 813 283 828 329
rect 752 270 828 283
rect 977 914 1045 925
rect 977 87 988 914
rect 865 79 988 87
rect 68 75 988 79
rect 68 68 877 75
rect 68 22 176 68
rect 880 22 988 23
rect 1034 22 1045 914
rect 1573 914 1641 925
rect 11 11 1045 22
rect 1115 179 1191 191
rect 1115 23 1127 179
rect 1179 23 1191 179
rect 1115 -81 1191 23
rect 1573 22 1584 914
rect 1630 79 1641 914
rect 1909 857 1985 1019
rect 1909 811 1924 857
rect 1970 811 1985 857
rect 1909 752 1985 811
rect 1909 706 1924 752
rect 1970 706 1985 752
rect 1909 647 1985 706
rect 1909 601 1924 647
rect 1970 601 1985 647
rect 1909 541 1985 601
rect 1909 495 1924 541
rect 1970 495 1985 541
rect 1909 435 1985 495
rect 1909 389 1924 435
rect 1970 389 1985 435
rect 1909 329 1985 389
rect 1909 283 1924 329
rect 1970 283 1985 329
rect 1909 270 1985 283
rect 2153 857 2229 870
rect 2153 811 2168 857
rect 2214 811 2229 857
rect 2153 752 2229 811
rect 2153 706 2168 752
rect 2214 706 2229 752
rect 2153 647 2229 706
rect 2153 601 2168 647
rect 2214 601 2229 647
rect 2153 541 2229 601
rect 2153 495 2168 541
rect 2214 495 2229 541
rect 2153 435 2229 495
rect 2153 389 2168 435
rect 2214 389 2229 435
rect 2153 329 2229 389
rect 2153 283 2168 329
rect 2214 283 2229 329
rect 2153 79 2229 283
rect 2397 857 2473 1371
rect 2633 1350 2644 2749
rect 2690 1350 2701 2806
rect 2633 1339 2701 1350
rect 2397 811 2412 857
rect 2458 811 2473 857
rect 2397 752 2473 811
rect 2397 706 2412 752
rect 2458 706 2473 752
rect 2397 647 2473 706
rect 2397 601 2412 647
rect 2458 601 2473 647
rect 2397 541 2473 601
rect 2397 495 2412 541
rect 2458 495 2473 541
rect 2397 435 2473 495
rect 2397 389 2412 435
rect 2458 389 2473 435
rect 2397 329 2473 389
rect 2397 283 2412 329
rect 2458 283 2473 329
rect 2397 270 2473 283
rect 2633 1008 2701 1019
rect 2633 79 2644 1008
rect 1630 68 2644 79
rect 1630 22 1738 68
rect 2536 22 2644 68
rect 2690 22 2701 1008
rect 1573 11 2701 22
rect 1115 -157 1671 -81
rect 1595 -231 1671 -157
rect 386 -243 1149 -231
rect 386 -399 398 -243
rect 450 -244 1149 -243
rect 450 -290 730 -244
rect 776 -290 850 -244
rect 896 -290 970 -244
rect 1016 -290 1090 -244
rect 1136 -290 1149 -244
rect 450 -303 1149 -290
rect 450 -364 789 -303
rect 450 -399 730 -364
rect 386 -410 730 -399
rect 776 -410 789 -364
rect 1077 -364 1149 -303
rect 386 -411 789 -410
rect 717 -484 789 -411
rect 717 -530 730 -484
rect 776 -530 789 -484
rect 885 -421 981 -399
rect 885 -473 907 -421
rect 959 -473 981 -421
rect 885 -495 981 -473
rect 1077 -410 1090 -364
rect 1136 -410 1149 -364
rect 1077 -484 1149 -410
rect 717 -591 789 -530
rect 1077 -530 1090 -484
rect 1136 -530 1149 -484
rect 1077 -591 1149 -530
rect 717 -604 1149 -591
rect 717 -650 730 -604
rect 776 -650 850 -604
rect 896 -650 970 -604
rect 1016 -650 1090 -604
rect 1136 -650 1149 -604
rect 717 -663 1149 -650
rect 1595 -244 2027 -231
rect 1595 -290 1608 -244
rect 1654 -290 1728 -244
rect 1774 -290 1848 -244
rect 1894 -290 1968 -244
rect 2014 -290 2027 -244
rect 1595 -303 2027 -290
rect 1595 -364 1667 -303
rect 1595 -410 1608 -364
rect 1654 -410 1667 -364
rect 1955 -364 2027 -303
rect 1595 -484 1667 -410
rect 1595 -530 1608 -484
rect 1654 -530 1667 -484
rect 1763 -421 1859 -399
rect 1763 -473 1785 -421
rect 1837 -473 1859 -421
rect 1763 -495 1859 -473
rect 1955 -410 1968 -364
rect 2014 -410 2027 -364
rect 1955 -484 2027 -410
rect 1595 -591 1667 -530
rect 1955 -530 1968 -484
rect 2014 -530 2027 -484
rect 1955 -591 2027 -530
rect 1595 -604 2027 -591
rect 1595 -650 1608 -604
rect 1654 -650 1728 -604
rect 1774 -650 1848 -604
rect 1894 -650 1968 -604
rect 2014 -650 2027 -604
rect 1595 -663 2027 -650
rect 895 -739 1953 -727
rect 895 -791 907 -739
rect 1063 -791 1785 -739
rect 1941 -791 1953 -739
rect 895 -803 1953 -791
<< via1 >>
rect 398 1537 450 1544
rect 398 1397 401 1537
rect 401 1397 447 1537
rect 447 1397 450 1537
rect 398 1388 450 1397
rect 642 1537 694 1544
rect 642 1397 645 1537
rect 645 1397 691 1537
rect 691 1397 694 1537
rect 642 1388 694 1397
rect 877 68 988 75
rect 877 23 880 68
rect 880 23 988 68
rect 988 23 1033 75
rect 1127 23 1179 179
rect 398 -399 450 -243
rect 907 -424 959 -421
rect 907 -470 910 -424
rect 910 -470 956 -424
rect 956 -470 959 -424
rect 907 -473 959 -470
rect 1785 -424 1837 -421
rect 1785 -470 1788 -424
rect 1788 -470 1834 -424
rect 1834 -470 1837 -424
rect 1785 -473 1837 -470
rect 907 -791 1063 -739
rect 1785 -791 1941 -739
<< metal2 >>
rect 386 1544 462 1556
rect 386 1388 398 1544
rect 450 1388 462 1544
rect 386 -243 462 1388
rect 630 1544 1191 1556
rect 630 1388 642 1544
rect 694 1388 1191 1544
rect 630 1376 1191 1388
rect 1115 179 1191 1376
rect 865 75 1045 87
rect 865 23 877 75
rect 1033 23 1045 75
rect 865 11 1045 23
rect 1115 23 1127 179
rect 1179 23 1191 179
rect 1115 11 1191 23
rect 386 -399 398 -243
rect 450 -399 462 -243
rect 386 -411 462 -399
rect 895 -421 971 11
rect 895 -473 907 -421
rect 959 -473 971 -421
rect 895 -727 971 -473
rect 1773 -421 1849 -409
rect 1773 -473 1785 -421
rect 1837 -473 1849 -421
rect 1773 -727 1849 -473
rect 895 -739 1075 -727
rect 895 -791 907 -739
rect 1063 -791 1075 -739
rect 895 -803 1075 -791
rect 1773 -739 1953 -727
rect 1773 -791 1785 -739
rect 1941 -791 1953 -739
rect 1773 -803 1953 -791
use M1_NWELL_CDNS_40661953145218  M1_NWELL_CDNS_40661953145218_0
timestamp 1749760379
transform 1 0 528 0 1 2783
box 0 0 1 1
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_0
timestamp 1749760379
transform 1 0 45 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_1
timestamp 1749760379
transform 1 0 2667 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_2
timestamp 1749760379
transform 1 0 1607 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_3
timestamp 1749760379
transform 1 0 1011 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145225  M1_NWELL_CDNS_40661953145225_0
timestamp 1749760379
transform 1 0 2137 0 1 2783
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_0
timestamp 1749760379
transform -1 0 424 0 1 1467
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_1
timestamp 1749760379
transform -1 0 668 0 1 1467
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_2
timestamp 1749760379
transform 1 0 2305 0 1 1108
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_3
timestamp 1749760379
transform 1 0 1825 0 1 1108
box 0 0 1 1
use M1_PSUB_CDNS_40661953145221  M1_PSUB_CDNS_40661953145221_0
timestamp 1749760379
transform 1 0 2137 0 -1 45
box 0 0 1 1
use M1_PSUB_CDNS_40661953145224  M1_PSUB_CDNS_40661953145224_0
timestamp 1749760379
transform 1 0 528 0 -1 45
box 0 0 1 1
use M1_PSUB_CDNS_40661953145226  M1_PSUB_CDNS_40661953145226_0
timestamp 1749760379
transform 1 0 2667 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661953145226  M1_PSUB_CDNS_40661953145226_1
timestamp 1749760379
transform 1 0 45 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661953145228  M1_PSUB_CDNS_40661953145228_0
timestamp 1749760379
transform 1 0 1607 0 -1 468
box 0 0 1 1
use M1_PSUB_CDNS_40661953145228  M1_PSUB_CDNS_40661953145228_1
timestamp 1749760379
transform 1 0 1011 0 -1 468
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_0
timestamp 1749760379
transform 0 -1 1153 1 0 101
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_1
timestamp 1749760379
transform 1 0 985 0 1 -765
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_2
timestamp 1749760379
transform 1 0 955 0 1 49
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_3
timestamp 1749760379
transform 1 0 1863 0 1 -765
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_0
timestamp 1749760379
transform 1 0 424 0 1 -321
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_1
timestamp 1749760379
transform 1 0 668 0 1 1466
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_2
timestamp 1749760379
transform 1 0 424 0 1 1466
box 0 0 1 1
use M2_M1_CDNS_40661953145227  M2_M1_CDNS_40661953145227_0
timestamp 1749760379
transform 1 0 1811 0 1 -447
box 0 0 1 1
use M2_M1_CDNS_40661953145227  M2_M1_CDNS_40661953145227_1
timestamp 1749760379
transform 1 0 933 0 1 -447
box 0 0 1 1
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_0
timestamp 1749760379
transform -1 0 494 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_1
timestamp 1749760379
transform -1 0 738 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_2
timestamp 1749760379
transform 1 0 2243 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_3
timestamp 1749760379
transform 1 0 1999 0 1 270
box 0 0 1 1
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1749760379
transform 1 0 354 0 1 1958
box 0 0 1 1
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_1
timestamp 1749760379
transform 1 0 598 0 1 1958
box 0 0 1 1
use pmos_6p0_CDNS_4066195314513  pmos_6p0_CDNS_4066195314513_0
timestamp 1749760379
transform -1 0 2383 0 1 1358
box 0 0 1 1
use pmos_6p0_CDNS_4066195314513  pmos_6p0_CDNS_4066195314513_1
timestamp 1749760379
transform -1 0 2139 0 1 1358
box 0 0 1 1
use pn_6p0_CDNS_4066195314510  pn_6p0_CDNS_4066195314510_0
timestamp 1749760379
transform -1 0 981 0 -1 -399
box 0 0 1 1
use pn_6p0_CDNS_4066195314510  pn_6p0_CDNS_4066195314510_1
timestamp 1749760379
transform -1 0 1859 0 -1 -399
box 0 0 1 1
<< labels >>
rlabel metal1 s 667 1468 667 1468 4 OE
port 1 nsew
rlabel metal1 s 421 1468 421 1468 4 PDRV
port 2 nsew
rlabel metal1 s 2435 1100 2435 1100 4 ENB
port 3 nsew
rlabel metal1 s 75 2788 75 2788 4 VDD
port 4 nsew
rlabel metal1 s 256 45 256 45 4 VSS
port 5 nsew
rlabel metal1 s 2283 2788 2283 2788 4 DVDD
port 6 nsew
rlabel metal1 s 2290 45 2290 45 4 DVSS
port 7 nsew
rlabel metal1 s 2112 1100 2112 1100 4 EN
port 8 nsew
<< properties >>
string GDS_END 1502664
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1497672
string path 48.675 6.750 48.675 63.950 
<< end >>
