magic
tech gf180mcuD
timestamp 1749760379
<< properties >>
string GDS_END 8989580
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 8988040
<< end >>
