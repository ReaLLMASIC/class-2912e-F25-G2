magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< isosubstrate >>
rect -257 10974 13760 27678
rect -39 -129 13470 10974
<< metal1 >>
rect -360 10764 61 10914
rect -360 9776 -280 10764
rect -20 9776 61 10764
rect 843 10815 1780 10854
rect 843 10763 1001 10815
rect 1053 10763 1125 10815
rect 1177 10763 1780 10815
rect 843 10691 1780 10763
rect 843 10639 1001 10691
rect 1053 10639 1125 10691
rect 1177 10639 1780 10691
rect 843 10567 1780 10639
rect 843 10515 1001 10567
rect 1053 10515 1125 10567
rect 1177 10515 1780 10567
rect 843 10443 1780 10515
rect 843 10391 1001 10443
rect 1053 10391 1125 10443
rect 1177 10391 1780 10443
rect 843 10319 1780 10391
rect 843 10267 1001 10319
rect 1053 10267 1125 10319
rect 1177 10267 1780 10319
rect 843 10195 1780 10267
rect 843 10143 1001 10195
rect 1053 10143 1125 10195
rect 1177 10143 1780 10195
rect 843 10071 1780 10143
rect 843 10058 1001 10071
rect -360 8855 61 9776
rect 989 10019 1001 10058
rect 1053 10019 1125 10071
rect 1177 10058 1780 10071
rect 11780 10815 12701 10854
rect 11780 10763 12319 10815
rect 12371 10763 12443 10815
rect 12495 10763 12701 10815
rect 11780 10691 12701 10763
rect 11780 10639 12319 10691
rect 12371 10639 12443 10691
rect 12495 10639 12701 10691
rect 11780 10567 12701 10639
rect 11780 10515 12319 10567
rect 12371 10515 12443 10567
rect 12495 10515 12701 10567
rect 11780 10443 12701 10515
rect 11780 10391 12319 10443
rect 12371 10391 12443 10443
rect 12495 10391 12701 10443
rect 11780 10319 12701 10391
rect 11780 10267 12319 10319
rect 12371 10267 12443 10319
rect 12495 10267 12701 10319
rect 11780 10195 12701 10267
rect 11780 10143 12319 10195
rect 12371 10143 12443 10195
rect 12495 10143 12701 10195
rect 11780 10071 12701 10143
rect 11780 10058 12319 10071
rect 1177 10019 1189 10058
rect 989 9947 1189 10019
rect 989 9895 1001 9947
rect 1053 9895 1125 9947
rect 1177 9895 1189 9947
rect 989 9823 1189 9895
rect 989 9771 1001 9823
rect 1053 9771 1125 9823
rect 1177 9771 1189 9823
rect 989 9759 1189 9771
rect 12307 10019 12319 10058
rect 12371 10019 12443 10071
rect 12495 10058 12701 10071
rect 13375 10764 13796 10914
rect 12495 10019 12507 10058
rect 12307 9947 12507 10019
rect 12307 9895 12319 9947
rect 12371 9895 12443 9947
rect 12495 9895 12507 9947
rect 12307 9823 12507 9895
rect 12307 9771 12319 9823
rect 12371 9771 12443 9823
rect 12495 9771 12507 9823
rect 12307 9759 12507 9771
rect 13375 9776 13462 10764
rect 13722 9776 13796 10764
rect 1026 9510 1206 9522
rect 1026 9458 1038 9510
rect 1194 9458 1206 9510
rect 1026 9446 1206 9458
rect 12305 9510 12485 9522
rect 12305 9458 12317 9510
rect 12473 9458 12485 9510
rect 12305 9446 12485 9458
rect 1026 9344 1206 9356
rect 1026 9292 1038 9344
rect 1194 9292 1206 9344
rect 1026 9280 1206 9292
rect 12305 9344 12485 9356
rect 12305 9292 12317 9344
rect 12473 9292 12485 9344
rect 12305 9280 12485 9292
rect 1026 9184 1206 9196
rect 1026 9132 1038 9184
rect 1194 9132 1206 9184
rect 1026 9120 1206 9132
rect 12305 9184 12485 9196
rect 12305 9132 12317 9184
rect 12473 9132 12485 9184
rect 12305 9120 12485 9132
rect 1026 9018 1206 9030
rect 1026 8966 1038 9018
rect 1194 8966 1206 9018
rect 1026 8954 1206 8966
rect 12305 9018 12485 9030
rect 12305 8966 12317 9018
rect 12473 8966 12485 9018
rect 12305 8954 12485 8966
rect 13375 8877 13796 9776
rect -360 8434 1108 8855
rect 1741 8819 2142 8863
rect 1741 6583 1753 8819
rect 1805 6583 2142 8819
rect 1741 6273 2142 6583
rect 1741 3413 1753 6273
rect 1805 3413 2142 6273
rect 1741 3086 2142 3413
rect 1741 538 1753 3086
rect 1805 1243 2142 3086
rect 11290 8819 11732 8863
rect 11290 6583 11627 8819
rect 11679 6583 11732 8819
rect 12368 8456 13796 8877
rect 11290 6273 11732 6583
rect 11290 3413 11627 6273
rect 11679 3413 11732 6273
rect 11290 3086 11732 3413
rect 11290 1243 11627 3086
rect 1805 538 2127 1243
rect 11316 770 11627 1243
rect 1741 510 2127 538
rect 11290 538 11627 770
rect 11679 538 11732 3086
rect 11290 510 11732 538
<< via1 >>
rect -280 9776 -20 10764
rect 1001 10763 1053 10815
rect 1125 10763 1177 10815
rect 1001 10639 1053 10691
rect 1125 10639 1177 10691
rect 1001 10515 1053 10567
rect 1125 10515 1177 10567
rect 1001 10391 1053 10443
rect 1125 10391 1177 10443
rect 1001 10267 1053 10319
rect 1125 10267 1177 10319
rect 1001 10143 1053 10195
rect 1125 10143 1177 10195
rect 1001 10019 1053 10071
rect 1125 10019 1177 10071
rect 12319 10763 12371 10815
rect 12443 10763 12495 10815
rect 12319 10639 12371 10691
rect 12443 10639 12495 10691
rect 12319 10515 12371 10567
rect 12443 10515 12495 10567
rect 12319 10391 12371 10443
rect 12443 10391 12495 10443
rect 12319 10267 12371 10319
rect 12443 10267 12495 10319
rect 12319 10143 12371 10195
rect 12443 10143 12495 10195
rect 1001 9895 1053 9947
rect 1125 9895 1177 9947
rect 1001 9771 1053 9823
rect 1125 9771 1177 9823
rect 12319 10019 12371 10071
rect 12443 10019 12495 10071
rect 12319 9895 12371 9947
rect 12443 9895 12495 9947
rect 12319 9771 12371 9823
rect 12443 9771 12495 9823
rect 13462 9776 13722 10764
rect 1038 9458 1194 9510
rect 12317 9458 12473 9510
rect 1038 9292 1194 9344
rect 12317 9292 12473 9344
rect 1038 9132 1194 9184
rect 12317 9132 12473 9184
rect 1038 8966 1194 9018
rect 12317 8966 12473 9018
rect 1753 6583 1805 8819
rect 1753 3413 1805 6273
rect 1753 538 1805 3086
rect 11627 6583 11679 8819
rect 11627 3413 11679 6273
rect 11627 538 11679 3086
<< metal2 >>
rect -326 10818 34 10828
rect -326 10762 -316 10818
rect -260 10764 -174 10818
rect -118 10764 -32 10818
rect 24 10762 34 10818
rect -326 10676 -280 10762
rect -20 10676 34 10762
rect -326 10620 -316 10676
rect 24 10620 34 10676
rect -326 10534 -280 10620
rect -20 10534 34 10620
rect -326 10478 -316 10534
rect 24 10478 34 10534
rect -326 10392 -280 10478
rect -20 10392 34 10478
rect -326 10336 -316 10392
rect 24 10336 34 10392
rect -326 10250 -280 10336
rect -20 10250 34 10336
rect -326 10194 -316 10250
rect 24 10194 34 10250
rect -326 10108 -280 10194
rect -20 10108 34 10194
rect -326 10052 -316 10108
rect 24 10052 34 10108
rect -326 9966 -280 10052
rect -20 9966 34 10052
rect -326 9910 -316 9966
rect 24 9910 34 9966
rect -326 9824 -280 9910
rect -20 9824 34 9910
rect -326 9768 -316 9824
rect -260 9768 -174 9776
rect -118 9768 -32 9776
rect 24 9768 34 9824
rect -326 9758 34 9768
rect 213 9051 313 26936
rect 393 9211 493 26936
rect 573 9371 673 26936
rect 753 9539 861 26936
rect 1697 26000 11781 26600
rect 1697 23319 2941 26000
rect 3465 23319 4709 26000
rect 5233 23319 6477 26000
rect 7001 23319 8245 26000
rect 8769 23319 10013 26000
rect 10537 23319 11781 26000
rect 1697 12658 2941 15319
rect 3465 12658 4709 15319
rect 5233 12658 6477 15319
rect 7001 12658 8245 15319
rect 8769 12658 10013 15319
rect 10537 12658 11781 15319
rect 980 10818 1198 10828
rect 980 10762 990 10818
rect 1046 10815 1132 10818
rect 1053 10763 1125 10815
rect 1046 10762 1132 10763
rect 1188 10762 1198 10818
rect 980 10691 1198 10762
rect 980 10676 1001 10691
rect 980 10620 990 10676
rect 1053 10639 1125 10691
rect 1177 10676 1198 10691
rect 1046 10620 1132 10639
rect 1188 10620 1198 10676
rect 980 10567 1198 10620
rect 980 10534 1001 10567
rect 980 10478 990 10534
rect 1053 10515 1125 10567
rect 1177 10534 1198 10567
rect 1046 10478 1132 10515
rect 1188 10478 1198 10534
rect 980 10443 1198 10478
rect 980 10392 1001 10443
rect 980 10336 990 10392
rect 1053 10391 1125 10443
rect 1177 10392 1198 10443
rect 1046 10336 1132 10391
rect 1188 10336 1198 10392
rect 980 10319 1198 10336
rect 980 10267 1001 10319
rect 1053 10267 1125 10319
rect 1177 10267 1198 10319
rect 980 10250 1198 10267
rect 980 10194 990 10250
rect 1046 10195 1132 10250
rect 980 10143 1001 10194
rect 1053 10143 1125 10195
rect 1188 10194 1198 10250
rect 1177 10143 1198 10194
rect 980 10108 1198 10143
rect 980 10052 990 10108
rect 1046 10071 1132 10108
rect 980 10019 1001 10052
rect 1053 10019 1125 10071
rect 1188 10052 1198 10108
rect 1177 10019 1198 10052
rect 980 9966 1198 10019
rect 980 9910 990 9966
rect 1046 9947 1132 9966
rect 980 9895 1001 9910
rect 1053 9895 1125 9947
rect 1188 9910 1198 9966
rect 1177 9895 1198 9910
rect 980 9824 1198 9895
rect 980 9768 990 9824
rect 1046 9823 1132 9824
rect 1053 9771 1125 9823
rect 1046 9768 1132 9771
rect 1188 9768 1198 9824
rect 980 9758 1198 9768
rect 753 9510 1206 9539
rect 753 9458 1038 9510
rect 1194 9458 1206 9510
rect 753 9431 1206 9458
rect 573 9344 1206 9371
rect 573 9292 1038 9344
rect 1194 9292 1206 9344
rect 573 9271 1206 9292
rect 393 9184 1206 9211
rect 393 9132 1038 9184
rect 1194 9132 1206 9184
rect 393 9111 1206 9132
rect 213 9018 1206 9051
rect 213 8966 1038 9018
rect 1194 8966 1206 9018
rect 213 8951 1206 8966
rect 1313 8943 12165 12658
rect 12298 10818 12516 10828
rect 12298 10762 12308 10818
rect 12364 10815 12450 10818
rect 12371 10763 12443 10815
rect 12364 10762 12450 10763
rect 12506 10762 12516 10818
rect 12298 10691 12516 10762
rect 12298 10676 12319 10691
rect 12298 10620 12308 10676
rect 12371 10639 12443 10691
rect 12495 10676 12516 10691
rect 12364 10620 12450 10639
rect 12506 10620 12516 10676
rect 12298 10567 12516 10620
rect 12298 10534 12319 10567
rect 12298 10478 12308 10534
rect 12371 10515 12443 10567
rect 12495 10534 12516 10567
rect 12364 10478 12450 10515
rect 12506 10478 12516 10534
rect 12298 10443 12516 10478
rect 12298 10392 12319 10443
rect 12298 10336 12308 10392
rect 12371 10391 12443 10443
rect 12495 10392 12516 10443
rect 12364 10336 12450 10391
rect 12506 10336 12516 10392
rect 12298 10319 12516 10336
rect 12298 10267 12319 10319
rect 12371 10267 12443 10319
rect 12495 10267 12516 10319
rect 12298 10250 12516 10267
rect 12298 10194 12308 10250
rect 12364 10195 12450 10250
rect 12298 10143 12319 10194
rect 12371 10143 12443 10195
rect 12506 10194 12516 10250
rect 12495 10143 12516 10194
rect 12298 10108 12516 10143
rect 12298 10052 12308 10108
rect 12364 10071 12450 10108
rect 12298 10019 12319 10052
rect 12371 10019 12443 10071
rect 12506 10052 12516 10108
rect 12495 10019 12516 10052
rect 12298 9966 12516 10019
rect 12298 9910 12308 9966
rect 12364 9947 12450 9966
rect 12298 9895 12319 9910
rect 12371 9895 12443 9947
rect 12506 9910 12516 9966
rect 12495 9895 12516 9910
rect 12298 9824 12516 9895
rect 12298 9768 12308 9824
rect 12364 9823 12450 9824
rect 12371 9771 12443 9823
rect 12364 9768 12450 9771
rect 12506 9768 12516 9824
rect 12298 9758 12516 9768
rect 12617 9539 12725 26936
rect 12305 9510 12725 9539
rect 12305 9458 12317 9510
rect 12473 9458 12725 9510
rect 12305 9431 12725 9458
rect 12805 9371 12905 26936
rect 12305 9344 12905 9371
rect 12305 9292 12317 9344
rect 12473 9292 12905 9344
rect 12305 9271 12905 9292
rect 12985 9211 13085 26936
rect 12305 9184 13085 9211
rect 12305 9132 12317 9184
rect 12473 9132 13085 9184
rect 12305 9111 13085 9132
rect 13165 9051 13265 26936
rect 13408 10818 13768 10828
rect 13408 10762 13418 10818
rect 13474 10764 13560 10818
rect 13616 10764 13702 10818
rect 13758 10762 13768 10818
rect 13408 10676 13462 10762
rect 13722 10676 13768 10762
rect 13408 10620 13418 10676
rect 13758 10620 13768 10676
rect 13408 10534 13462 10620
rect 13722 10534 13768 10620
rect 13408 10478 13418 10534
rect 13758 10478 13768 10534
rect 13408 10392 13462 10478
rect 13722 10392 13768 10478
rect 13408 10336 13418 10392
rect 13758 10336 13768 10392
rect 13408 10250 13462 10336
rect 13722 10250 13768 10336
rect 13408 10194 13418 10250
rect 13758 10194 13768 10250
rect 13408 10108 13462 10194
rect 13722 10108 13768 10194
rect 13408 10052 13418 10108
rect 13758 10052 13768 10108
rect 13408 9966 13462 10052
rect 13722 9966 13768 10052
rect 13408 9910 13418 9966
rect 13758 9910 13768 9966
rect 13408 9824 13462 9910
rect 13722 9824 13768 9910
rect 13408 9768 13418 9824
rect 13474 9768 13560 9776
rect 13616 9768 13702 9776
rect 13758 9768 13768 9824
rect 13408 9758 13768 9768
rect 12305 9018 13265 9051
rect 12305 8966 12317 9018
rect 12473 8966 13265 9018
rect 12305 8951 13265 8966
rect 1313 -1210 1663 8943
rect 1741 8819 2142 8863
rect 1741 8504 1753 8819
rect 1805 8504 2142 8819
rect 1741 6888 1751 8504
rect 1807 6888 2142 8504
rect 1741 6583 1753 6888
rect 1805 6583 2142 6888
rect 1741 6273 2142 6583
rect 1741 5902 1753 6273
rect 1805 5902 2142 6273
rect 1741 3766 1751 5902
rect 1807 3766 2142 5902
rect 1741 3413 1753 3766
rect 1805 3413 2142 3766
rect 1741 3086 2142 3413
rect 1741 2691 1753 3086
rect 1805 2691 2142 3086
rect 1741 971 1751 2691
rect 1807 971 2142 2691
rect 1741 538 1753 971
rect 1805 538 2142 971
rect 1741 510 2142 538
rect 2372 -1210 4016 8943
rect 4720 -1210 6364 8943
rect 7069 -1210 8713 8943
rect 9416 -1210 11060 8943
rect 11290 8819 11732 8863
rect 11290 8504 11627 8819
rect 11679 8504 11732 8819
rect 11290 6888 11625 8504
rect 11681 6888 11732 8504
rect 11290 6583 11627 6888
rect 11679 6583 11732 6888
rect 11290 6273 11732 6583
rect 11290 5902 11627 6273
rect 11679 5902 11732 6273
rect 11290 3766 11625 5902
rect 11681 3766 11732 5902
rect 11290 3413 11627 3766
rect 11679 3413 11732 3766
rect 11290 3086 11732 3413
rect 11290 2691 11627 3086
rect 11679 2691 11732 3086
rect 11290 971 11625 2691
rect 11681 971 11732 2691
rect 11290 538 11627 971
rect 11679 538 11732 971
rect 11290 510 11732 538
rect 11831 -1465 12165 8943
<< via2 >>
rect -316 10764 -260 10818
rect -174 10764 -118 10818
rect -32 10764 24 10818
rect -316 10762 -280 10764
rect -280 10762 -260 10764
rect -174 10762 -118 10764
rect -32 10762 -20 10764
rect -20 10762 24 10764
rect -316 10620 -280 10676
rect -280 10620 -260 10676
rect -174 10620 -118 10676
rect -32 10620 -20 10676
rect -20 10620 24 10676
rect -316 10478 -280 10534
rect -280 10478 -260 10534
rect -174 10478 -118 10534
rect -32 10478 -20 10534
rect -20 10478 24 10534
rect -316 10336 -280 10392
rect -280 10336 -260 10392
rect -174 10336 -118 10392
rect -32 10336 -20 10392
rect -20 10336 24 10392
rect -316 10194 -280 10250
rect -280 10194 -260 10250
rect -174 10194 -118 10250
rect -32 10194 -20 10250
rect -20 10194 24 10250
rect -316 10052 -280 10108
rect -280 10052 -260 10108
rect -174 10052 -118 10108
rect -32 10052 -20 10108
rect -20 10052 24 10108
rect -316 9910 -280 9966
rect -280 9910 -260 9966
rect -174 9910 -118 9966
rect -32 9910 -20 9966
rect -20 9910 24 9966
rect -316 9776 -280 9824
rect -280 9776 -260 9824
rect -174 9776 -118 9824
rect -32 9776 -20 9824
rect -20 9776 24 9824
rect -316 9768 -260 9776
rect -174 9768 -118 9776
rect -32 9768 24 9776
rect 990 10815 1046 10818
rect 1132 10815 1188 10818
rect 990 10763 1001 10815
rect 1001 10763 1046 10815
rect 1132 10763 1177 10815
rect 1177 10763 1188 10815
rect 990 10762 1046 10763
rect 1132 10762 1188 10763
rect 990 10639 1001 10676
rect 1001 10639 1046 10676
rect 1132 10639 1177 10676
rect 1177 10639 1188 10676
rect 990 10620 1046 10639
rect 1132 10620 1188 10639
rect 990 10515 1001 10534
rect 1001 10515 1046 10534
rect 1132 10515 1177 10534
rect 1177 10515 1188 10534
rect 990 10478 1046 10515
rect 1132 10478 1188 10515
rect 990 10391 1001 10392
rect 1001 10391 1046 10392
rect 1132 10391 1177 10392
rect 1177 10391 1188 10392
rect 990 10336 1046 10391
rect 1132 10336 1188 10391
rect 990 10195 1046 10250
rect 1132 10195 1188 10250
rect 990 10194 1001 10195
rect 1001 10194 1046 10195
rect 1132 10194 1177 10195
rect 1177 10194 1188 10195
rect 990 10071 1046 10108
rect 1132 10071 1188 10108
rect 990 10052 1001 10071
rect 1001 10052 1046 10071
rect 1132 10052 1177 10071
rect 1177 10052 1188 10071
rect 990 9947 1046 9966
rect 1132 9947 1188 9966
rect 990 9910 1001 9947
rect 1001 9910 1046 9947
rect 1132 9910 1177 9947
rect 1177 9910 1188 9947
rect 990 9823 1046 9824
rect 1132 9823 1188 9824
rect 990 9771 1001 9823
rect 1001 9771 1046 9823
rect 1132 9771 1177 9823
rect 1177 9771 1188 9823
rect 990 9768 1046 9771
rect 1132 9768 1188 9771
rect 12308 10815 12364 10818
rect 12450 10815 12506 10818
rect 12308 10763 12319 10815
rect 12319 10763 12364 10815
rect 12450 10763 12495 10815
rect 12495 10763 12506 10815
rect 12308 10762 12364 10763
rect 12450 10762 12506 10763
rect 12308 10639 12319 10676
rect 12319 10639 12364 10676
rect 12450 10639 12495 10676
rect 12495 10639 12506 10676
rect 12308 10620 12364 10639
rect 12450 10620 12506 10639
rect 12308 10515 12319 10534
rect 12319 10515 12364 10534
rect 12450 10515 12495 10534
rect 12495 10515 12506 10534
rect 12308 10478 12364 10515
rect 12450 10478 12506 10515
rect 12308 10391 12319 10392
rect 12319 10391 12364 10392
rect 12450 10391 12495 10392
rect 12495 10391 12506 10392
rect 12308 10336 12364 10391
rect 12450 10336 12506 10391
rect 12308 10195 12364 10250
rect 12450 10195 12506 10250
rect 12308 10194 12319 10195
rect 12319 10194 12364 10195
rect 12450 10194 12495 10195
rect 12495 10194 12506 10195
rect 12308 10071 12364 10108
rect 12450 10071 12506 10108
rect 12308 10052 12319 10071
rect 12319 10052 12364 10071
rect 12450 10052 12495 10071
rect 12495 10052 12506 10071
rect 12308 9947 12364 9966
rect 12450 9947 12506 9966
rect 12308 9910 12319 9947
rect 12319 9910 12364 9947
rect 12450 9910 12495 9947
rect 12495 9910 12506 9947
rect 12308 9823 12364 9824
rect 12450 9823 12506 9824
rect 12308 9771 12319 9823
rect 12319 9771 12364 9823
rect 12450 9771 12495 9823
rect 12495 9771 12506 9823
rect 12308 9768 12364 9771
rect 12450 9768 12506 9771
rect 13418 10764 13474 10818
rect 13560 10764 13616 10818
rect 13702 10764 13758 10818
rect 13418 10762 13462 10764
rect 13462 10762 13474 10764
rect 13560 10762 13616 10764
rect 13702 10762 13722 10764
rect 13722 10762 13758 10764
rect 13418 10620 13462 10676
rect 13462 10620 13474 10676
rect 13560 10620 13616 10676
rect 13702 10620 13722 10676
rect 13722 10620 13758 10676
rect 13418 10478 13462 10534
rect 13462 10478 13474 10534
rect 13560 10478 13616 10534
rect 13702 10478 13722 10534
rect 13722 10478 13758 10534
rect 13418 10336 13462 10392
rect 13462 10336 13474 10392
rect 13560 10336 13616 10392
rect 13702 10336 13722 10392
rect 13722 10336 13758 10392
rect 13418 10194 13462 10250
rect 13462 10194 13474 10250
rect 13560 10194 13616 10250
rect 13702 10194 13722 10250
rect 13722 10194 13758 10250
rect 13418 10052 13462 10108
rect 13462 10052 13474 10108
rect 13560 10052 13616 10108
rect 13702 10052 13722 10108
rect 13722 10052 13758 10108
rect 13418 9910 13462 9966
rect 13462 9910 13474 9966
rect 13560 9910 13616 9966
rect 13702 9910 13722 9966
rect 13722 9910 13758 9966
rect 13418 9776 13462 9824
rect 13462 9776 13474 9824
rect 13560 9776 13616 9824
rect 13702 9776 13722 9824
rect 13722 9776 13758 9824
rect 13418 9768 13474 9776
rect 13560 9768 13616 9776
rect 13702 9768 13758 9776
rect 1751 6888 1753 8504
rect 1753 6888 1805 8504
rect 1805 6888 1807 8504
rect 1751 3766 1753 5902
rect 1753 3766 1805 5902
rect 1805 3766 1807 5902
rect 1751 971 1753 2691
rect 1753 971 1805 2691
rect 1805 971 1807 2691
rect 11625 6888 11627 8504
rect 11627 6888 11679 8504
rect 11679 6888 11681 8504
rect 11625 3766 11627 5902
rect 11627 3766 11679 5902
rect 11679 3766 11681 5902
rect 11625 971 11627 2691
rect 11627 971 11679 2691
rect 11679 971 11681 2691
<< metal3 >>
rect -326 10818 34 10828
rect -326 10762 -316 10818
rect -260 10762 -174 10818
rect -118 10762 -32 10818
rect 24 10762 34 10818
rect -326 10676 34 10762
rect -326 10620 -316 10676
rect -260 10620 -174 10676
rect -118 10620 -32 10676
rect 24 10620 34 10676
rect -326 10534 34 10620
rect -326 10478 -316 10534
rect -260 10478 -174 10534
rect -118 10478 -32 10534
rect 24 10478 34 10534
rect -326 10392 34 10478
rect -326 10336 -316 10392
rect -260 10336 -174 10392
rect -118 10336 -32 10392
rect 24 10336 34 10392
rect -326 10250 34 10336
rect -326 10194 -316 10250
rect -260 10194 -174 10250
rect -118 10194 -32 10250
rect 24 10194 34 10250
rect -326 10108 34 10194
rect -326 10052 -316 10108
rect -260 10052 -174 10108
rect -118 10052 -32 10108
rect 24 10052 34 10108
rect -326 9966 34 10052
rect -326 9910 -316 9966
rect -260 9910 -174 9966
rect -118 9910 -32 9966
rect 24 9910 34 9966
rect -326 9824 34 9910
rect -326 9768 -316 9824
rect -260 9768 -174 9824
rect -118 9768 -32 9824
rect 24 9768 34 9824
rect -326 9758 34 9768
rect 980 10818 1198 10828
rect 980 10762 990 10818
rect 1046 10762 1132 10818
rect 1188 10762 1198 10818
rect 980 10676 1198 10762
rect 980 10620 990 10676
rect 1046 10620 1132 10676
rect 1188 10620 1198 10676
rect 980 10534 1198 10620
rect 980 10478 990 10534
rect 1046 10478 1132 10534
rect 1188 10478 1198 10534
rect 980 10392 1198 10478
rect 980 10336 990 10392
rect 1046 10336 1132 10392
rect 1188 10336 1198 10392
rect 980 10250 1198 10336
rect 980 10194 990 10250
rect 1046 10194 1132 10250
rect 1188 10194 1198 10250
rect 980 10108 1198 10194
rect 980 10052 990 10108
rect 1046 10052 1132 10108
rect 1188 10052 1198 10108
rect 980 9966 1198 10052
rect 980 9910 990 9966
rect 1046 9910 1132 9966
rect 1188 9910 1198 9966
rect 980 9824 1198 9910
rect 980 9768 990 9824
rect 1046 9768 1132 9824
rect 1188 9768 1198 9824
rect 980 9758 1198 9768
rect 12298 10818 12516 10828
rect 12298 10762 12308 10818
rect 12364 10762 12450 10818
rect 12506 10762 12516 10818
rect 12298 10676 12516 10762
rect 12298 10620 12308 10676
rect 12364 10620 12450 10676
rect 12506 10620 12516 10676
rect 12298 10534 12516 10620
rect 12298 10478 12308 10534
rect 12364 10478 12450 10534
rect 12506 10478 12516 10534
rect 12298 10392 12516 10478
rect 12298 10336 12308 10392
rect 12364 10336 12450 10392
rect 12506 10336 12516 10392
rect 12298 10250 12516 10336
rect 12298 10194 12308 10250
rect 12364 10194 12450 10250
rect 12506 10194 12516 10250
rect 12298 10108 12516 10194
rect 12298 10052 12308 10108
rect 12364 10052 12450 10108
rect 12506 10052 12516 10108
rect 12298 9966 12516 10052
rect 12298 9910 12308 9966
rect 12364 9910 12450 9966
rect 12506 9910 12516 9966
rect 12298 9824 12516 9910
rect 12298 9768 12308 9824
rect 12364 9768 12450 9824
rect 12506 9768 12516 9824
rect 12298 9758 12516 9768
rect 13408 10818 13768 10828
rect 13408 10762 13418 10818
rect 13474 10762 13560 10818
rect 13616 10762 13702 10818
rect 13758 10762 13768 10818
rect 13408 10676 13768 10762
rect 13408 10620 13418 10676
rect 13474 10620 13560 10676
rect 13616 10620 13702 10676
rect 13758 10620 13768 10676
rect 13408 10534 13768 10620
rect 13408 10478 13418 10534
rect 13474 10478 13560 10534
rect 13616 10478 13702 10534
rect 13758 10478 13768 10534
rect 13408 10392 13768 10478
rect 13408 10336 13418 10392
rect 13474 10336 13560 10392
rect 13616 10336 13702 10392
rect 13758 10336 13768 10392
rect 13408 10250 13768 10336
rect 13408 10194 13418 10250
rect 13474 10194 13560 10250
rect 13616 10194 13702 10250
rect 13758 10194 13768 10250
rect 13408 10108 13768 10194
rect 13408 10052 13418 10108
rect 13474 10052 13560 10108
rect 13616 10052 13702 10108
rect 13758 10052 13768 10108
rect 13408 9966 13768 10052
rect 13408 9910 13418 9966
rect 13474 9910 13560 9966
rect 13616 9910 13702 9966
rect 13758 9910 13768 9966
rect 13408 9824 13768 9910
rect 13408 9768 13418 9824
rect 13474 9768 13560 9824
rect 13616 9768 13702 9824
rect 13758 9768 13768 9824
rect 13408 9758 13768 9768
rect 1741 8504 1817 8514
rect 1741 6888 1751 8504
rect 1807 6888 1817 8504
rect 1741 6878 1817 6888
rect 11615 8504 11691 8514
rect 11615 6888 11625 8504
rect 11681 6888 11691 8504
rect 11615 6878 11691 6888
rect 1741 5902 1817 5912
rect 1741 3766 1751 5902
rect 1807 3766 1817 5902
rect 1741 3756 1817 3766
rect 11615 5902 11691 5912
rect 11615 3766 11625 5902
rect 11681 3766 11691 5902
rect 11615 3756 11691 3766
rect 1741 2691 1817 2701
rect 1741 971 1751 2691
rect 1807 971 1817 2691
rect 1741 961 1817 971
rect 11615 2691 11691 2701
rect 11615 971 11625 2691
rect 11681 971 11691 2691
rect 11615 961 11691 971
use comp018green_out_paddrv_4T_NMOS_GROUP  comp018green_out_paddrv_4T_NMOS_GROUP_0
timestamp 1749760379
transform 1 0 1339 0 1 31
box -1367 -147 12129 10917
use comp018green_out_paddrv_4T_PMOS_GROUP  comp018green_out_paddrv_4T_PMOS_GROUP_0
timestamp 1749760379
transform 1 0 548 0 1 12347
box -767 -1312 13147 15294
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_0
timestamp 1749760379
transform 0 1 12395 1 0 9484
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_1
timestamp 1749760379
transform 0 1 12395 1 0 9318
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_2
timestamp 1749760379
transform 0 1 12395 1 0 9158
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_3
timestamp 1749760379
transform 0 1 12395 1 0 8992
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_4
timestamp 1749760379
transform 0 -1 1116 1 0 9484
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_5
timestamp 1749760379
transform 0 -1 1116 1 0 8992
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_6
timestamp 1749760379
transform 0 -1 1116 1 0 9158
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_7
timestamp 1749760379
transform 0 -1 1116 1 0 9318
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_0
timestamp 1749760379
transform -1 0 11653 0 1 7701
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_1
timestamp 1749760379
transform 1 0 1779 0 1 7701
box 0 0 1 1
use M2_M1_CDNS_40661953145279  M2_M1_CDNS_40661953145279_0
timestamp 1749760379
transform -1 0 11653 0 1 4843
box 0 0 1 1
use M2_M1_CDNS_40661953145279  M2_M1_CDNS_40661953145279_1
timestamp 1749760379
transform 1 0 1779 0 1 4843
box 0 0 1 1
use M2_M1_CDNS_40661953145280  M2_M1_CDNS_40661953145280_0
timestamp 1749760379
transform -1 0 11653 0 1 1812
box 0 0 1 1
use M2_M1_CDNS_40661953145280  M2_M1_CDNS_40661953145280_1
timestamp 1749760379
transform 1 0 1779 0 1 1812
box 0 0 1 1
use M2_M1_CDNS_40661953145343  M2_M1_CDNS_40661953145343_0
timestamp 1749760379
transform 1 0 12407 0 1 10293
box 0 0 1 1
use M2_M1_CDNS_40661953145343  M2_M1_CDNS_40661953145343_1
timestamp 1749760379
transform 1 0 1089 0 1 10293
box 0 0 1 1
use M2_M1_CDNS_40661953145344  M2_M1_CDNS_40661953145344_0
timestamp 1749760379
transform -1 0 13592 0 1 10270
box 0 0 1 1
use M2_M1_CDNS_40661953145344  M2_M1_CDNS_40661953145344_1
timestamp 1749760379
transform 1 0 -150 0 1 10270
box 0 0 1 1
use M3_M2_CDNS_40661953145263  M3_M2_CDNS_40661953145263_0
timestamp 1749760379
transform -1 0 13588 0 1 10293
box 0 0 1 1
use M3_M2_CDNS_40661953145263  M3_M2_CDNS_40661953145263_1
timestamp 1749760379
transform 1 0 -146 0 1 10293
box 0 0 1 1
use M3_M2_CDNS_40661953145278  M3_M2_CDNS_40661953145278_0
timestamp 1749760379
transform 1 0 12407 0 1 10293
box 0 0 1 1
use M3_M2_CDNS_40661953145278  M3_M2_CDNS_40661953145278_1
timestamp 1749760379
transform 1 0 1089 0 1 10293
box 0 0 1 1
use M3_M2_CDNS_40661953145340  M3_M2_CDNS_40661953145340_0
timestamp 1749760379
transform -1 0 11653 0 1 7696
box 0 0 1 1
use M3_M2_CDNS_40661953145340  M3_M2_CDNS_40661953145340_1
timestamp 1749760379
transform 1 0 1779 0 1 7696
box 0 0 1 1
use M3_M2_CDNS_40661953145341  M3_M2_CDNS_40661953145341_0
timestamp 1749760379
transform -1 0 11653 0 1 4834
box 0 0 1 1
use M3_M2_CDNS_40661953145341  M3_M2_CDNS_40661953145341_1
timestamp 1749760379
transform 1 0 1779 0 1 4834
box 0 0 1 1
use M3_M2_CDNS_40661953145342  M3_M2_CDNS_40661953145342_0
timestamp 1749760379
transform -1 0 11653 0 1 1831
box 0 0 1 1
use M3_M2_CDNS_40661953145342  M3_M2_CDNS_40661953145342_1
timestamp 1749760379
transform 1 0 1779 0 1 1831
box 0 0 1 1
<< properties >>
string GDS_END 3554048
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 3548770
string path 42.425 657.500 294.525 657.500 
<< end >>
