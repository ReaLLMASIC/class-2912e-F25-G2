magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 453 2438 1094
<< pwell >>
rect -86 -86 2438 453
<< mvnmos >>
rect 128 69 248 333
rect 352 69 472 333
rect 576 69 696 333
rect 760 69 880 333
rect 1128 69 1248 333
rect 1352 69 1472 333
rect 1576 69 1696 333
rect 1848 69 1968 333
rect 2072 69 2192 333
<< mvpmos >>
rect 138 573 238 939
rect 362 573 462 939
rect 576 573 676 939
rect 780 573 880 939
rect 1148 573 1248 939
rect 1362 573 1462 939
rect 1576 573 1676 939
rect 1868 573 1968 939
rect 2082 573 2182 939
<< mvndiff >>
rect 40 305 128 333
rect 40 165 53 305
rect 99 165 128 305
rect 40 69 128 165
rect 248 305 352 333
rect 248 165 277 305
rect 323 165 352 305
rect 248 69 352 165
rect 472 305 576 333
rect 472 165 501 305
rect 547 165 576 305
rect 472 69 576 165
rect 696 69 760 333
rect 880 305 968 333
rect 880 165 909 305
rect 955 165 968 305
rect 880 69 968 165
rect 1040 305 1128 333
rect 1040 165 1053 305
rect 1099 165 1128 305
rect 1040 69 1128 165
rect 1248 285 1352 333
rect 1248 239 1277 285
rect 1323 239 1352 285
rect 1248 69 1352 239
rect 1472 211 1576 333
rect 1472 165 1501 211
rect 1547 165 1576 211
rect 1472 69 1576 165
rect 1696 305 1848 333
rect 1696 165 1773 305
rect 1819 165 1848 305
rect 1696 69 1848 165
rect 1968 305 2072 333
rect 1968 165 1997 305
rect 2043 165 2072 305
rect 1968 69 2072 165
rect 2192 305 2280 333
rect 2192 165 2221 305
rect 2267 165 2280 305
rect 2192 69 2280 165
<< mvpdiff >>
rect 50 926 138 939
rect 50 786 63 926
rect 109 786 138 926
rect 50 573 138 786
rect 238 860 362 939
rect 238 720 277 860
rect 323 720 362 860
rect 238 573 362 720
rect 462 926 576 939
rect 462 786 491 926
rect 537 786 576 926
rect 462 573 576 786
rect 676 854 780 939
rect 676 714 705 854
rect 751 714 780 854
rect 676 573 780 714
rect 880 926 968 939
rect 880 786 909 926
rect 955 786 968 926
rect 880 573 968 786
rect 1060 926 1148 939
rect 1060 786 1073 926
rect 1119 786 1148 926
rect 1060 573 1148 786
rect 1248 573 1362 939
rect 1462 832 1576 939
rect 1462 786 1501 832
rect 1547 786 1576 832
rect 1462 573 1576 786
rect 1676 926 1868 939
rect 1676 786 1773 926
rect 1819 786 1868 926
rect 1676 573 1868 786
rect 1968 860 2082 939
rect 1968 720 1997 860
rect 2043 720 2082 860
rect 1968 573 2082 720
rect 2182 926 2270 939
rect 2182 786 2211 926
rect 2257 786 2270 926
rect 2182 573 2270 786
<< mvndiffc >>
rect 53 165 99 305
rect 277 165 323 305
rect 501 165 547 305
rect 909 165 955 305
rect 1053 165 1099 305
rect 1277 239 1323 285
rect 1501 165 1547 211
rect 1773 165 1819 305
rect 1997 165 2043 305
rect 2221 165 2267 305
<< mvpdiffc >>
rect 63 786 109 926
rect 277 720 323 860
rect 491 786 537 926
rect 705 714 751 854
rect 909 786 955 926
rect 1073 786 1119 926
rect 1501 786 1547 832
rect 1773 786 1819 926
rect 1997 720 2043 860
rect 2211 786 2257 926
<< polysilicon >>
rect 138 939 238 983
rect 362 939 462 983
rect 576 939 676 983
rect 780 939 880 983
rect 1148 939 1248 983
rect 1362 939 1462 983
rect 1576 939 1676 983
rect 1868 939 1968 983
rect 2082 939 2182 983
rect 138 513 238 573
rect 362 522 462 573
rect 362 513 403 522
rect 138 441 403 513
rect 138 377 248 441
rect 128 333 248 377
rect 352 382 403 441
rect 449 382 462 522
rect 352 377 462 382
rect 576 500 676 573
rect 576 454 617 500
rect 663 454 676 500
rect 576 377 676 454
rect 780 513 880 573
rect 1148 513 1248 573
rect 780 500 1248 513
rect 780 454 814 500
rect 860 454 1248 500
rect 780 441 1248 454
rect 780 377 880 441
rect 352 333 472 377
rect 576 333 696 377
rect 760 333 880 377
rect 1128 333 1248 441
rect 1362 500 1462 573
rect 1362 454 1375 500
rect 1421 454 1462 500
rect 1362 377 1462 454
rect 1576 529 1676 573
rect 1576 389 1589 529
rect 1635 389 1676 529
rect 1576 377 1676 389
rect 1868 518 1968 573
rect 1868 378 1881 518
rect 1927 513 1968 518
rect 2082 513 2182 573
rect 1927 441 2182 513
rect 1927 378 1968 441
rect 1868 377 1968 378
rect 1352 333 1472 377
rect 1576 333 1696 377
rect 1848 333 1968 377
rect 2072 377 2182 441
rect 2072 333 2192 377
rect 128 25 248 69
rect 352 25 472 69
rect 576 25 696 69
rect 760 25 880 69
rect 1128 25 1248 69
rect 1352 25 1472 69
rect 1576 25 1696 69
rect 1848 25 1968 69
rect 2072 25 2192 69
<< polycontact >>
rect 403 382 449 522
rect 617 454 663 500
rect 814 454 860 500
rect 1375 454 1421 500
rect 1589 389 1635 529
rect 1881 378 1927 518
<< metal1 >>
rect 0 926 2352 1098
rect 0 918 63 926
rect 109 918 491 926
rect 63 775 109 786
rect 254 860 323 871
rect 254 720 277 860
rect 537 918 909 926
rect 491 775 537 786
rect 705 854 751 865
rect 53 305 99 316
rect 53 90 99 165
rect 254 305 323 720
rect 514 714 705 726
rect 955 918 1073 926
rect 909 775 955 786
rect 1119 918 1773 926
rect 1073 775 1119 786
rect 1501 832 1727 843
rect 1547 786 1727 832
rect 1501 775 1727 786
rect 1819 918 2211 926
rect 1773 775 1819 786
rect 1997 860 2043 871
rect 751 714 1635 726
rect 514 680 1635 714
rect 514 533 560 680
rect 403 522 560 533
rect 449 477 560 522
rect 722 588 1202 634
rect 722 500 768 588
rect 606 454 617 500
rect 663 454 768 500
rect 814 500 866 542
rect 860 454 866 500
rect 1150 500 1202 588
rect 1589 529 1635 680
rect 1150 454 1375 500
rect 1421 454 1432 500
rect 814 430 866 454
rect 403 371 449 382
rect 909 389 1589 408
rect 909 362 1635 389
rect 1681 529 1727 775
rect 2257 918 2352 926
rect 2211 775 2257 786
rect 1681 518 1927 529
rect 1681 454 1881 518
rect 254 165 277 305
rect 254 154 323 165
rect 501 305 547 316
rect 501 90 547 165
rect 909 305 955 362
rect 909 154 955 165
rect 1053 305 1099 316
rect 1681 314 1727 454
rect 1880 378 1881 454
rect 1880 367 1927 378
rect 1997 318 2043 720
rect 1277 285 1727 314
rect 1323 268 1727 285
rect 1773 305 1819 316
rect 1277 228 1323 239
rect 1501 211 1547 222
rect 1099 165 1501 182
rect 1053 136 1547 165
rect 1773 90 1819 165
rect 1997 305 2098 318
rect 2043 165 2098 305
rect 1997 154 2098 165
rect 2221 305 2267 316
rect 2221 90 2267 165
rect 0 -90 2352 90
<< labels >>
flabel metal1 s 722 588 1202 634 0 FreeSans 200 0 0 0 A
port 1 nsew default input
flabel metal1 s 814 430 866 542 0 FreeSans 200 0 0 0 B
port 2 nsew default input
flabel metal1 s 254 154 323 871 0 FreeSans 200 0 0 0 CO
port 3 nsew default output
flabel metal1 s 1997 318 2043 871 0 FreeSans 200 0 0 0 S
port 4 nsew default output
flabel metal1 s 0 918 2352 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 2221 90 2267 316 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 1150 500 1202 588 1 A
port 1 nsew default input
rlabel metal1 s 722 500 768 588 1 A
port 1 nsew default input
rlabel metal1 s 1150 454 1432 500 1 A
port 1 nsew default input
rlabel metal1 s 606 454 768 500 1 A
port 1 nsew default input
rlabel metal1 s 1997 154 2098 318 1 S
port 4 nsew default output
rlabel metal1 s 2211 775 2257 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1773 775 1819 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1073 775 1119 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 909 775 955 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 491 775 537 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 63 775 109 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1773 90 1819 316 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 501 90 547 316 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 53 90 99 316 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2352 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2352 1008
string GDS_END 1115666
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1109232
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
