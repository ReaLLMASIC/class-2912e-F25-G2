magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect 13512 13500 70089 70434
<< obsm1 >>
rect 13108 13108 71000 71000
<< obsm2 >>
rect 13606 13594 70901 70890
<< metal3 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70800 52400 71000 53800
rect 70800 50800 71000 52200
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70412 42800 70488 45799
rect 70800 41200 71000 42600
rect 70800 39600 71000 41000
rect 70800 36400 71000 39400
rect 70800 33200 71000 36200
rect 70800 30000 71000 33000
rect 70800 26800 71000 29800
rect 70800 25200 71000 26600
rect 70800 23600 71000 25000
rect 70800 20400 71000 23400
rect 70800 17200 71000 20200
rect 70800 14000 71000 17000
<< obsm3 >>
rect 17060 70740 17140 70890
rect 20260 70740 20340 70890
rect 23460 70740 23540 70890
rect 25060 70740 25140 70890
rect 26660 70740 26740 70890
rect 29860 70740 29940 70890
rect 33060 70740 33140 70890
rect 36260 70740 36340 70890
rect 39460 70740 39540 70890
rect 41060 70740 41140 70890
rect 42660 70740 42740 70890
rect 45860 70740 45940 70890
rect 49060 70740 49140 70890
rect 50660 70740 50740 70890
rect 52260 70740 52340 70890
rect 53860 70740 53940 70890
rect 55460 70740 55540 70890
rect 57060 70740 57140 70890
rect 58660 70740 58740 70890
rect 60260 70740 60340 70890
rect 61860 70740 61940 70890
rect 63460 70740 63540 70890
rect 65060 70740 65140 70890
rect 66660 70740 66740 70890
rect 68260 70740 68340 70890
rect 69738 70740 71000 70890
rect 14000 69738 71000 70740
rect 14000 68340 70740 69738
rect 14000 68260 71000 68340
rect 14000 66740 70740 68260
rect 14000 66660 71000 66740
rect 14000 65140 70740 66660
rect 14000 65060 71000 65140
rect 14000 63540 70740 65060
rect 14000 63460 71000 63540
rect 14000 61940 70740 63460
rect 14000 61860 71000 61940
rect 14000 60340 70740 61860
rect 14000 60260 71000 60340
rect 14000 58740 70740 60260
rect 14000 58660 71000 58740
rect 14000 57140 70740 58660
rect 14000 57060 71000 57140
rect 14000 55540 70740 57060
rect 14000 55460 71000 55540
rect 14000 53940 70740 55460
rect 14000 53860 71000 53940
rect 14000 52340 70740 53860
rect 14000 52260 71000 52340
rect 14000 50740 70740 52260
rect 14000 50660 71000 50740
rect 14000 49140 70740 50660
rect 14000 49060 71000 49140
rect 14000 45940 70740 49060
rect 14000 45859 71000 45940
rect 14000 42740 70352 45859
rect 70548 42740 71000 45859
rect 14000 42660 71000 42740
rect 14000 41140 70740 42660
rect 14000 41060 71000 41140
rect 14000 39540 70740 41060
rect 14000 39460 71000 39540
rect 14000 36340 70740 39460
rect 14000 36260 71000 36340
rect 14000 33140 70740 36260
rect 14000 33060 71000 33140
rect 14000 29940 70740 33060
rect 14000 29860 71000 29940
rect 14000 26740 70740 29860
rect 14000 26660 71000 26740
rect 14000 25140 70740 26660
rect 14000 25060 71000 25140
rect 14000 23540 70740 25060
rect 14000 23460 71000 23540
rect 14000 20340 70740 23460
rect 14000 20260 71000 20340
rect 14000 17140 70740 20260
rect 14000 17060 71000 17140
rect 14000 14000 70740 17060
<< metal4 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 34408 70196 34464 70252
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70390 53138 70446 53194
rect 70800 52400 71000 53800
rect 70517 51406 70573 51462
rect 70800 50800 71000 52200
rect 70516 49938 70572 49994
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70412 42800 70488 45799
rect 70800 41200 71000 42600
rect 70800 39600 71000 41000
rect 70800 36400 71000 39400
rect 70800 33200 71000 36200
rect 70800 30000 71000 33000
rect 70800 26800 71000 29800
rect 70800 25200 71000 26600
rect 70800 23600 71000 25000
rect 70800 20400 71000 23400
rect 70800 17200 71000 20200
rect 70800 14000 71000 17000
<< obsm4 >>
rect 17060 70740 17140 70800
rect 20260 70740 20340 70800
rect 23460 70740 23540 70800
rect 25060 70740 25140 70800
rect 26660 70740 26740 70800
rect 29860 70740 29940 70800
rect 33060 70740 33140 70800
rect 36260 70740 36340 70800
rect 39460 70740 39540 70800
rect 41060 70740 41140 70800
rect 42660 70740 42740 70800
rect 45860 70740 45940 70800
rect 49060 70740 49140 70800
rect 50660 70740 50740 70800
rect 52260 70740 52340 70800
rect 53860 70740 53940 70800
rect 55460 70740 55540 70800
rect 57060 70740 57140 70800
rect 58660 70740 58740 70800
rect 60260 70740 60340 70800
rect 61860 70740 61940 70800
rect 63460 70740 63540 70800
rect 65060 70740 65140 70800
rect 66660 70740 66740 70800
rect 68260 70740 68340 70800
rect 69738 70740 71000 70800
rect 14000 70252 71000 70740
rect 14000 70196 34408 70252
rect 34464 70196 71000 70252
rect 14000 69738 71000 70196
rect 14000 68340 70740 69738
rect 14000 68260 71000 68340
rect 14000 66740 70740 68260
rect 14000 66660 71000 66740
rect 14000 65140 70740 66660
rect 14000 65060 71000 65140
rect 14000 63540 70740 65060
rect 14000 63460 71000 63540
rect 14000 61940 70740 63460
rect 14000 61860 71000 61940
rect 14000 60340 70740 61860
rect 14000 60260 71000 60340
rect 14000 58740 70740 60260
rect 14000 58660 71000 58740
rect 14000 57140 70740 58660
rect 14000 57060 71000 57140
rect 14000 55540 70740 57060
rect 14000 55460 71000 55540
rect 14000 53940 70740 55460
rect 14000 53860 71000 53940
rect 14000 53194 70740 53860
rect 14000 53138 70390 53194
rect 70446 53138 70740 53194
rect 14000 52340 70740 53138
rect 14000 52260 71000 52340
rect 14000 51462 70740 52260
rect 14000 51406 70517 51462
rect 70573 51406 70740 51462
rect 14000 50740 70740 51406
rect 14000 50660 71000 50740
rect 14000 49994 70740 50660
rect 14000 49938 70516 49994
rect 70572 49938 70740 49994
rect 14000 49140 70740 49938
rect 14000 49060 71000 49140
rect 14000 45940 70740 49060
rect 14000 45859 71000 45940
rect 14000 42740 70352 45859
rect 70548 42740 71000 45859
rect 14000 42660 71000 42740
rect 14000 41140 70740 42660
rect 14000 41060 71000 41140
rect 14000 39540 70740 41060
rect 14000 39460 71000 39540
rect 14000 36340 70740 39460
rect 14000 36260 71000 36340
rect 14000 33140 70740 36260
rect 14000 33060 71000 33140
rect 14000 29940 70740 33060
rect 14000 29860 71000 29940
rect 14000 26740 70740 29860
rect 14000 26660 71000 26740
rect 14000 25140 70740 26660
rect 14000 25060 71000 25140
rect 14000 23540 70740 25060
rect 14000 23460 71000 23540
rect 14000 20340 70740 23460
rect 14000 20260 71000 20340
rect 14000 17140 70740 20260
rect 14000 17060 71000 17140
rect 14000 14000 70740 17060
<< metal5 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 15396 47287 15472 70800
rect 18596 48623 18672 70800
rect 20400 70151 23400 70227
rect 23600 70160 25000 70236
rect 25200 70164 26600 70240
rect 28064 52629 28140 70800
rect 31264 53967 31340 70800
rect 34408 70196 34464 70252
rect 37664 56640 37740 70800
rect 40262 57314 40338 70800
rect 41862 57986 41938 70800
rect 42800 70148 45800 70224
rect 46000 70171 49000 70247
rect 49200 70176 50600 70252
rect 51462 62015 51538 70800
rect 53062 62683 53138 70800
rect 54662 63349 54738 70800
rect 56262 64012 56338 70800
rect 57862 64675 57938 70800
rect 59462 65342 59538 70800
rect 61062 66007 61138 70800
rect 62662 66670 62738 70800
rect 64262 67342 64338 70800
rect 65867 68000 65943 70800
rect 67462 68669 67538 70800
rect 69001 69258 69077 70800
rect 70395 68400 70471 69678
rect 70800 68400 71000 69678
rect 70402 66800 70478 68200
rect 70800 66800 71000 68200
rect 70400 65200 70476 66600
rect 70800 65200 71000 66600
rect 70399 63600 70475 65000
rect 70800 63600 71000 65000
rect 70393 62000 70469 63400
rect 70800 62000 71000 63400
rect 70391 60400 70467 61800
rect 70800 60400 71000 61800
rect 70389 58800 70465 60200
rect 70800 58800 71000 60200
rect 70386 57200 70462 58600
rect 70800 57200 71000 58600
rect 70384 55600 70460 57000
rect 70800 55600 71000 57000
rect 70382 54000 70458 55400
rect 70800 54000 71000 55400
rect 70390 53138 70446 53194
rect 70800 52400 71000 53800
rect 70517 51406 70573 51462
rect 70800 50800 71000 52200
rect 70516 49938 70572 49994
rect 70800 49200 71000 50600
rect 70800 47604 71000 49000
rect 60617 47528 71000 47604
rect 70800 46000 71000 47528
rect 70412 42800 70488 45799
rect 70407 41200 70483 42600
rect 70800 41200 71000 42600
rect 70401 39600 70477 41000
rect 70800 39600 71000 41000
rect 70394 36400 70470 39400
rect 70800 36400 71000 39400
rect 70384 33200 70460 36200
rect 70800 33200 71000 36200
rect 70800 31604 71000 33000
rect 58681 31528 71000 31604
rect 70800 30000 71000 31528
rect 70800 28404 71000 29800
rect 58681 28328 71000 28404
rect 70800 26800 71000 28328
rect 70800 26070 71000 26600
rect 51296 25994 71000 26070
rect 70800 25200 71000 25994
rect 70424 23600 70500 25000
rect 70800 23600 71000 25000
rect 70415 20400 70491 23400
rect 70800 20400 71000 23400
rect 70800 18936 71000 20200
rect 58405 18860 71000 18936
rect 70800 17200 71000 18860
rect 70404 14000 70480 17000
rect 70800 14000 71000 17000
<< obsm5 >>
rect 14000 47187 15296 70700
rect 15572 48523 18496 70700
rect 18772 70340 27964 70700
rect 18772 70336 25100 70340
rect 18772 70327 23500 70336
rect 18772 70051 20300 70327
rect 26700 70064 27964 70340
rect 25100 70060 27964 70064
rect 23500 70051 27964 70060
rect 18772 52529 27964 70051
rect 28240 53867 31164 70700
rect 31440 70352 37564 70700
rect 31440 70096 34308 70352
rect 34564 70096 37564 70352
rect 31440 56540 37564 70096
rect 37840 57214 40162 70700
rect 40438 57886 41762 70700
rect 42038 70352 51362 70700
rect 42038 70347 49100 70352
rect 42038 70324 45900 70347
rect 42038 70048 42700 70324
rect 50700 70076 51362 70352
rect 49100 70071 51362 70076
rect 45900 70048 51362 70071
rect 42038 61915 51362 70048
rect 51638 62583 52962 70700
rect 53238 63249 54562 70700
rect 54838 63912 56162 70700
rect 56438 64575 57762 70700
rect 58038 65242 59362 70700
rect 59638 65907 60962 70700
rect 61238 66570 62562 70700
rect 62838 67242 64162 70700
rect 64438 67900 65767 70700
rect 66043 68569 67362 70700
rect 67638 69158 68901 70700
rect 69778 70700 71000 70800
rect 69177 69778 71000 70700
rect 69177 69158 70295 69778
rect 67638 68569 70295 69158
rect 66043 68300 70295 68569
rect 70571 68300 70700 69778
rect 66043 67900 70302 68300
rect 64438 67242 70302 67900
rect 62838 66700 70302 67242
rect 70578 66700 70700 68300
rect 62838 66570 70300 66700
rect 61238 65907 70300 66570
rect 59638 65242 70300 65907
rect 58038 65100 70300 65242
rect 70576 65100 70700 66700
rect 58038 64575 70299 65100
rect 56438 63912 70299 64575
rect 54838 63500 70299 63912
rect 70575 63500 70700 65100
rect 54838 63249 70293 63500
rect 53238 62583 70293 63249
rect 51638 61915 70293 62583
rect 42038 61900 70293 61915
rect 70569 61900 70700 63500
rect 42038 60300 70291 61900
rect 70567 60300 70700 61900
rect 42038 58700 70289 60300
rect 70565 58700 70700 60300
rect 42038 57886 70286 58700
rect 40438 57214 70286 57886
rect 37840 57100 70286 57214
rect 70562 57100 70700 58700
rect 37840 56540 70284 57100
rect 31440 55500 70284 56540
rect 70560 55500 70700 57100
rect 31440 53900 70282 55500
rect 70558 53900 70700 55500
rect 31440 53867 70700 53900
rect 28240 53294 70700 53867
rect 28240 53038 70290 53294
rect 70546 53038 70700 53294
rect 28240 52529 70700 53038
rect 18772 51562 70700 52529
rect 18772 51306 70417 51562
rect 70673 51306 70700 51562
rect 18772 50094 70700 51306
rect 18772 49838 70416 50094
rect 70672 49838 70700 50094
rect 18772 48523 70700 49838
rect 15572 47704 70700 48523
rect 15572 47428 60517 47704
rect 15572 47187 70700 47428
rect 14000 45900 70700 47187
rect 14000 45899 71000 45900
rect 14000 42700 70312 45899
rect 70588 42700 71000 45899
rect 14000 41100 70307 42700
rect 70583 41100 70700 42700
rect 14000 39500 70301 41100
rect 70577 39500 70700 41100
rect 14000 36300 70294 39500
rect 70570 36300 70700 39500
rect 14000 33100 70284 36300
rect 70560 33100 70700 36300
rect 14000 31704 70700 33100
rect 14000 31428 58581 31704
rect 14000 28504 70700 31428
rect 14000 28228 58581 28504
rect 14000 26170 70700 28228
rect 14000 25894 51196 26170
rect 14000 25100 70700 25894
rect 14000 23500 70324 25100
rect 70600 23500 70700 25100
rect 14000 20300 70315 23500
rect 70591 20300 70700 23500
rect 14000 19036 70700 20300
rect 14000 18760 58305 19036
rect 14000 17100 70700 18760
rect 14000 14000 70304 17100
rect 70580 14000 70700 17100
<< labels >>
rlabel metal3 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 55600 70800 57000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70412 42800 70488 45799 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 55600 70800 57000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70412 42800 70488 45799 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 55600 70800 57000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 54662 63349 54738 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 67462 68669 67538 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70412 42800 70488 45799 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70390 53138 70446 53194 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70390 53138 70446 53194 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70382 54000 70458 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70384 55600 70460 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70389 58800 70465 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70402 66800 70478 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 42800 70148 45800 70224 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 53062 62683 53138 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 56262 64012 56338 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 59462 65342 59538 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 41862 57986 41938 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 37664 56640 37740 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 23600 70160 25000 70236 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 28064 52629 28140 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 31264 53967 31340 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 34408 70196 34464 70252 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 34408 70196 34464 70252 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70394 36400 70470 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70407 41200 70483 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 58681 31528 70800 31604 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70384 33200 70460 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70424 23600 70500 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 58681 28328 70800 28404 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 69001 69258 69077 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 60617 47528 70800 47604 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70386 57200 70462 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70391 60400 70467 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70400 65200 70476 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70395 68400 70471 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 46000 70171 49000 70247 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 57862 64675 57938 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 61062 66007 61138 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 65867 68000 65943 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 40262 57314 40338 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 15396 47287 15472 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 18596 48623 18672 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 20400 70151 23400 70227 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 25200 70164 26600 70240 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 58405 18860 70800 18936 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70404 14000 70480 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70415 20400 70491 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 51296 25994 70800 26070 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70401 39600 70477 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70517 51406 70573 51462 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70517 51406 70573 51462 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70393 62000 70469 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 51462 62015 51538 70800 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 62662 66670 62738 70800 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70516 49938 70572 49994 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70516 49938 70572 49994 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70399 63600 70475 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 49200 70176 50600 70252 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 64262 67342 64338 70800 6 VSS
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string LEFclass ENDCAP BOTTOMLEFT
string LEFsite GF_COR_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 17524782
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17514044
<< end >>
