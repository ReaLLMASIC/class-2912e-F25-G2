magic
tech gf180mcuD
timestamp 1749760379
<< properties >>
string GDS_END 2756302
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2753866
<< end >>
