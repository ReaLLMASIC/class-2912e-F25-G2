magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 453 5126 1094
<< pwell >>
rect -86 -86 5126 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 978 68 1098 332
rect 1202 68 1322 332
rect 1426 68 1546 332
rect 1650 68 1770 332
rect 1874 68 1994 332
rect 2098 68 2218 332
rect 2322 68 2442 332
rect 2546 68 2666 332
rect 2770 68 2890 332
rect 2994 68 3114 332
rect 3218 68 3338 332
rect 3442 68 3562 332
rect 3666 68 3786 332
rect 3890 68 4010 332
rect 4114 68 4234 332
rect 4338 68 4458 332
rect 4562 68 4682 332
rect 4786 68 4906 332
<< mvpmos >>
rect 172 573 272 933
rect 376 573 476 933
rect 660 573 760 933
rect 1098 580 1198 940
rect 1302 580 1402 940
rect 1506 580 1606 940
rect 1710 580 1810 940
rect 1914 580 2014 940
rect 2118 580 2218 940
rect 2322 580 2422 940
rect 2526 580 2626 940
rect 2730 580 2830 940
rect 2934 580 3034 940
rect 3138 580 3238 940
rect 3342 580 3442 940
rect 3546 580 3646 940
rect 3750 580 3850 940
rect 3954 580 4054 940
rect 4158 580 4258 940
rect 4362 580 4462 940
rect 4566 580 4666 940
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 69 124 274
rect 244 128 348 333
rect 244 82 273 128
rect 319 82 348 128
rect 244 69 348 82
rect 468 287 572 333
rect 468 147 497 287
rect 543 147 572 287
rect 468 69 572 147
rect 692 320 780 333
rect 692 274 721 320
rect 767 274 780 320
rect 692 69 780 274
rect 852 125 978 332
rect 852 79 865 125
rect 911 79 978 125
rect 852 68 978 79
rect 1098 228 1202 332
rect 1098 182 1127 228
rect 1173 182 1202 228
rect 1098 68 1202 182
rect 1322 127 1426 332
rect 1322 81 1351 127
rect 1397 81 1426 127
rect 1322 68 1426 81
rect 1546 287 1650 332
rect 1546 147 1575 287
rect 1621 147 1650 287
rect 1546 68 1650 147
rect 1770 127 1874 332
rect 1770 81 1799 127
rect 1845 81 1874 127
rect 1770 68 1874 81
rect 1994 287 2098 332
rect 1994 147 2023 287
rect 2069 147 2098 287
rect 1994 68 2098 147
rect 2218 127 2322 332
rect 2218 81 2247 127
rect 2293 81 2322 127
rect 2218 68 2322 81
rect 2442 272 2546 332
rect 2442 226 2471 272
rect 2517 226 2546 272
rect 2442 68 2546 226
rect 2666 127 2770 332
rect 2666 81 2695 127
rect 2741 81 2770 127
rect 2666 68 2770 81
rect 2890 319 2994 332
rect 2890 179 2919 319
rect 2965 179 2994 319
rect 2890 68 2994 179
rect 3114 127 3218 332
rect 3114 81 3143 127
rect 3189 81 3218 127
rect 3114 68 3218 81
rect 3338 319 3442 332
rect 3338 179 3367 319
rect 3413 179 3442 319
rect 3338 68 3442 179
rect 3562 127 3666 332
rect 3562 81 3591 127
rect 3637 81 3666 127
rect 3562 68 3666 81
rect 3786 319 3890 332
rect 3786 179 3815 319
rect 3861 179 3890 319
rect 3786 68 3890 179
rect 4010 127 4114 332
rect 4010 81 4039 127
rect 4085 81 4114 127
rect 4010 68 4114 81
rect 4234 319 4338 332
rect 4234 179 4263 319
rect 4309 179 4338 319
rect 4234 68 4338 179
rect 4458 127 4562 332
rect 4458 81 4487 127
rect 4533 81 4562 127
rect 4458 68 4562 81
rect 4682 272 4786 332
rect 4682 226 4711 272
rect 4757 226 4786 272
rect 4682 68 4786 226
rect 4906 221 4994 332
rect 4906 81 4935 221
rect 4981 81 4994 221
rect 4906 68 4994 81
rect 852 66 918 68
<< mvpdiff >>
rect 84 739 172 933
rect 84 599 97 739
rect 143 599 172 739
rect 84 573 172 599
rect 272 920 376 933
rect 272 780 301 920
rect 347 780 376 920
rect 272 573 376 780
rect 476 840 660 933
rect 476 700 585 840
rect 631 700 660 840
rect 476 573 660 700
rect 760 632 848 933
rect 760 586 789 632
rect 835 586 848 632
rect 760 573 848 586
rect 1010 927 1098 940
rect 1010 787 1023 927
rect 1069 787 1098 927
rect 1010 580 1098 787
rect 1198 639 1302 940
rect 1198 593 1227 639
rect 1273 593 1302 639
rect 1198 580 1302 593
rect 1402 927 1506 940
rect 1402 787 1431 927
rect 1477 787 1506 927
rect 1402 580 1506 787
rect 1606 639 1710 940
rect 1606 593 1635 639
rect 1681 593 1710 639
rect 1606 580 1710 593
rect 1810 927 1914 940
rect 1810 787 1839 927
rect 1885 787 1914 927
rect 1810 580 1914 787
rect 2014 777 2118 940
rect 2014 637 2043 777
rect 2089 637 2118 777
rect 2014 580 2118 637
rect 2218 927 2322 940
rect 2218 787 2247 927
rect 2293 787 2322 927
rect 2218 580 2322 787
rect 2422 824 2526 940
rect 2422 684 2451 824
rect 2497 684 2526 824
rect 2422 580 2526 684
rect 2626 927 2730 940
rect 2626 881 2655 927
rect 2701 881 2730 927
rect 2626 580 2730 881
rect 2830 824 2934 940
rect 2830 684 2859 824
rect 2905 684 2934 824
rect 2830 580 2934 684
rect 3034 927 3138 940
rect 3034 881 3063 927
rect 3109 881 3138 927
rect 3034 580 3138 881
rect 3238 824 3342 940
rect 3238 684 3267 824
rect 3313 684 3342 824
rect 3238 580 3342 684
rect 3442 927 3546 940
rect 3442 881 3471 927
rect 3517 881 3546 927
rect 3442 580 3546 881
rect 3646 824 3750 940
rect 3646 684 3675 824
rect 3721 684 3750 824
rect 3646 580 3750 684
rect 3850 927 3954 940
rect 3850 881 3879 927
rect 3925 881 3954 927
rect 3850 580 3954 881
rect 4054 824 4158 940
rect 4054 684 4083 824
rect 4129 684 4158 824
rect 4054 580 4158 684
rect 4258 927 4362 940
rect 4258 881 4287 927
rect 4333 881 4362 927
rect 4258 580 4362 881
rect 4462 824 4566 940
rect 4462 684 4491 824
rect 4537 684 4566 824
rect 4462 580 4566 684
rect 4666 927 4754 940
rect 4666 787 4695 927
rect 4741 787 4754 927
rect 4666 580 4754 787
<< mvndiffc >>
rect 49 274 95 320
rect 273 82 319 128
rect 497 147 543 287
rect 721 274 767 320
rect 865 79 911 125
rect 1127 182 1173 228
rect 1351 81 1397 127
rect 1575 147 1621 287
rect 1799 81 1845 127
rect 2023 147 2069 287
rect 2247 81 2293 127
rect 2471 226 2517 272
rect 2695 81 2741 127
rect 2919 179 2965 319
rect 3143 81 3189 127
rect 3367 179 3413 319
rect 3591 81 3637 127
rect 3815 179 3861 319
rect 4039 81 4085 127
rect 4263 179 4309 319
rect 4487 81 4533 127
rect 4711 226 4757 272
rect 4935 81 4981 221
<< mvpdiffc >>
rect 97 599 143 739
rect 301 780 347 920
rect 585 700 631 840
rect 789 586 835 632
rect 1023 787 1069 927
rect 1227 593 1273 639
rect 1431 787 1477 927
rect 1635 593 1681 639
rect 1839 787 1885 927
rect 2043 637 2089 777
rect 2247 787 2293 927
rect 2451 684 2497 824
rect 2655 881 2701 927
rect 2859 684 2905 824
rect 3063 881 3109 927
rect 3267 684 3313 824
rect 3471 881 3517 927
rect 3675 684 3721 824
rect 3879 881 3925 927
rect 4083 684 4129 824
rect 4287 881 4333 927
rect 4491 684 4537 824
rect 4695 787 4741 927
<< polysilicon >>
rect 172 933 272 977
rect 376 933 476 977
rect 660 933 760 977
rect 1098 940 1198 984
rect 1302 940 1402 984
rect 1506 940 1606 984
rect 1710 940 1810 984
rect 1914 940 2014 984
rect 2118 940 2218 984
rect 2322 940 2422 984
rect 2526 940 2626 984
rect 2730 940 2830 984
rect 2934 940 3034 984
rect 3138 940 3238 984
rect 3342 940 3442 984
rect 3546 940 3646 984
rect 3750 940 3850 984
rect 3954 940 4054 984
rect 4158 940 4258 984
rect 4362 940 4462 984
rect 4566 940 4666 984
rect 172 523 272 573
rect 172 477 185 523
rect 231 513 272 523
rect 376 513 476 573
rect 660 540 760 573
rect 231 477 612 513
rect 660 494 673 540
rect 719 494 760 540
rect 660 481 760 494
rect 1098 520 1198 580
rect 1302 520 1402 580
rect 1506 520 1606 580
rect 1710 520 1810 580
rect 1914 520 2014 580
rect 2118 520 2218 580
rect 172 473 612 477
rect 172 377 244 473
rect 124 333 244 377
rect 348 412 468 425
rect 348 366 361 412
rect 407 366 468 412
rect 348 333 468 366
rect 572 377 612 473
rect 1098 480 2218 520
rect 2322 547 2422 580
rect 2322 501 2363 547
rect 2409 520 2422 547
rect 2526 547 2626 580
rect 2526 520 2552 547
rect 2409 501 2552 520
rect 2598 520 2626 547
rect 2730 547 2830 580
rect 2730 520 2757 547
rect 2598 501 2757 520
rect 2803 520 2830 547
rect 2934 547 3034 580
rect 2934 520 2959 547
rect 2803 501 2959 520
rect 3005 520 3034 547
rect 3138 547 3238 580
rect 3138 520 3163 547
rect 3005 501 3163 520
rect 3209 520 3238 547
rect 3342 547 3442 580
rect 3342 520 3368 547
rect 3209 501 3368 520
rect 3414 520 3442 547
rect 3546 547 3646 580
rect 3546 520 3573 547
rect 3414 501 3573 520
rect 3619 520 3646 547
rect 3750 547 3850 580
rect 3750 520 3778 547
rect 3619 501 3778 520
rect 3824 520 3850 547
rect 3954 547 4054 580
rect 3954 520 3981 547
rect 3824 501 3981 520
rect 4027 520 4054 547
rect 4158 547 4258 580
rect 4158 520 4185 547
rect 4027 501 4185 520
rect 4231 520 4258 547
rect 4362 520 4462 580
rect 4566 520 4666 580
rect 4231 501 4666 520
rect 2322 480 4666 501
rect 1098 432 1322 480
rect 978 414 1322 432
rect 978 392 1238 414
rect 572 333 692 377
rect 978 332 1098 392
rect 1202 368 1238 392
rect 1284 368 1322 414
rect 1202 332 1322 368
rect 1426 411 1546 480
rect 1426 365 1458 411
rect 1504 365 1546 411
rect 1426 332 1546 365
rect 1650 411 1770 480
rect 1650 365 1688 411
rect 1734 365 1770 411
rect 1650 332 1770 365
rect 1874 411 1994 480
rect 1874 365 1912 411
rect 1958 365 1994 411
rect 1874 332 1994 365
rect 2098 411 2218 480
rect 2098 365 2134 411
rect 2180 365 2218 411
rect 2098 332 2218 365
rect 2322 419 4906 432
rect 2322 373 2335 419
rect 2381 392 2581 419
rect 2381 373 2442 392
rect 2322 332 2442 373
rect 2546 373 2581 392
rect 2627 392 2806 419
rect 2627 373 2666 392
rect 2546 332 2666 373
rect 2770 373 2806 392
rect 2852 392 3032 419
rect 2852 373 2890 392
rect 2770 332 2890 373
rect 2994 373 3032 392
rect 3078 392 3255 419
rect 3078 373 3114 392
rect 2994 332 3114 373
rect 3218 373 3255 392
rect 3301 392 3479 419
rect 3301 373 3338 392
rect 3218 332 3338 373
rect 3442 373 3479 392
rect 3525 392 3702 419
rect 3525 373 3562 392
rect 3442 332 3562 373
rect 3666 373 3702 392
rect 3748 392 3927 419
rect 3748 373 3786 392
rect 3666 332 3786 373
rect 3890 373 3927 392
rect 3973 392 4150 419
rect 3973 373 4010 392
rect 3890 332 4010 373
rect 4114 373 4150 392
rect 4196 392 4906 419
rect 4196 373 4234 392
rect 4114 332 4234 373
rect 4338 332 4458 392
rect 4562 332 4682 392
rect 4786 332 4906 392
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 978 24 1098 68
rect 1202 24 1322 68
rect 1426 24 1546 68
rect 1650 24 1770 68
rect 1874 24 1994 68
rect 2098 24 2218 68
rect 2322 24 2442 68
rect 2546 24 2666 68
rect 2770 24 2890 68
rect 2994 24 3114 68
rect 3218 24 3338 68
rect 3442 24 3562 68
rect 3666 24 3786 68
rect 3890 24 4010 68
rect 4114 24 4234 68
rect 4338 24 4458 68
rect 4562 24 4682 68
rect 4786 24 4906 68
<< polycontact >>
rect 185 477 231 523
rect 673 494 719 540
rect 361 366 407 412
rect 2363 501 2409 547
rect 2552 501 2598 547
rect 2757 501 2803 547
rect 2959 501 3005 547
rect 3163 501 3209 547
rect 3368 501 3414 547
rect 3573 501 3619 547
rect 3778 501 3824 547
rect 3981 501 4027 547
rect 4185 501 4231 547
rect 1238 368 1284 414
rect 1458 365 1504 411
rect 1688 365 1734 411
rect 1912 365 1958 411
rect 2134 365 2180 411
rect 2335 373 2381 419
rect 2581 373 2627 419
rect 2806 373 2852 419
rect 3032 373 3078 419
rect 3255 373 3301 419
rect 3479 373 3525 419
rect 3702 373 3748 419
rect 3927 373 3973 419
rect 4150 373 4196 419
<< metal1 >>
rect 0 927 5040 1098
rect 0 920 1023 927
rect 0 918 301 920
rect 347 918 1023 920
rect 301 769 347 780
rect 585 840 631 851
rect 97 739 143 750
rect 1069 918 1431 927
rect 1023 776 1069 787
rect 1477 918 1839 927
rect 1431 776 1477 787
rect 1885 918 2247 927
rect 1839 776 1885 787
rect 2043 777 2089 788
rect 631 700 927 735
rect 585 689 927 700
rect 881 672 927 689
rect 143 599 719 634
rect 97 588 719 599
rect 142 523 315 542
rect 142 477 185 523
rect 231 477 315 523
rect 142 466 315 477
rect 361 412 407 588
rect 673 540 719 588
rect 673 483 719 494
rect 789 632 835 643
rect 789 437 835 586
rect 361 320 407 366
rect 38 274 49 320
rect 95 274 407 320
rect 629 391 835 437
rect 881 639 2043 672
rect 881 593 1227 639
rect 1273 593 1635 639
rect 1681 637 2043 639
rect 2293 918 2655 927
rect 2644 881 2655 918
rect 2701 918 3063 927
rect 2701 881 2712 918
rect 3052 881 3063 918
rect 3109 918 3471 927
rect 3109 881 3120 918
rect 3460 881 3471 918
rect 3517 918 3879 927
rect 3517 881 3528 918
rect 3868 881 3879 918
rect 3925 918 4287 927
rect 3925 881 3936 918
rect 4276 881 4287 918
rect 4333 918 4695 927
rect 4333 881 4344 918
rect 2247 776 2293 787
rect 2451 824 4537 835
rect 2497 684 2859 824
rect 2905 684 3267 824
rect 3313 684 3675 824
rect 3721 684 4083 824
rect 4129 684 4491 824
rect 4741 918 5040 927
rect 4695 776 4741 787
rect 2451 673 4537 684
rect 1681 628 2089 637
rect 1681 593 2339 628
rect 881 582 2339 593
rect 629 298 675 391
rect 881 331 927 582
rect 2293 558 2339 582
rect 2293 547 4242 558
rect 2293 501 2363 547
rect 2409 501 2552 547
rect 2598 501 2757 547
rect 2803 501 2959 547
rect 3005 501 3163 547
rect 3209 501 3368 547
rect 3414 501 3573 547
rect 3619 501 3778 547
rect 3824 501 3981 547
rect 4027 501 4185 547
rect 4231 501 4242 547
rect 2293 490 4242 501
rect 1208 414 2210 430
rect 1208 368 1238 414
rect 1284 411 2210 414
rect 1284 368 1458 411
rect 1208 365 1458 368
rect 1504 365 1688 411
rect 1734 365 1912 411
rect 1958 365 2134 411
rect 2180 365 2210 411
rect 1208 354 2210 365
rect 2335 419 4207 430
rect 2381 373 2581 419
rect 2627 373 2806 419
rect 2852 373 3032 419
rect 3078 373 3255 419
rect 3301 373 3479 419
rect 3525 373 3702 419
rect 3748 373 3927 419
rect 3973 373 4150 419
rect 4196 373 4207 419
rect 2335 366 4207 373
rect 497 287 675 298
rect 543 217 675 287
rect 721 320 927 331
rect 767 274 927 320
rect 2335 298 2381 366
rect 4416 330 4537 673
rect 4416 320 4757 330
rect 721 263 927 274
rect 1127 287 2381 298
rect 1127 228 1575 287
rect 543 182 1127 217
rect 1173 182 1575 228
rect 543 173 1575 182
rect 543 171 1173 173
rect 273 128 319 139
rect 497 136 543 147
rect 1621 252 2023 287
rect 1575 136 1621 147
rect 2069 252 2381 287
rect 2471 319 4757 320
rect 2471 272 2919 319
rect 2517 226 2919 272
rect 2471 179 2919 226
rect 2965 179 3367 319
rect 3413 179 3815 319
rect 3861 179 4263 319
rect 4309 272 4757 319
rect 4309 226 4711 272
rect 4309 179 4757 226
rect 2471 173 4757 179
rect 4935 221 4981 232
rect 2023 136 2069 147
rect 0 82 273 90
rect 854 90 865 125
rect 319 82 865 90
rect 0 79 865 82
rect 911 90 922 125
rect 1340 90 1351 127
rect 911 81 1351 90
rect 1397 90 1408 127
rect 1788 90 1799 127
rect 1397 81 1799 90
rect 1845 90 1856 127
rect 2236 90 2247 127
rect 1845 81 2247 90
rect 2293 90 2304 127
rect 2684 90 2695 127
rect 2293 81 2695 90
rect 2741 90 2752 127
rect 3132 90 3143 127
rect 2741 81 3143 90
rect 3189 90 3200 127
rect 3580 90 3591 127
rect 3189 81 3591 90
rect 3637 90 3648 127
rect 4028 90 4039 127
rect 3637 81 4039 90
rect 4085 90 4096 127
rect 4476 90 4487 127
rect 4085 81 4487 90
rect 4533 90 4544 127
rect 4533 81 4935 90
rect 4981 81 5040 90
rect 911 79 5040 81
rect 0 -90 5040 79
<< labels >>
flabel metal1 s 142 466 315 542 0 FreeSans 200 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1208 354 2210 430 0 FreeSans 200 0 0 0 I
port 2 nsew default input
flabel metal1 s 0 918 5040 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 4935 139 4981 232 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 2451 673 4537 835 0 FreeSans 200 0 0 0 Z
port 3 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 4416 330 4537 673 1 Z
port 3 nsew default output
rlabel metal1 s 4416 320 4757 330 1 Z
port 3 nsew default output
rlabel metal1 s 2471 173 4757 320 1 Z
port 3 nsew default output
rlabel metal1 s 4695 881 4741 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4276 881 4344 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3868 881 3936 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3460 881 3528 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3052 881 3120 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2644 881 2712 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2247 881 2293 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1839 881 1885 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1431 881 1477 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1023 881 1069 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 881 347 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4695 776 4741 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2247 776 2293 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1839 776 1885 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1431 776 1477 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1023 776 1069 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 776 347 881 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 769 347 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4935 127 4981 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 127 319 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4935 125 4981 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4476 125 4544 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4028 125 4096 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3580 125 3648 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3132 125 3200 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2684 125 2752 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2236 125 2304 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1788 125 1856 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1340 125 1408 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 125 319 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4935 90 4981 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4476 90 4544 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4028 90 4096 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3580 90 3648 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3132 90 3200 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2684 90 2752 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2236 90 2304 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1788 90 1856 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1340 90 1408 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 854 90 922 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 5040 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5040 1008
string GDS_END 1367650
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1356782
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
