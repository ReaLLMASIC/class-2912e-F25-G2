magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 355 3558 870
rect -86 352 947 355
rect 2176 352 3558 355
<< pwell >>
rect 947 352 2176 355
rect -86 -86 3558 352
<< metal1 >>
rect 0 724 3472 844
rect 69 496 115 724
rect 464 430 546 674
rect 1260 558 1306 724
rect 54 354 314 430
rect 369 354 546 430
rect 262 60 330 212
rect 1213 60 1281 215
rect 1822 494 1868 724
rect 1821 60 1889 215
rect 2560 492 2606 724
rect 2805 336 2851 439
rect 2714 318 2851 336
rect 2362 290 2851 318
rect 3069 485 3137 724
rect 2362 242 2773 290
rect 2533 60 2601 152
rect 2981 60 3049 152
rect 3136 60 3182 219
rect 3260 126 3407 654
rect 0 -60 3472 60
<< obsm1 >>
rect 762 512 808 625
rect 1362 632 1758 678
rect 1362 512 1408 632
rect 600 466 1408 512
rect 38 258 423 304
rect 38 169 106 258
rect 377 215 423 258
rect 600 215 646 466
rect 1464 420 1510 580
rect 692 374 1510 420
rect 692 284 738 374
rect 377 169 554 215
rect 600 169 778 215
rect 1464 156 1510 374
rect 1608 315 1654 580
rect 1712 364 1758 632
rect 2036 632 2514 678
rect 1608 268 1982 315
rect 1608 156 1654 268
rect 2036 156 2102 632
rect 2356 499 2402 586
rect 2172 452 2402 499
rect 2172 152 2218 452
rect 2468 428 2514 632
rect 2468 382 2726 428
rect 2912 426 2958 636
rect 2912 358 3214 426
rect 2912 244 2958 358
rect 2868 198 2958 244
rect 2868 152 2914 198
rect 2172 106 2395 152
rect 2757 106 2914 152
<< labels >>
rlabel metal1 s 2362 242 2773 290 6 CLKN
port 1 nsew clock input
rlabel metal1 s 2362 290 2851 318 6 CLKN
port 1 nsew clock input
rlabel metal1 s 2714 318 2851 336 6 CLKN
port 1 nsew clock input
rlabel metal1 s 2805 336 2851 439 6 CLKN
port 1 nsew clock input
rlabel metal1 s 369 354 546 430 6 E
port 2 nsew default input
rlabel metal1 s 464 430 546 674 6 E
port 2 nsew default input
rlabel metal1 s 54 354 314 430 6 TE
port 3 nsew default input
rlabel metal1 s 3260 126 3407 654 6 Q
port 4 nsew default output
rlabel metal1 s 3069 485 3137 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2560 492 2606 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1822 494 1868 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1260 558 1306 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 496 115 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 724 3472 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel nwell s 2176 352 3558 355 6 VNW
port 6 nsew power bidirectional
rlabel nwell s -86 352 947 355 6 VNW
port 6 nsew power bidirectional
rlabel nwell s -86 355 3558 870 6 VNW
port 6 nsew power bidirectional
rlabel pwell s -86 -86 3558 352 6 VPW
port 7 nsew ground bidirectional
rlabel pwell s 947 352 2176 355 6 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 0 -60 3472 60 8 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3136 60 3182 219 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2981 60 3049 152 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2533 60 2601 152 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1821 60 1889 215 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1213 60 1281 215 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 212 6 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3472 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 433888
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 426350
<< end >>
