magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< deepnwell >>
rect -680 -680 788 2280
<< pbase >>
rect -180 -180 288 1780
<< ndiff >>
rect 0 1528 108 1600
rect 0 72 31 1528
rect 77 72 108 1528
rect 0 0 108 72
<< ndiffc >>
rect 31 72 77 1528
<< psubdiff >>
rect -1264 2845 1372 2864
rect -1264 2799 -1097 2845
rect 1205 2799 1372 2845
rect -1264 2780 1372 2799
rect -1264 2703 -1180 2780
rect -1264 -1103 -1245 2703
rect -1199 -1103 -1180 2703
rect 1288 2703 1372 2780
rect -148 1729 256 1748
rect -148 1683 -109 1729
rect 219 1683 256 1729
rect -148 1664 256 1683
rect -148 1622 -64 1664
rect -148 -22 -129 1622
rect -83 -22 -64 1622
rect 172 1622 256 1664
rect -148 -64 -64 -22
rect 172 -22 191 1622
rect 237 -22 256 1622
rect 172 -64 256 -22
rect -148 -148 256 -64
rect -1264 -1180 -1180 -1103
rect 1288 -1103 1307 2703
rect 1353 -1103 1372 2703
rect 1288 -1180 1372 -1103
rect -1264 -1199 1372 -1180
rect -1264 -1245 -1097 -1199
rect -769 -1245 877 -1199
rect 1205 -1245 1372 -1199
rect -1264 -1264 1372 -1245
<< nsubdiff >>
rect -296 1877 404 1896
rect -296 1831 -251 1877
rect 359 1831 404 1877
rect -296 1812 404 1831
rect -296 1763 -212 1812
rect -296 -163 -277 1763
rect -231 -163 -212 1763
rect 320 1763 404 1812
rect -296 -212 -212 -163
rect 320 -163 339 1763
rect 385 -163 404 1763
rect 320 -212 404 -163
rect -296 -296 404 -212
<< psubdiffcont >>
rect -1097 2799 1205 2845
rect -1245 -1103 -1199 2703
rect -109 1683 219 1729
rect -129 -22 -83 1622
rect 191 -22 237 1622
rect 1307 -1103 1353 2703
rect -1097 -1245 -769 -1199
rect 877 -1245 1205 -1199
<< nsubdiffcont >>
rect -251 1831 359 1877
rect -277 -163 -231 1763
rect 339 -163 385 1763
<< metal1 >>
rect -1264 2845 1372 2864
rect -1264 2799 -1097 2845
rect 1205 2799 1372 2845
rect -1264 2780 1372 2799
rect -1264 2703 -1180 2780
rect -1264 -1103 -1245 2703
rect -1199 -1103 -1180 2703
rect 1288 2703 1372 2780
rect -296 1877 404 1896
rect -296 1831 -251 1877
rect 359 1831 404 1877
rect -296 1812 404 1831
rect -296 1763 -212 1812
rect -296 -163 -277 1763
rect -231 -163 -212 1763
rect 320 1763 404 1812
rect -148 1729 256 1748
rect -148 1683 -109 1729
rect 219 1683 256 1729
rect -148 1664 256 1683
rect -148 1622 -64 1664
rect -148 -22 -129 1622
rect -83 -22 -64 1622
rect 172 1622 256 1664
rect 0 1528 108 1600
rect 0 72 31 1528
rect 77 72 108 1528
rect 0 0 108 72
rect -148 -148 -64 -22
rect 172 -22 191 1622
rect 237 -22 256 1622
rect 172 -148 256 -22
rect -296 -296 -212 -163
rect 320 -163 339 1763
rect 385 -163 404 1763
rect 320 -296 404 -163
rect -1264 -1180 -1180 -1103
rect 1288 -1103 1307 2703
rect 1353 -1103 1372 2703
rect 1288 -1180 1372 -1103
rect -1264 -1199 -680 -1180
rect -1264 -1245 -1097 -1199
rect -769 -1245 -680 -1199
rect -1264 -1264 -680 -1245
rect 788 -1199 1372 -1180
rect 788 -1245 877 -1199
rect 1205 -1245 1372 -1199
rect 788 -1264 1372 -1245
<< labels >>
flabel ndiffc 54 900 54 900 0 FreeSans 400 0 0 0 E
flabel metal1 -108 -106 -108 -106 0 FreeSans 400 0 0 0 B
flabel metal1 208 -100 208 -100 0 FreeSans 400 0 0 0 B
flabel psubdiffcont 213 1703 213 1703 0 FreeSans 400 0 0 0 B
flabel metal1 362 -255 362 -255 0 FreeSans 400 0 0 0 C
flabel metal1 365 1857 365 1857 0 FreeSans 400 0 0 0 C
flabel metal1 -252 -251 -252 -251 0 FreeSans 400 0 0 0 C
flabel metal1 1332 -1219 1332 -1219 0 FreeSans 400 0 0 0 S
flabel metal1 1332 -1219 1332 -1219 0 FreeSans 400 0 0 0 S
flabel metal1 1333 2824 1333 2824 0 FreeSans 400 0 0 0 S
flabel metal1 -1220 -1222 -1220 -1222 0 FreeSans 400 0 0 0 S
flabel metal1 -1220 -1222 -1220 -1222 0 FreeSans 400 0 0 0 S
<< properties >>
string GDS_END 17388
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/npn_00p54x08p00.gds
string GDS_START 112
string gencell npn_00p54x08p00
<< end >>
