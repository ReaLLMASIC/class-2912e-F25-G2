magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -27 702 7407 2956
<< mvnmos >>
rect 252 3214 372 3614
rect 476 3214 596 3614
rect 700 3214 820 3614
rect 2023 3214 2143 3598
rect 2247 3214 2367 3598
rect 2471 3214 2591 3598
rect 2695 3214 2815 3598
rect 2919 3214 3039 3598
rect 3143 3214 3263 3598
rect 3367 3214 3487 3598
rect 3591 3214 3711 3598
rect 3815 3214 3935 3598
rect 4039 3214 4159 3598
rect 4669 3214 4789 3598
rect 4893 3214 5013 3598
rect 5117 3214 5237 3598
rect 5341 3214 5461 3598
rect 5565 3214 5685 3598
rect 5789 3214 5909 3598
rect 6013 3214 6133 3598
rect 6237 3214 6357 3598
rect 6461 3214 6581 3598
rect 6685 3214 6805 3598
rect 509 213 629 405
rect 733 213 853 405
rect 1181 295 1301 487
rect 1688 109 1808 563
rect 2150 372 2270 564
rect 2374 372 2494 564
rect 2822 372 2942 564
rect 3293 324 3413 564
rect 3517 324 3637 564
rect 3950 109 4070 563
rect 4174 109 4294 563
rect 4618 248 4738 440
rect 4842 248 4962 440
rect 5307 381 5427 559
rect 5531 381 5651 559
rect 5755 381 5875 559
rect 5979 381 6099 559
rect 6203 381 6323 559
rect 6427 381 6547 559
rect 6651 381 6771 559
<< mvpmos >>
rect 252 1884 372 2380
rect 476 1884 596 2380
rect 700 1884 820 2380
rect 924 1884 1044 2380
rect 1148 1884 1268 2380
rect 1372 1884 1492 2380
rect 2023 1884 2143 2828
rect 2247 1884 2367 2828
rect 2471 1884 2591 2828
rect 2695 1884 2815 2828
rect 2919 1884 3039 2828
rect 3143 1884 3263 2828
rect 3367 1884 3487 2828
rect 3591 1884 3711 2828
rect 3815 1884 3935 2828
rect 4039 1884 4159 2828
rect 4669 1884 4789 2828
rect 4893 1884 5013 2828
rect 5117 1884 5237 2828
rect 5341 1884 5461 2828
rect 5565 1884 5685 2828
rect 5789 1884 5909 2828
rect 6013 1884 6133 2828
rect 6237 1884 6357 2828
rect 6461 1884 6581 2828
rect 6685 1884 6805 2828
rect 509 843 629 1297
rect 733 843 853 1297
rect 1181 843 1301 1297
rect 1688 843 1808 1297
rect 2036 843 2156 1035
rect 2374 843 2494 1297
rect 2822 843 2942 1297
rect 3293 843 3413 1411
rect 3517 843 3637 1411
rect 3950 843 4070 1297
rect 4174 843 4294 1297
rect 4510 1105 4630 1297
rect 4842 843 4962 1297
rect 5307 843 5427 1283
rect 5531 843 5651 1283
rect 5755 843 5875 1283
rect 5979 843 6099 1283
rect 6203 843 6323 1283
rect 6427 843 6547 1283
rect 6651 843 6771 1283
<< ndiff >>
rect 79 484 233 541
rect 79 438 133 484
rect 179 438 233 484
rect 79 320 233 438
rect 79 274 133 320
rect 179 274 233 320
rect 79 218 233 274
<< mvndiff >>
rect 164 3601 252 3614
rect 164 3555 177 3601
rect 223 3555 252 3601
rect 164 3492 252 3555
rect 164 3446 177 3492
rect 223 3446 252 3492
rect 164 3383 252 3446
rect 164 3337 177 3383
rect 223 3337 252 3383
rect 164 3273 252 3337
rect 164 3227 177 3273
rect 223 3227 252 3273
rect 164 3214 252 3227
rect 372 3601 476 3614
rect 372 3555 401 3601
rect 447 3555 476 3601
rect 372 3492 476 3555
rect 372 3446 401 3492
rect 447 3446 476 3492
rect 372 3383 476 3446
rect 372 3337 401 3383
rect 447 3337 476 3383
rect 372 3273 476 3337
rect 372 3227 401 3273
rect 447 3227 476 3273
rect 372 3214 476 3227
rect 596 3601 700 3614
rect 596 3555 625 3601
rect 671 3555 700 3601
rect 596 3492 700 3555
rect 596 3446 625 3492
rect 671 3446 700 3492
rect 596 3383 700 3446
rect 596 3337 625 3383
rect 671 3337 700 3383
rect 596 3273 700 3337
rect 596 3227 625 3273
rect 671 3227 700 3273
rect 596 3214 700 3227
rect 820 3601 908 3614
rect 820 3555 849 3601
rect 895 3555 908 3601
rect 820 3492 908 3555
rect 1935 3585 2023 3598
rect 820 3446 849 3492
rect 895 3446 908 3492
rect 820 3383 908 3446
rect 820 3337 849 3383
rect 895 3337 908 3383
rect 820 3273 908 3337
rect 820 3227 849 3273
rect 895 3227 908 3273
rect 1935 3539 1948 3585
rect 1994 3539 2023 3585
rect 1935 3481 2023 3539
rect 1935 3435 1948 3481
rect 1994 3435 2023 3481
rect 1935 3377 2023 3435
rect 1935 3331 1948 3377
rect 1994 3331 2023 3377
rect 1935 3273 2023 3331
rect 820 3214 908 3227
rect 1935 3227 1948 3273
rect 1994 3227 2023 3273
rect 1935 3214 2023 3227
rect 2143 3585 2247 3598
rect 2143 3539 2172 3585
rect 2218 3539 2247 3585
rect 2143 3481 2247 3539
rect 2143 3435 2172 3481
rect 2218 3435 2247 3481
rect 2143 3377 2247 3435
rect 2143 3331 2172 3377
rect 2218 3331 2247 3377
rect 2143 3273 2247 3331
rect 2143 3227 2172 3273
rect 2218 3227 2247 3273
rect 2143 3214 2247 3227
rect 2367 3585 2471 3598
rect 2367 3539 2396 3585
rect 2442 3539 2471 3585
rect 2367 3481 2471 3539
rect 2367 3435 2396 3481
rect 2442 3435 2471 3481
rect 2367 3377 2471 3435
rect 2367 3331 2396 3377
rect 2442 3331 2471 3377
rect 2367 3273 2471 3331
rect 2367 3227 2396 3273
rect 2442 3227 2471 3273
rect 2367 3214 2471 3227
rect 2591 3585 2695 3598
rect 2591 3539 2620 3585
rect 2666 3539 2695 3585
rect 2591 3481 2695 3539
rect 2591 3435 2620 3481
rect 2666 3435 2695 3481
rect 2591 3377 2695 3435
rect 2591 3331 2620 3377
rect 2666 3331 2695 3377
rect 2591 3273 2695 3331
rect 2591 3227 2620 3273
rect 2666 3227 2695 3273
rect 2591 3214 2695 3227
rect 2815 3585 2919 3598
rect 2815 3539 2844 3585
rect 2890 3539 2919 3585
rect 2815 3481 2919 3539
rect 2815 3435 2844 3481
rect 2890 3435 2919 3481
rect 2815 3377 2919 3435
rect 2815 3331 2844 3377
rect 2890 3331 2919 3377
rect 2815 3273 2919 3331
rect 2815 3227 2844 3273
rect 2890 3227 2919 3273
rect 2815 3214 2919 3227
rect 3039 3585 3143 3598
rect 3039 3539 3068 3585
rect 3114 3539 3143 3585
rect 3039 3481 3143 3539
rect 3039 3435 3068 3481
rect 3114 3435 3143 3481
rect 3039 3377 3143 3435
rect 3039 3331 3068 3377
rect 3114 3331 3143 3377
rect 3039 3273 3143 3331
rect 3039 3227 3068 3273
rect 3114 3227 3143 3273
rect 3039 3214 3143 3227
rect 3263 3585 3367 3598
rect 3263 3539 3292 3585
rect 3338 3539 3367 3585
rect 3263 3481 3367 3539
rect 3263 3435 3292 3481
rect 3338 3435 3367 3481
rect 3263 3377 3367 3435
rect 3263 3331 3292 3377
rect 3338 3331 3367 3377
rect 3263 3273 3367 3331
rect 3263 3227 3292 3273
rect 3338 3227 3367 3273
rect 3263 3214 3367 3227
rect 3487 3585 3591 3598
rect 3487 3539 3516 3585
rect 3562 3539 3591 3585
rect 3487 3481 3591 3539
rect 3487 3435 3516 3481
rect 3562 3435 3591 3481
rect 3487 3377 3591 3435
rect 3487 3331 3516 3377
rect 3562 3331 3591 3377
rect 3487 3273 3591 3331
rect 3487 3227 3516 3273
rect 3562 3227 3591 3273
rect 3487 3214 3591 3227
rect 3711 3585 3815 3598
rect 3711 3539 3740 3585
rect 3786 3539 3815 3585
rect 3711 3481 3815 3539
rect 3711 3435 3740 3481
rect 3786 3435 3815 3481
rect 3711 3377 3815 3435
rect 3711 3331 3740 3377
rect 3786 3331 3815 3377
rect 3711 3273 3815 3331
rect 3711 3227 3740 3273
rect 3786 3227 3815 3273
rect 3711 3214 3815 3227
rect 3935 3585 4039 3598
rect 3935 3539 3964 3585
rect 4010 3539 4039 3585
rect 3935 3481 4039 3539
rect 3935 3435 3964 3481
rect 4010 3435 4039 3481
rect 3935 3377 4039 3435
rect 3935 3331 3964 3377
rect 4010 3331 4039 3377
rect 3935 3273 4039 3331
rect 3935 3227 3964 3273
rect 4010 3227 4039 3273
rect 3935 3214 4039 3227
rect 4159 3585 4247 3598
rect 4159 3539 4188 3585
rect 4234 3539 4247 3585
rect 4581 3585 4669 3598
rect 4159 3481 4247 3539
rect 4159 3435 4188 3481
rect 4234 3435 4247 3481
rect 4159 3377 4247 3435
rect 4159 3331 4188 3377
rect 4234 3331 4247 3377
rect 4159 3273 4247 3331
rect 4159 3227 4188 3273
rect 4234 3227 4247 3273
rect 4581 3539 4594 3585
rect 4640 3539 4669 3585
rect 4581 3481 4669 3539
rect 4581 3435 4594 3481
rect 4640 3435 4669 3481
rect 4581 3377 4669 3435
rect 4581 3331 4594 3377
rect 4640 3331 4669 3377
rect 4581 3273 4669 3331
rect 4159 3214 4247 3227
rect 4581 3227 4594 3273
rect 4640 3227 4669 3273
rect 4581 3214 4669 3227
rect 4789 3585 4893 3598
rect 4789 3539 4818 3585
rect 4864 3539 4893 3585
rect 4789 3481 4893 3539
rect 4789 3435 4818 3481
rect 4864 3435 4893 3481
rect 4789 3377 4893 3435
rect 4789 3331 4818 3377
rect 4864 3331 4893 3377
rect 4789 3273 4893 3331
rect 4789 3227 4818 3273
rect 4864 3227 4893 3273
rect 4789 3214 4893 3227
rect 5013 3585 5117 3598
rect 5013 3539 5042 3585
rect 5088 3539 5117 3585
rect 5013 3481 5117 3539
rect 5013 3435 5042 3481
rect 5088 3435 5117 3481
rect 5013 3377 5117 3435
rect 5013 3331 5042 3377
rect 5088 3331 5117 3377
rect 5013 3273 5117 3331
rect 5013 3227 5042 3273
rect 5088 3227 5117 3273
rect 5013 3214 5117 3227
rect 5237 3585 5341 3598
rect 5237 3539 5266 3585
rect 5312 3539 5341 3585
rect 5237 3481 5341 3539
rect 5237 3435 5266 3481
rect 5312 3435 5341 3481
rect 5237 3377 5341 3435
rect 5237 3331 5266 3377
rect 5312 3331 5341 3377
rect 5237 3273 5341 3331
rect 5237 3227 5266 3273
rect 5312 3227 5341 3273
rect 5237 3214 5341 3227
rect 5461 3585 5565 3598
rect 5461 3539 5490 3585
rect 5536 3539 5565 3585
rect 5461 3481 5565 3539
rect 5461 3435 5490 3481
rect 5536 3435 5565 3481
rect 5461 3377 5565 3435
rect 5461 3331 5490 3377
rect 5536 3331 5565 3377
rect 5461 3273 5565 3331
rect 5461 3227 5490 3273
rect 5536 3227 5565 3273
rect 5461 3214 5565 3227
rect 5685 3585 5789 3598
rect 5685 3539 5714 3585
rect 5760 3539 5789 3585
rect 5685 3481 5789 3539
rect 5685 3435 5714 3481
rect 5760 3435 5789 3481
rect 5685 3377 5789 3435
rect 5685 3331 5714 3377
rect 5760 3331 5789 3377
rect 5685 3273 5789 3331
rect 5685 3227 5714 3273
rect 5760 3227 5789 3273
rect 5685 3214 5789 3227
rect 5909 3585 6013 3598
rect 5909 3539 5938 3585
rect 5984 3539 6013 3585
rect 5909 3481 6013 3539
rect 5909 3435 5938 3481
rect 5984 3435 6013 3481
rect 5909 3377 6013 3435
rect 5909 3331 5938 3377
rect 5984 3331 6013 3377
rect 5909 3273 6013 3331
rect 5909 3227 5938 3273
rect 5984 3227 6013 3273
rect 5909 3214 6013 3227
rect 6133 3585 6237 3598
rect 6133 3539 6162 3585
rect 6208 3539 6237 3585
rect 6133 3481 6237 3539
rect 6133 3435 6162 3481
rect 6208 3435 6237 3481
rect 6133 3377 6237 3435
rect 6133 3331 6162 3377
rect 6208 3331 6237 3377
rect 6133 3273 6237 3331
rect 6133 3227 6162 3273
rect 6208 3227 6237 3273
rect 6133 3214 6237 3227
rect 6357 3585 6461 3598
rect 6357 3539 6386 3585
rect 6432 3539 6461 3585
rect 6357 3481 6461 3539
rect 6357 3435 6386 3481
rect 6432 3435 6461 3481
rect 6357 3377 6461 3435
rect 6357 3331 6386 3377
rect 6432 3331 6461 3377
rect 6357 3273 6461 3331
rect 6357 3227 6386 3273
rect 6432 3227 6461 3273
rect 6357 3214 6461 3227
rect 6581 3585 6685 3598
rect 6581 3539 6610 3585
rect 6656 3539 6685 3585
rect 6581 3481 6685 3539
rect 6581 3435 6610 3481
rect 6656 3435 6685 3481
rect 6581 3377 6685 3435
rect 6581 3331 6610 3377
rect 6656 3331 6685 3377
rect 6581 3273 6685 3331
rect 6581 3227 6610 3273
rect 6656 3227 6685 3273
rect 6581 3214 6685 3227
rect 6805 3585 6893 3598
rect 6805 3539 6834 3585
rect 6880 3539 6893 3585
rect 6805 3481 6893 3539
rect 6805 3435 6834 3481
rect 6880 3435 6893 3481
rect 6805 3377 6893 3435
rect 6805 3331 6834 3377
rect 6880 3331 6893 3377
rect 6805 3273 6893 3331
rect 6805 3227 6834 3273
rect 6880 3227 6893 3273
rect 6805 3214 6893 3227
rect 1600 550 1688 563
rect 1600 504 1613 550
rect 1659 504 1688 550
rect 1093 474 1181 487
rect 1093 428 1106 474
rect 1152 428 1181 474
rect 421 392 509 405
rect 421 346 434 392
rect 480 346 509 392
rect 421 272 509 346
rect 421 226 434 272
rect 480 226 509 272
rect 421 213 509 226
rect 629 392 733 405
rect 629 346 658 392
rect 704 346 733 392
rect 629 272 733 346
rect 629 226 658 272
rect 704 226 733 272
rect 629 213 733 226
rect 853 392 941 405
rect 853 346 882 392
rect 928 346 941 392
rect 853 272 941 346
rect 1093 354 1181 428
rect 1093 308 1106 354
rect 1152 308 1181 354
rect 1093 295 1181 308
rect 1301 474 1389 487
rect 1301 428 1330 474
rect 1376 428 1389 474
rect 1301 354 1389 428
rect 1301 308 1330 354
rect 1376 308 1389 354
rect 1301 295 1389 308
rect 1600 423 1688 504
rect 1600 377 1613 423
rect 1659 377 1688 423
rect 1600 296 1688 377
rect 853 226 882 272
rect 928 226 941 272
rect 853 213 941 226
rect 1600 250 1613 296
rect 1659 250 1688 296
rect 1600 168 1688 250
rect 1600 122 1613 168
rect 1659 122 1688 168
rect 1600 109 1688 122
rect 1808 550 1896 563
rect 1808 504 1837 550
rect 1883 504 1896 550
rect 1808 423 1896 504
rect 1808 377 1837 423
rect 1883 377 1896 423
rect 1808 296 1896 377
rect 2062 551 2150 564
rect 2062 505 2075 551
rect 2121 505 2150 551
rect 2062 431 2150 505
rect 2062 385 2075 431
rect 2121 385 2150 431
rect 2062 372 2150 385
rect 2270 551 2374 564
rect 2270 505 2299 551
rect 2345 505 2374 551
rect 2270 431 2374 505
rect 2270 385 2299 431
rect 2345 385 2374 431
rect 2270 372 2374 385
rect 2494 551 2582 564
rect 2494 505 2523 551
rect 2569 505 2582 551
rect 2494 431 2582 505
rect 2494 385 2523 431
rect 2569 385 2582 431
rect 2494 372 2582 385
rect 2734 551 2822 564
rect 2734 505 2747 551
rect 2793 505 2822 551
rect 2734 431 2822 505
rect 2734 385 2747 431
rect 2793 385 2822 431
rect 2734 372 2822 385
rect 2942 551 3030 564
rect 2942 505 2971 551
rect 3017 505 3030 551
rect 2942 431 3030 505
rect 2942 385 2971 431
rect 3017 385 3030 431
rect 2942 372 3030 385
rect 3205 551 3293 564
rect 3205 505 3218 551
rect 3264 505 3293 551
rect 3205 383 3293 505
rect 1808 250 1837 296
rect 1883 250 1896 296
rect 1808 168 1896 250
rect 1808 122 1837 168
rect 1883 122 1896 168
rect 1808 109 1896 122
rect 3205 337 3218 383
rect 3264 337 3293 383
rect 3205 324 3293 337
rect 3413 551 3517 564
rect 3413 505 3442 551
rect 3488 505 3517 551
rect 3413 383 3517 505
rect 3413 337 3442 383
rect 3488 337 3517 383
rect 3413 324 3517 337
rect 3637 551 3725 564
rect 3637 505 3666 551
rect 3712 505 3725 551
rect 3637 383 3725 505
rect 3637 337 3666 383
rect 3712 337 3725 383
rect 3637 324 3725 337
rect 3862 550 3950 563
rect 3862 504 3875 550
rect 3921 504 3950 550
rect 3862 423 3950 504
rect 3862 377 3875 423
rect 3921 377 3950 423
rect 3862 296 3950 377
rect 3862 250 3875 296
rect 3921 250 3950 296
rect 3862 168 3950 250
rect 3862 122 3875 168
rect 3921 122 3950 168
rect 3862 109 3950 122
rect 4070 550 4174 563
rect 4070 504 4099 550
rect 4145 504 4174 550
rect 4070 423 4174 504
rect 4070 377 4099 423
rect 4145 377 4174 423
rect 4070 296 4174 377
rect 4070 250 4099 296
rect 4145 250 4174 296
rect 4070 168 4174 250
rect 4070 122 4099 168
rect 4145 122 4174 168
rect 4070 109 4174 122
rect 4294 550 4382 563
rect 4294 504 4323 550
rect 4369 504 4382 550
rect 4294 423 4382 504
rect 5219 546 5307 559
rect 5219 500 5232 546
rect 5278 500 5307 546
rect 5219 440 5307 500
rect 4294 377 4323 423
rect 4369 377 4382 423
rect 4294 296 4382 377
rect 4294 250 4323 296
rect 4369 250 4382 296
rect 4294 168 4382 250
rect 4530 427 4618 440
rect 4530 381 4543 427
rect 4589 381 4618 427
rect 4530 307 4618 381
rect 4530 261 4543 307
rect 4589 261 4618 307
rect 4530 248 4618 261
rect 4738 427 4842 440
rect 4738 381 4767 427
rect 4813 381 4842 427
rect 4738 307 4842 381
rect 4738 261 4767 307
rect 4813 261 4842 307
rect 4738 248 4842 261
rect 4962 427 5050 440
rect 4962 381 4991 427
rect 5037 381 5050 427
rect 5219 394 5232 440
rect 5278 394 5307 440
rect 5219 381 5307 394
rect 5427 546 5531 559
rect 5427 500 5456 546
rect 5502 500 5531 546
rect 5427 440 5531 500
rect 5427 394 5456 440
rect 5502 394 5531 440
rect 5427 381 5531 394
rect 5651 546 5755 559
rect 5651 500 5680 546
rect 5726 500 5755 546
rect 5651 440 5755 500
rect 5651 394 5680 440
rect 5726 394 5755 440
rect 5651 381 5755 394
rect 5875 546 5979 559
rect 5875 500 5904 546
rect 5950 500 5979 546
rect 5875 440 5979 500
rect 5875 394 5904 440
rect 5950 394 5979 440
rect 5875 381 5979 394
rect 6099 546 6203 559
rect 6099 500 6128 546
rect 6174 500 6203 546
rect 6099 440 6203 500
rect 6099 394 6128 440
rect 6174 394 6203 440
rect 6099 381 6203 394
rect 6323 546 6427 559
rect 6323 500 6352 546
rect 6398 500 6427 546
rect 6323 440 6427 500
rect 6323 394 6352 440
rect 6398 394 6427 440
rect 6323 381 6427 394
rect 6547 546 6651 559
rect 6547 500 6576 546
rect 6622 500 6651 546
rect 6547 440 6651 500
rect 6547 394 6576 440
rect 6622 394 6651 440
rect 6547 381 6651 394
rect 6771 546 6859 559
rect 6771 500 6800 546
rect 6846 500 6859 546
rect 6771 440 6859 500
rect 6771 394 6800 440
rect 6846 394 6859 440
rect 6771 381 6859 394
rect 4962 307 5050 381
rect 4962 261 4991 307
rect 5037 261 5050 307
rect 4962 248 5050 261
rect 4294 122 4323 168
rect 4369 122 4382 168
rect 4294 109 4382 122
<< mvpdiff >>
rect 1935 2815 2023 2828
rect 1935 2769 1948 2815
rect 1994 2769 2023 2815
rect 1935 2706 2023 2769
rect 1935 2660 1948 2706
rect 1994 2660 2023 2706
rect 1935 2597 2023 2660
rect 1935 2551 1948 2597
rect 1994 2551 2023 2597
rect 1935 2488 2023 2551
rect 1935 2442 1948 2488
rect 1994 2442 2023 2488
rect 164 2367 252 2380
rect 164 2321 177 2367
rect 223 2321 252 2367
rect 164 2261 252 2321
rect 164 2215 177 2261
rect 223 2215 252 2261
rect 164 2155 252 2215
rect 164 2109 177 2155
rect 223 2109 252 2155
rect 164 2049 252 2109
rect 164 2003 177 2049
rect 223 2003 252 2049
rect 164 1943 252 2003
rect 164 1897 177 1943
rect 223 1897 252 1943
rect 164 1884 252 1897
rect 372 2367 476 2380
rect 372 2321 401 2367
rect 447 2321 476 2367
rect 372 2261 476 2321
rect 372 2215 401 2261
rect 447 2215 476 2261
rect 372 2155 476 2215
rect 372 2109 401 2155
rect 447 2109 476 2155
rect 372 2049 476 2109
rect 372 2003 401 2049
rect 447 2003 476 2049
rect 372 1943 476 2003
rect 372 1897 401 1943
rect 447 1897 476 1943
rect 372 1884 476 1897
rect 596 2367 700 2380
rect 596 2321 625 2367
rect 671 2321 700 2367
rect 596 2261 700 2321
rect 596 2215 625 2261
rect 671 2215 700 2261
rect 596 2155 700 2215
rect 596 2109 625 2155
rect 671 2109 700 2155
rect 596 2049 700 2109
rect 596 2003 625 2049
rect 671 2003 700 2049
rect 596 1943 700 2003
rect 596 1897 625 1943
rect 671 1897 700 1943
rect 596 1884 700 1897
rect 820 2367 924 2380
rect 820 2321 849 2367
rect 895 2321 924 2367
rect 820 2261 924 2321
rect 820 2215 849 2261
rect 895 2215 924 2261
rect 820 2155 924 2215
rect 820 2109 849 2155
rect 895 2109 924 2155
rect 820 2049 924 2109
rect 820 2003 849 2049
rect 895 2003 924 2049
rect 820 1943 924 2003
rect 820 1897 849 1943
rect 895 1897 924 1943
rect 820 1884 924 1897
rect 1044 2367 1148 2380
rect 1044 2321 1073 2367
rect 1119 2321 1148 2367
rect 1044 2261 1148 2321
rect 1044 2215 1073 2261
rect 1119 2215 1148 2261
rect 1044 2155 1148 2215
rect 1044 2109 1073 2155
rect 1119 2109 1148 2155
rect 1044 2049 1148 2109
rect 1044 2003 1073 2049
rect 1119 2003 1148 2049
rect 1044 1943 1148 2003
rect 1044 1897 1073 1943
rect 1119 1897 1148 1943
rect 1044 1884 1148 1897
rect 1268 2367 1372 2380
rect 1268 2321 1297 2367
rect 1343 2321 1372 2367
rect 1268 2261 1372 2321
rect 1268 2215 1297 2261
rect 1343 2215 1372 2261
rect 1268 2155 1372 2215
rect 1268 2109 1297 2155
rect 1343 2109 1372 2155
rect 1268 2049 1372 2109
rect 1268 2003 1297 2049
rect 1343 2003 1372 2049
rect 1268 1943 1372 2003
rect 1268 1897 1297 1943
rect 1343 1897 1372 1943
rect 1268 1884 1372 1897
rect 1492 2367 1580 2380
rect 1492 2321 1521 2367
rect 1567 2321 1580 2367
rect 1492 2261 1580 2321
rect 1935 2379 2023 2442
rect 1935 2333 1948 2379
rect 1994 2333 2023 2379
rect 1935 2270 2023 2333
rect 1492 2215 1521 2261
rect 1567 2215 1580 2261
rect 1492 2155 1580 2215
rect 1492 2109 1521 2155
rect 1567 2109 1580 2155
rect 1492 2049 1580 2109
rect 1492 2003 1521 2049
rect 1567 2003 1580 2049
rect 1492 1943 1580 2003
rect 1935 2224 1948 2270
rect 1994 2224 2023 2270
rect 1935 2161 2023 2224
rect 1935 2115 1948 2161
rect 1994 2115 2023 2161
rect 1935 2052 2023 2115
rect 1935 2006 1948 2052
rect 1994 2006 2023 2052
rect 1492 1897 1521 1943
rect 1567 1897 1580 1943
rect 1492 1884 1580 1897
rect 1935 1943 2023 2006
rect 1935 1897 1948 1943
rect 1994 1897 2023 1943
rect 1935 1884 2023 1897
rect 2143 2815 2247 2828
rect 2143 2769 2172 2815
rect 2218 2769 2247 2815
rect 2143 2706 2247 2769
rect 2143 2660 2172 2706
rect 2218 2660 2247 2706
rect 2143 2597 2247 2660
rect 2143 2551 2172 2597
rect 2218 2551 2247 2597
rect 2143 2488 2247 2551
rect 2143 2442 2172 2488
rect 2218 2442 2247 2488
rect 2143 2379 2247 2442
rect 2143 2333 2172 2379
rect 2218 2333 2247 2379
rect 2143 2270 2247 2333
rect 2143 2224 2172 2270
rect 2218 2224 2247 2270
rect 2143 2161 2247 2224
rect 2143 2115 2172 2161
rect 2218 2115 2247 2161
rect 2143 2052 2247 2115
rect 2143 2006 2172 2052
rect 2218 2006 2247 2052
rect 2143 1943 2247 2006
rect 2143 1897 2172 1943
rect 2218 1897 2247 1943
rect 2143 1884 2247 1897
rect 2367 2815 2471 2828
rect 2367 2769 2396 2815
rect 2442 2769 2471 2815
rect 2367 2706 2471 2769
rect 2367 2660 2396 2706
rect 2442 2660 2471 2706
rect 2367 2597 2471 2660
rect 2367 2551 2396 2597
rect 2442 2551 2471 2597
rect 2367 2488 2471 2551
rect 2367 2442 2396 2488
rect 2442 2442 2471 2488
rect 2367 2379 2471 2442
rect 2367 2333 2396 2379
rect 2442 2333 2471 2379
rect 2367 2270 2471 2333
rect 2367 2224 2396 2270
rect 2442 2224 2471 2270
rect 2367 2161 2471 2224
rect 2367 2115 2396 2161
rect 2442 2115 2471 2161
rect 2367 2052 2471 2115
rect 2367 2006 2396 2052
rect 2442 2006 2471 2052
rect 2367 1943 2471 2006
rect 2367 1897 2396 1943
rect 2442 1897 2471 1943
rect 2367 1884 2471 1897
rect 2591 2815 2695 2828
rect 2591 2769 2620 2815
rect 2666 2769 2695 2815
rect 2591 2706 2695 2769
rect 2591 2660 2620 2706
rect 2666 2660 2695 2706
rect 2591 2597 2695 2660
rect 2591 2551 2620 2597
rect 2666 2551 2695 2597
rect 2591 2488 2695 2551
rect 2591 2442 2620 2488
rect 2666 2442 2695 2488
rect 2591 2379 2695 2442
rect 2591 2333 2620 2379
rect 2666 2333 2695 2379
rect 2591 2270 2695 2333
rect 2591 2224 2620 2270
rect 2666 2224 2695 2270
rect 2591 2161 2695 2224
rect 2591 2115 2620 2161
rect 2666 2115 2695 2161
rect 2591 2052 2695 2115
rect 2591 2006 2620 2052
rect 2666 2006 2695 2052
rect 2591 1943 2695 2006
rect 2591 1897 2620 1943
rect 2666 1897 2695 1943
rect 2591 1884 2695 1897
rect 2815 2815 2919 2828
rect 2815 2769 2844 2815
rect 2890 2769 2919 2815
rect 2815 2706 2919 2769
rect 2815 2660 2844 2706
rect 2890 2660 2919 2706
rect 2815 2597 2919 2660
rect 2815 2551 2844 2597
rect 2890 2551 2919 2597
rect 2815 2488 2919 2551
rect 2815 2442 2844 2488
rect 2890 2442 2919 2488
rect 2815 2379 2919 2442
rect 2815 2333 2844 2379
rect 2890 2333 2919 2379
rect 2815 2270 2919 2333
rect 2815 2224 2844 2270
rect 2890 2224 2919 2270
rect 2815 2161 2919 2224
rect 2815 2115 2844 2161
rect 2890 2115 2919 2161
rect 2815 2052 2919 2115
rect 2815 2006 2844 2052
rect 2890 2006 2919 2052
rect 2815 1943 2919 2006
rect 2815 1897 2844 1943
rect 2890 1897 2919 1943
rect 2815 1884 2919 1897
rect 3039 2815 3143 2828
rect 3039 2769 3068 2815
rect 3114 2769 3143 2815
rect 3039 2706 3143 2769
rect 3039 2660 3068 2706
rect 3114 2660 3143 2706
rect 3039 2597 3143 2660
rect 3039 2551 3068 2597
rect 3114 2551 3143 2597
rect 3039 2488 3143 2551
rect 3039 2442 3068 2488
rect 3114 2442 3143 2488
rect 3039 2379 3143 2442
rect 3039 2333 3068 2379
rect 3114 2333 3143 2379
rect 3039 2270 3143 2333
rect 3039 2224 3068 2270
rect 3114 2224 3143 2270
rect 3039 2161 3143 2224
rect 3039 2115 3068 2161
rect 3114 2115 3143 2161
rect 3039 2052 3143 2115
rect 3039 2006 3068 2052
rect 3114 2006 3143 2052
rect 3039 1943 3143 2006
rect 3039 1897 3068 1943
rect 3114 1897 3143 1943
rect 3039 1884 3143 1897
rect 3263 2815 3367 2828
rect 3263 2769 3292 2815
rect 3338 2769 3367 2815
rect 3263 2706 3367 2769
rect 3263 2660 3292 2706
rect 3338 2660 3367 2706
rect 3263 2597 3367 2660
rect 3263 2551 3292 2597
rect 3338 2551 3367 2597
rect 3263 2488 3367 2551
rect 3263 2442 3292 2488
rect 3338 2442 3367 2488
rect 3263 2379 3367 2442
rect 3263 2333 3292 2379
rect 3338 2333 3367 2379
rect 3263 2270 3367 2333
rect 3263 2224 3292 2270
rect 3338 2224 3367 2270
rect 3263 2161 3367 2224
rect 3263 2115 3292 2161
rect 3338 2115 3367 2161
rect 3263 2052 3367 2115
rect 3263 2006 3292 2052
rect 3338 2006 3367 2052
rect 3263 1943 3367 2006
rect 3263 1897 3292 1943
rect 3338 1897 3367 1943
rect 3263 1884 3367 1897
rect 3487 2815 3591 2828
rect 3487 2769 3516 2815
rect 3562 2769 3591 2815
rect 3487 2706 3591 2769
rect 3487 2660 3516 2706
rect 3562 2660 3591 2706
rect 3487 2597 3591 2660
rect 3487 2551 3516 2597
rect 3562 2551 3591 2597
rect 3487 2488 3591 2551
rect 3487 2442 3516 2488
rect 3562 2442 3591 2488
rect 3487 2379 3591 2442
rect 3487 2333 3516 2379
rect 3562 2333 3591 2379
rect 3487 2270 3591 2333
rect 3487 2224 3516 2270
rect 3562 2224 3591 2270
rect 3487 2161 3591 2224
rect 3487 2115 3516 2161
rect 3562 2115 3591 2161
rect 3487 2052 3591 2115
rect 3487 2006 3516 2052
rect 3562 2006 3591 2052
rect 3487 1943 3591 2006
rect 3487 1897 3516 1943
rect 3562 1897 3591 1943
rect 3487 1884 3591 1897
rect 3711 2815 3815 2828
rect 3711 2769 3740 2815
rect 3786 2769 3815 2815
rect 3711 2706 3815 2769
rect 3711 2660 3740 2706
rect 3786 2660 3815 2706
rect 3711 2597 3815 2660
rect 3711 2551 3740 2597
rect 3786 2551 3815 2597
rect 3711 2488 3815 2551
rect 3711 2442 3740 2488
rect 3786 2442 3815 2488
rect 3711 2379 3815 2442
rect 3711 2333 3740 2379
rect 3786 2333 3815 2379
rect 3711 2270 3815 2333
rect 3711 2224 3740 2270
rect 3786 2224 3815 2270
rect 3711 2161 3815 2224
rect 3711 2115 3740 2161
rect 3786 2115 3815 2161
rect 3711 2052 3815 2115
rect 3711 2006 3740 2052
rect 3786 2006 3815 2052
rect 3711 1943 3815 2006
rect 3711 1897 3740 1943
rect 3786 1897 3815 1943
rect 3711 1884 3815 1897
rect 3935 2815 4039 2828
rect 3935 2769 3964 2815
rect 4010 2769 4039 2815
rect 3935 2706 4039 2769
rect 3935 2660 3964 2706
rect 4010 2660 4039 2706
rect 3935 2597 4039 2660
rect 3935 2551 3964 2597
rect 4010 2551 4039 2597
rect 3935 2488 4039 2551
rect 3935 2442 3964 2488
rect 4010 2442 4039 2488
rect 3935 2379 4039 2442
rect 3935 2333 3964 2379
rect 4010 2333 4039 2379
rect 3935 2270 4039 2333
rect 3935 2224 3964 2270
rect 4010 2224 4039 2270
rect 3935 2161 4039 2224
rect 3935 2115 3964 2161
rect 4010 2115 4039 2161
rect 3935 2052 4039 2115
rect 3935 2006 3964 2052
rect 4010 2006 4039 2052
rect 3935 1943 4039 2006
rect 3935 1897 3964 1943
rect 4010 1897 4039 1943
rect 3935 1884 4039 1897
rect 4159 2815 4247 2828
rect 4159 2769 4188 2815
rect 4234 2769 4247 2815
rect 4159 2706 4247 2769
rect 4159 2660 4188 2706
rect 4234 2660 4247 2706
rect 4159 2597 4247 2660
rect 4159 2551 4188 2597
rect 4234 2551 4247 2597
rect 4159 2488 4247 2551
rect 4159 2442 4188 2488
rect 4234 2442 4247 2488
rect 4159 2379 4247 2442
rect 4159 2333 4188 2379
rect 4234 2333 4247 2379
rect 4159 2270 4247 2333
rect 4159 2224 4188 2270
rect 4234 2224 4247 2270
rect 4581 2815 4669 2828
rect 4581 2769 4594 2815
rect 4640 2769 4669 2815
rect 4581 2706 4669 2769
rect 4581 2660 4594 2706
rect 4640 2660 4669 2706
rect 4581 2597 4669 2660
rect 4581 2551 4594 2597
rect 4640 2551 4669 2597
rect 4581 2488 4669 2551
rect 4581 2442 4594 2488
rect 4640 2442 4669 2488
rect 4581 2379 4669 2442
rect 4581 2333 4594 2379
rect 4640 2333 4669 2379
rect 4581 2270 4669 2333
rect 4159 2161 4247 2224
rect 4159 2115 4188 2161
rect 4234 2115 4247 2161
rect 4159 2052 4247 2115
rect 4159 2006 4188 2052
rect 4234 2006 4247 2052
rect 4159 1943 4247 2006
rect 4581 2224 4594 2270
rect 4640 2224 4669 2270
rect 4581 2161 4669 2224
rect 4581 2115 4594 2161
rect 4640 2115 4669 2161
rect 4581 2052 4669 2115
rect 4581 2006 4594 2052
rect 4640 2006 4669 2052
rect 4159 1897 4188 1943
rect 4234 1897 4247 1943
rect 4159 1884 4247 1897
rect 4581 1943 4669 2006
rect 4581 1897 4594 1943
rect 4640 1897 4669 1943
rect 4581 1884 4669 1897
rect 4789 2815 4893 2828
rect 4789 2769 4818 2815
rect 4864 2769 4893 2815
rect 4789 2706 4893 2769
rect 4789 2660 4818 2706
rect 4864 2660 4893 2706
rect 4789 2597 4893 2660
rect 4789 2551 4818 2597
rect 4864 2551 4893 2597
rect 4789 2488 4893 2551
rect 4789 2442 4818 2488
rect 4864 2442 4893 2488
rect 4789 2379 4893 2442
rect 4789 2333 4818 2379
rect 4864 2333 4893 2379
rect 4789 2270 4893 2333
rect 4789 2224 4818 2270
rect 4864 2224 4893 2270
rect 4789 2161 4893 2224
rect 4789 2115 4818 2161
rect 4864 2115 4893 2161
rect 4789 2052 4893 2115
rect 4789 2006 4818 2052
rect 4864 2006 4893 2052
rect 4789 1943 4893 2006
rect 4789 1897 4818 1943
rect 4864 1897 4893 1943
rect 4789 1884 4893 1897
rect 5013 2815 5117 2828
rect 5013 2769 5042 2815
rect 5088 2769 5117 2815
rect 5013 2706 5117 2769
rect 5013 2660 5042 2706
rect 5088 2660 5117 2706
rect 5013 2597 5117 2660
rect 5013 2551 5042 2597
rect 5088 2551 5117 2597
rect 5013 2488 5117 2551
rect 5013 2442 5042 2488
rect 5088 2442 5117 2488
rect 5013 2379 5117 2442
rect 5013 2333 5042 2379
rect 5088 2333 5117 2379
rect 5013 2270 5117 2333
rect 5013 2224 5042 2270
rect 5088 2224 5117 2270
rect 5013 2161 5117 2224
rect 5013 2115 5042 2161
rect 5088 2115 5117 2161
rect 5013 2052 5117 2115
rect 5013 2006 5042 2052
rect 5088 2006 5117 2052
rect 5013 1943 5117 2006
rect 5013 1897 5042 1943
rect 5088 1897 5117 1943
rect 5013 1884 5117 1897
rect 5237 2815 5341 2828
rect 5237 2769 5266 2815
rect 5312 2769 5341 2815
rect 5237 2706 5341 2769
rect 5237 2660 5266 2706
rect 5312 2660 5341 2706
rect 5237 2597 5341 2660
rect 5237 2551 5266 2597
rect 5312 2551 5341 2597
rect 5237 2488 5341 2551
rect 5237 2442 5266 2488
rect 5312 2442 5341 2488
rect 5237 2379 5341 2442
rect 5237 2333 5266 2379
rect 5312 2333 5341 2379
rect 5237 2270 5341 2333
rect 5237 2224 5266 2270
rect 5312 2224 5341 2270
rect 5237 2161 5341 2224
rect 5237 2115 5266 2161
rect 5312 2115 5341 2161
rect 5237 2052 5341 2115
rect 5237 2006 5266 2052
rect 5312 2006 5341 2052
rect 5237 1943 5341 2006
rect 5237 1897 5266 1943
rect 5312 1897 5341 1943
rect 5237 1884 5341 1897
rect 5461 2815 5565 2828
rect 5461 2769 5490 2815
rect 5536 2769 5565 2815
rect 5461 2706 5565 2769
rect 5461 2660 5490 2706
rect 5536 2660 5565 2706
rect 5461 2597 5565 2660
rect 5461 2551 5490 2597
rect 5536 2551 5565 2597
rect 5461 2488 5565 2551
rect 5461 2442 5490 2488
rect 5536 2442 5565 2488
rect 5461 2379 5565 2442
rect 5461 2333 5490 2379
rect 5536 2333 5565 2379
rect 5461 2270 5565 2333
rect 5461 2224 5490 2270
rect 5536 2224 5565 2270
rect 5461 2161 5565 2224
rect 5461 2115 5490 2161
rect 5536 2115 5565 2161
rect 5461 2052 5565 2115
rect 5461 2006 5490 2052
rect 5536 2006 5565 2052
rect 5461 1943 5565 2006
rect 5461 1897 5490 1943
rect 5536 1897 5565 1943
rect 5461 1884 5565 1897
rect 5685 2815 5789 2828
rect 5685 2769 5714 2815
rect 5760 2769 5789 2815
rect 5685 2706 5789 2769
rect 5685 2660 5714 2706
rect 5760 2660 5789 2706
rect 5685 2597 5789 2660
rect 5685 2551 5714 2597
rect 5760 2551 5789 2597
rect 5685 2488 5789 2551
rect 5685 2442 5714 2488
rect 5760 2442 5789 2488
rect 5685 2379 5789 2442
rect 5685 2333 5714 2379
rect 5760 2333 5789 2379
rect 5685 2270 5789 2333
rect 5685 2224 5714 2270
rect 5760 2224 5789 2270
rect 5685 2161 5789 2224
rect 5685 2115 5714 2161
rect 5760 2115 5789 2161
rect 5685 2052 5789 2115
rect 5685 2006 5714 2052
rect 5760 2006 5789 2052
rect 5685 1943 5789 2006
rect 5685 1897 5714 1943
rect 5760 1897 5789 1943
rect 5685 1884 5789 1897
rect 5909 2815 6013 2828
rect 5909 2769 5938 2815
rect 5984 2769 6013 2815
rect 5909 2706 6013 2769
rect 5909 2660 5938 2706
rect 5984 2660 6013 2706
rect 5909 2597 6013 2660
rect 5909 2551 5938 2597
rect 5984 2551 6013 2597
rect 5909 2488 6013 2551
rect 5909 2442 5938 2488
rect 5984 2442 6013 2488
rect 5909 2379 6013 2442
rect 5909 2333 5938 2379
rect 5984 2333 6013 2379
rect 5909 2270 6013 2333
rect 5909 2224 5938 2270
rect 5984 2224 6013 2270
rect 5909 2161 6013 2224
rect 5909 2115 5938 2161
rect 5984 2115 6013 2161
rect 5909 2052 6013 2115
rect 5909 2006 5938 2052
rect 5984 2006 6013 2052
rect 5909 1943 6013 2006
rect 5909 1897 5938 1943
rect 5984 1897 6013 1943
rect 5909 1884 6013 1897
rect 6133 2815 6237 2828
rect 6133 2769 6162 2815
rect 6208 2769 6237 2815
rect 6133 2706 6237 2769
rect 6133 2660 6162 2706
rect 6208 2660 6237 2706
rect 6133 2597 6237 2660
rect 6133 2551 6162 2597
rect 6208 2551 6237 2597
rect 6133 2488 6237 2551
rect 6133 2442 6162 2488
rect 6208 2442 6237 2488
rect 6133 2379 6237 2442
rect 6133 2333 6162 2379
rect 6208 2333 6237 2379
rect 6133 2270 6237 2333
rect 6133 2224 6162 2270
rect 6208 2224 6237 2270
rect 6133 2161 6237 2224
rect 6133 2115 6162 2161
rect 6208 2115 6237 2161
rect 6133 2052 6237 2115
rect 6133 2006 6162 2052
rect 6208 2006 6237 2052
rect 6133 1943 6237 2006
rect 6133 1897 6162 1943
rect 6208 1897 6237 1943
rect 6133 1884 6237 1897
rect 6357 2815 6461 2828
rect 6357 2769 6386 2815
rect 6432 2769 6461 2815
rect 6357 2706 6461 2769
rect 6357 2660 6386 2706
rect 6432 2660 6461 2706
rect 6357 2597 6461 2660
rect 6357 2551 6386 2597
rect 6432 2551 6461 2597
rect 6357 2488 6461 2551
rect 6357 2442 6386 2488
rect 6432 2442 6461 2488
rect 6357 2379 6461 2442
rect 6357 2333 6386 2379
rect 6432 2333 6461 2379
rect 6357 2270 6461 2333
rect 6357 2224 6386 2270
rect 6432 2224 6461 2270
rect 6357 2161 6461 2224
rect 6357 2115 6386 2161
rect 6432 2115 6461 2161
rect 6357 2052 6461 2115
rect 6357 2006 6386 2052
rect 6432 2006 6461 2052
rect 6357 1943 6461 2006
rect 6357 1897 6386 1943
rect 6432 1897 6461 1943
rect 6357 1884 6461 1897
rect 6581 2815 6685 2828
rect 6581 2769 6610 2815
rect 6656 2769 6685 2815
rect 6581 2706 6685 2769
rect 6581 2660 6610 2706
rect 6656 2660 6685 2706
rect 6581 2597 6685 2660
rect 6581 2551 6610 2597
rect 6656 2551 6685 2597
rect 6581 2488 6685 2551
rect 6581 2442 6610 2488
rect 6656 2442 6685 2488
rect 6581 2379 6685 2442
rect 6581 2333 6610 2379
rect 6656 2333 6685 2379
rect 6581 2270 6685 2333
rect 6581 2224 6610 2270
rect 6656 2224 6685 2270
rect 6581 2161 6685 2224
rect 6581 2115 6610 2161
rect 6656 2115 6685 2161
rect 6581 2052 6685 2115
rect 6581 2006 6610 2052
rect 6656 2006 6685 2052
rect 6581 1943 6685 2006
rect 6581 1897 6610 1943
rect 6656 1897 6685 1943
rect 6581 1884 6685 1897
rect 6805 2815 6893 2828
rect 6805 2769 6834 2815
rect 6880 2769 6893 2815
rect 6805 2706 6893 2769
rect 6805 2660 6834 2706
rect 6880 2660 6893 2706
rect 6805 2597 6893 2660
rect 6805 2551 6834 2597
rect 6880 2551 6893 2597
rect 6805 2488 6893 2551
rect 6805 2442 6834 2488
rect 6880 2442 6893 2488
rect 6805 2379 6893 2442
rect 6805 2333 6834 2379
rect 6880 2333 6893 2379
rect 6805 2270 6893 2333
rect 6805 2224 6834 2270
rect 6880 2224 6893 2270
rect 6805 2161 6893 2224
rect 6805 2115 6834 2161
rect 6880 2115 6893 2161
rect 6805 2052 6893 2115
rect 6805 2006 6834 2052
rect 6880 2006 6893 2052
rect 6805 1943 6893 2006
rect 6805 1897 6834 1943
rect 6880 1897 6893 1943
rect 6805 1884 6893 1897
rect 421 1284 509 1297
rect 421 1238 434 1284
rect 480 1238 509 1284
rect 421 1157 509 1238
rect 421 1111 434 1157
rect 480 1111 509 1157
rect 421 1030 509 1111
rect 421 984 434 1030
rect 480 984 509 1030
rect 421 902 509 984
rect 421 856 434 902
rect 480 856 509 902
rect 421 843 509 856
rect 629 1284 733 1297
rect 629 1238 658 1284
rect 704 1238 733 1284
rect 629 1157 733 1238
rect 629 1111 658 1157
rect 704 1111 733 1157
rect 629 1030 733 1111
rect 629 984 658 1030
rect 704 984 733 1030
rect 629 902 733 984
rect 629 856 658 902
rect 704 856 733 902
rect 629 843 733 856
rect 853 1284 941 1297
rect 853 1238 882 1284
rect 928 1238 941 1284
rect 853 1157 941 1238
rect 853 1111 882 1157
rect 928 1111 941 1157
rect 853 1030 941 1111
rect 853 984 882 1030
rect 928 984 941 1030
rect 853 902 941 984
rect 853 856 882 902
rect 928 856 941 902
rect 853 843 941 856
rect 1093 1284 1181 1297
rect 1093 1238 1106 1284
rect 1152 1238 1181 1284
rect 1093 1157 1181 1238
rect 1093 1111 1106 1157
rect 1152 1111 1181 1157
rect 1093 1030 1181 1111
rect 1093 984 1106 1030
rect 1152 984 1181 1030
rect 1093 902 1181 984
rect 1093 856 1106 902
rect 1152 856 1181 902
rect 1093 843 1181 856
rect 1301 1284 1389 1297
rect 1301 1238 1330 1284
rect 1376 1238 1389 1284
rect 1301 1157 1389 1238
rect 1301 1111 1330 1157
rect 1376 1111 1389 1157
rect 1301 1030 1389 1111
rect 1301 984 1330 1030
rect 1376 984 1389 1030
rect 1301 902 1389 984
rect 1301 856 1330 902
rect 1376 856 1389 902
rect 1301 843 1389 856
rect 1600 1284 1688 1297
rect 1600 1238 1613 1284
rect 1659 1238 1688 1284
rect 1600 1157 1688 1238
rect 1600 1111 1613 1157
rect 1659 1111 1688 1157
rect 1600 1030 1688 1111
rect 1600 984 1613 1030
rect 1659 984 1688 1030
rect 1600 902 1688 984
rect 1600 856 1613 902
rect 1659 856 1688 902
rect 1600 843 1688 856
rect 1808 1284 1896 1297
rect 1808 1238 1837 1284
rect 1883 1238 1896 1284
rect 1808 1157 1896 1238
rect 1808 1111 1837 1157
rect 1883 1111 1896 1157
rect 1808 1035 1896 1111
rect 3205 1398 3293 1411
rect 3205 1352 3218 1398
rect 3264 1352 3293 1398
rect 2286 1284 2374 1297
rect 2286 1238 2299 1284
rect 2345 1238 2374 1284
rect 2286 1157 2374 1238
rect 2286 1111 2299 1157
rect 2345 1111 2374 1157
rect 2286 1035 2374 1111
rect 1808 1030 2036 1035
rect 1808 984 1837 1030
rect 1883 1022 2036 1030
rect 1883 984 1961 1022
rect 1808 976 1961 984
rect 2007 976 2036 1022
rect 1808 902 2036 976
rect 1808 856 1837 902
rect 1883 856 1961 902
rect 2007 856 2036 902
rect 1808 843 2036 856
rect 2156 1030 2374 1035
rect 2156 1022 2299 1030
rect 2156 976 2185 1022
rect 2231 984 2299 1022
rect 2345 984 2374 1030
rect 2231 976 2374 984
rect 2156 902 2374 976
rect 2156 856 2185 902
rect 2231 856 2299 902
rect 2345 856 2374 902
rect 2156 843 2374 856
rect 2494 1284 2582 1297
rect 2494 1238 2523 1284
rect 2569 1238 2582 1284
rect 2494 1157 2582 1238
rect 2494 1111 2523 1157
rect 2569 1111 2582 1157
rect 2494 1030 2582 1111
rect 2494 984 2523 1030
rect 2569 984 2582 1030
rect 2494 902 2582 984
rect 2494 856 2523 902
rect 2569 856 2582 902
rect 2494 843 2582 856
rect 2734 1284 2822 1297
rect 2734 1238 2747 1284
rect 2793 1238 2822 1284
rect 2734 1157 2822 1238
rect 2734 1111 2747 1157
rect 2793 1111 2822 1157
rect 2734 1030 2822 1111
rect 2734 984 2747 1030
rect 2793 984 2822 1030
rect 2734 902 2822 984
rect 2734 856 2747 902
rect 2793 856 2822 902
rect 2734 843 2822 856
rect 2942 1284 3030 1297
rect 2942 1238 2971 1284
rect 3017 1238 3030 1284
rect 2942 1157 3030 1238
rect 2942 1111 2971 1157
rect 3017 1111 3030 1157
rect 2942 1030 3030 1111
rect 2942 984 2971 1030
rect 3017 984 3030 1030
rect 2942 902 3030 984
rect 2942 856 2971 902
rect 3017 856 3030 902
rect 2942 843 3030 856
rect 3205 1274 3293 1352
rect 3205 1228 3218 1274
rect 3264 1228 3293 1274
rect 3205 1150 3293 1228
rect 3205 1104 3218 1150
rect 3264 1104 3293 1150
rect 3205 1026 3293 1104
rect 3205 980 3218 1026
rect 3264 980 3293 1026
rect 3205 902 3293 980
rect 3205 856 3218 902
rect 3264 856 3293 902
rect 3205 843 3293 856
rect 3413 1398 3517 1411
rect 3413 1352 3442 1398
rect 3488 1352 3517 1398
rect 3413 1274 3517 1352
rect 3413 1228 3442 1274
rect 3488 1228 3517 1274
rect 3413 1150 3517 1228
rect 3413 1104 3442 1150
rect 3488 1104 3517 1150
rect 3413 1026 3517 1104
rect 3413 980 3442 1026
rect 3488 980 3517 1026
rect 3413 902 3517 980
rect 3413 856 3442 902
rect 3488 856 3517 902
rect 3413 843 3517 856
rect 3637 1398 3725 1411
rect 3637 1352 3666 1398
rect 3712 1352 3725 1398
rect 3637 1274 3725 1352
rect 3637 1228 3666 1274
rect 3712 1228 3725 1274
rect 3637 1150 3725 1228
rect 3637 1104 3666 1150
rect 3712 1104 3725 1150
rect 3637 1026 3725 1104
rect 3637 980 3666 1026
rect 3712 980 3725 1026
rect 3637 902 3725 980
rect 3637 856 3666 902
rect 3712 856 3725 902
rect 3637 843 3725 856
rect 3862 1284 3950 1297
rect 3862 1238 3875 1284
rect 3921 1238 3950 1284
rect 3862 1157 3950 1238
rect 3862 1111 3875 1157
rect 3921 1111 3950 1157
rect 3862 1030 3950 1111
rect 3862 984 3875 1030
rect 3921 984 3950 1030
rect 3862 902 3950 984
rect 3862 856 3875 902
rect 3921 856 3950 902
rect 3862 843 3950 856
rect 4070 1284 4174 1297
rect 4070 1238 4099 1284
rect 4145 1238 4174 1284
rect 4070 1157 4174 1238
rect 4070 1111 4099 1157
rect 4145 1111 4174 1157
rect 4070 1030 4174 1111
rect 4070 984 4099 1030
rect 4145 984 4174 1030
rect 4070 902 4174 984
rect 4070 856 4099 902
rect 4145 856 4174 902
rect 4070 843 4174 856
rect 4294 1284 4510 1297
rect 4294 1238 4323 1284
rect 4369 1238 4435 1284
rect 4481 1238 4510 1284
rect 4294 1164 4510 1238
rect 4294 1157 4435 1164
rect 4294 1111 4323 1157
rect 4369 1118 4435 1157
rect 4481 1118 4510 1164
rect 4369 1111 4510 1118
rect 4294 1105 4510 1111
rect 4630 1284 4842 1297
rect 4630 1238 4659 1284
rect 4705 1238 4767 1284
rect 4813 1238 4842 1284
rect 4630 1164 4842 1238
rect 4630 1118 4659 1164
rect 4705 1156 4842 1164
rect 4705 1118 4767 1156
rect 4630 1110 4767 1118
rect 4813 1110 4842 1156
rect 4630 1105 4842 1110
rect 4294 1030 4382 1105
rect 4294 984 4323 1030
rect 4369 984 4382 1030
rect 4294 902 4382 984
rect 4294 856 4323 902
rect 4369 856 4382 902
rect 4294 843 4382 856
rect 4754 1029 4842 1105
rect 4754 983 4767 1029
rect 4813 983 4842 1029
rect 4754 902 4842 983
rect 4754 856 4767 902
rect 4813 856 4842 902
rect 4754 843 4842 856
rect 4962 1284 5050 1297
rect 4962 1238 4991 1284
rect 5037 1238 5050 1284
rect 4962 1156 5050 1238
rect 4962 1110 4991 1156
rect 5037 1110 5050 1156
rect 4962 1029 5050 1110
rect 4962 983 4991 1029
rect 5037 983 5050 1029
rect 4962 902 5050 983
rect 4962 856 4991 902
rect 5037 856 5050 902
rect 4962 843 5050 856
rect 5219 1270 5307 1283
rect 5219 1224 5232 1270
rect 5278 1224 5307 1270
rect 5219 1148 5307 1224
rect 5219 1102 5232 1148
rect 5278 1102 5307 1148
rect 5219 1025 5307 1102
rect 5219 979 5232 1025
rect 5278 979 5307 1025
rect 5219 902 5307 979
rect 5219 856 5232 902
rect 5278 856 5307 902
rect 5219 843 5307 856
rect 5427 1270 5531 1283
rect 5427 1224 5456 1270
rect 5502 1224 5531 1270
rect 5427 1148 5531 1224
rect 5427 1102 5456 1148
rect 5502 1102 5531 1148
rect 5427 1025 5531 1102
rect 5427 979 5456 1025
rect 5502 979 5531 1025
rect 5427 902 5531 979
rect 5427 856 5456 902
rect 5502 856 5531 902
rect 5427 843 5531 856
rect 5651 1270 5755 1283
rect 5651 1224 5680 1270
rect 5726 1224 5755 1270
rect 5651 1148 5755 1224
rect 5651 1102 5680 1148
rect 5726 1102 5755 1148
rect 5651 1025 5755 1102
rect 5651 979 5680 1025
rect 5726 979 5755 1025
rect 5651 902 5755 979
rect 5651 856 5680 902
rect 5726 856 5755 902
rect 5651 843 5755 856
rect 5875 1270 5979 1283
rect 5875 1224 5904 1270
rect 5950 1224 5979 1270
rect 5875 1148 5979 1224
rect 5875 1102 5904 1148
rect 5950 1102 5979 1148
rect 5875 1025 5979 1102
rect 5875 979 5904 1025
rect 5950 979 5979 1025
rect 5875 902 5979 979
rect 5875 856 5904 902
rect 5950 856 5979 902
rect 5875 843 5979 856
rect 6099 1270 6203 1283
rect 6099 1224 6128 1270
rect 6174 1224 6203 1270
rect 6099 1148 6203 1224
rect 6099 1102 6128 1148
rect 6174 1102 6203 1148
rect 6099 1025 6203 1102
rect 6099 979 6128 1025
rect 6174 979 6203 1025
rect 6099 902 6203 979
rect 6099 856 6128 902
rect 6174 856 6203 902
rect 6099 843 6203 856
rect 6323 1270 6427 1283
rect 6323 1224 6352 1270
rect 6398 1224 6427 1270
rect 6323 1148 6427 1224
rect 6323 1102 6352 1148
rect 6398 1102 6427 1148
rect 6323 1025 6427 1102
rect 6323 979 6352 1025
rect 6398 979 6427 1025
rect 6323 902 6427 979
rect 6323 856 6352 902
rect 6398 856 6427 902
rect 6323 843 6427 856
rect 6547 1270 6651 1283
rect 6547 1224 6576 1270
rect 6622 1224 6651 1270
rect 6547 1148 6651 1224
rect 6547 1102 6576 1148
rect 6622 1102 6651 1148
rect 6547 1025 6651 1102
rect 6547 979 6576 1025
rect 6622 979 6651 1025
rect 6547 902 6651 979
rect 6547 856 6576 902
rect 6622 856 6651 902
rect 6547 843 6651 856
rect 6771 1270 6859 1283
rect 6771 1224 6800 1270
rect 6846 1224 6859 1270
rect 6771 1148 6859 1224
rect 6771 1102 6800 1148
rect 6846 1102 6859 1148
rect 6771 1025 6859 1102
rect 6771 979 6800 1025
rect 6846 979 6859 1025
rect 6771 902 6859 979
rect 6771 856 6800 902
rect 6846 856 6859 902
rect 6771 843 6859 856
<< ndiffc >>
rect 133 438 179 484
rect 133 274 179 320
<< mvndiffc >>
rect 177 3555 223 3601
rect 177 3446 223 3492
rect 177 3337 223 3383
rect 177 3227 223 3273
rect 401 3555 447 3601
rect 401 3446 447 3492
rect 401 3337 447 3383
rect 401 3227 447 3273
rect 625 3555 671 3601
rect 625 3446 671 3492
rect 625 3337 671 3383
rect 625 3227 671 3273
rect 849 3555 895 3601
rect 849 3446 895 3492
rect 849 3337 895 3383
rect 849 3227 895 3273
rect 1948 3539 1994 3585
rect 1948 3435 1994 3481
rect 1948 3331 1994 3377
rect 1948 3227 1994 3273
rect 2172 3539 2218 3585
rect 2172 3435 2218 3481
rect 2172 3331 2218 3377
rect 2172 3227 2218 3273
rect 2396 3539 2442 3585
rect 2396 3435 2442 3481
rect 2396 3331 2442 3377
rect 2396 3227 2442 3273
rect 2620 3539 2666 3585
rect 2620 3435 2666 3481
rect 2620 3331 2666 3377
rect 2620 3227 2666 3273
rect 2844 3539 2890 3585
rect 2844 3435 2890 3481
rect 2844 3331 2890 3377
rect 2844 3227 2890 3273
rect 3068 3539 3114 3585
rect 3068 3435 3114 3481
rect 3068 3331 3114 3377
rect 3068 3227 3114 3273
rect 3292 3539 3338 3585
rect 3292 3435 3338 3481
rect 3292 3331 3338 3377
rect 3292 3227 3338 3273
rect 3516 3539 3562 3585
rect 3516 3435 3562 3481
rect 3516 3331 3562 3377
rect 3516 3227 3562 3273
rect 3740 3539 3786 3585
rect 3740 3435 3786 3481
rect 3740 3331 3786 3377
rect 3740 3227 3786 3273
rect 3964 3539 4010 3585
rect 3964 3435 4010 3481
rect 3964 3331 4010 3377
rect 3964 3227 4010 3273
rect 4188 3539 4234 3585
rect 4188 3435 4234 3481
rect 4188 3331 4234 3377
rect 4188 3227 4234 3273
rect 4594 3539 4640 3585
rect 4594 3435 4640 3481
rect 4594 3331 4640 3377
rect 4594 3227 4640 3273
rect 4818 3539 4864 3585
rect 4818 3435 4864 3481
rect 4818 3331 4864 3377
rect 4818 3227 4864 3273
rect 5042 3539 5088 3585
rect 5042 3435 5088 3481
rect 5042 3331 5088 3377
rect 5042 3227 5088 3273
rect 5266 3539 5312 3585
rect 5266 3435 5312 3481
rect 5266 3331 5312 3377
rect 5266 3227 5312 3273
rect 5490 3539 5536 3585
rect 5490 3435 5536 3481
rect 5490 3331 5536 3377
rect 5490 3227 5536 3273
rect 5714 3539 5760 3585
rect 5714 3435 5760 3481
rect 5714 3331 5760 3377
rect 5714 3227 5760 3273
rect 5938 3539 5984 3585
rect 5938 3435 5984 3481
rect 5938 3331 5984 3377
rect 5938 3227 5984 3273
rect 6162 3539 6208 3585
rect 6162 3435 6208 3481
rect 6162 3331 6208 3377
rect 6162 3227 6208 3273
rect 6386 3539 6432 3585
rect 6386 3435 6432 3481
rect 6386 3331 6432 3377
rect 6386 3227 6432 3273
rect 6610 3539 6656 3585
rect 6610 3435 6656 3481
rect 6610 3331 6656 3377
rect 6610 3227 6656 3273
rect 6834 3539 6880 3585
rect 6834 3435 6880 3481
rect 6834 3331 6880 3377
rect 6834 3227 6880 3273
rect 1613 504 1659 550
rect 1106 428 1152 474
rect 434 346 480 392
rect 434 226 480 272
rect 658 346 704 392
rect 658 226 704 272
rect 882 346 928 392
rect 1106 308 1152 354
rect 1330 428 1376 474
rect 1330 308 1376 354
rect 1613 377 1659 423
rect 882 226 928 272
rect 1613 250 1659 296
rect 1613 122 1659 168
rect 1837 504 1883 550
rect 1837 377 1883 423
rect 2075 505 2121 551
rect 2075 385 2121 431
rect 2299 505 2345 551
rect 2299 385 2345 431
rect 2523 505 2569 551
rect 2523 385 2569 431
rect 2747 505 2793 551
rect 2747 385 2793 431
rect 2971 505 3017 551
rect 2971 385 3017 431
rect 3218 505 3264 551
rect 1837 250 1883 296
rect 1837 122 1883 168
rect 3218 337 3264 383
rect 3442 505 3488 551
rect 3442 337 3488 383
rect 3666 505 3712 551
rect 3666 337 3712 383
rect 3875 504 3921 550
rect 3875 377 3921 423
rect 3875 250 3921 296
rect 3875 122 3921 168
rect 4099 504 4145 550
rect 4099 377 4145 423
rect 4099 250 4145 296
rect 4099 122 4145 168
rect 4323 504 4369 550
rect 5232 500 5278 546
rect 4323 377 4369 423
rect 4323 250 4369 296
rect 4543 381 4589 427
rect 4543 261 4589 307
rect 4767 381 4813 427
rect 4767 261 4813 307
rect 4991 381 5037 427
rect 5232 394 5278 440
rect 5456 500 5502 546
rect 5456 394 5502 440
rect 5680 500 5726 546
rect 5680 394 5726 440
rect 5904 500 5950 546
rect 5904 394 5950 440
rect 6128 500 6174 546
rect 6128 394 6174 440
rect 6352 500 6398 546
rect 6352 394 6398 440
rect 6576 500 6622 546
rect 6576 394 6622 440
rect 6800 500 6846 546
rect 6800 394 6846 440
rect 4991 261 5037 307
rect 4323 122 4369 168
<< mvpdiffc >>
rect 1948 2769 1994 2815
rect 1948 2660 1994 2706
rect 1948 2551 1994 2597
rect 1948 2442 1994 2488
rect 177 2321 223 2367
rect 177 2215 223 2261
rect 177 2109 223 2155
rect 177 2003 223 2049
rect 177 1897 223 1943
rect 401 2321 447 2367
rect 401 2215 447 2261
rect 401 2109 447 2155
rect 401 2003 447 2049
rect 401 1897 447 1943
rect 625 2321 671 2367
rect 625 2215 671 2261
rect 625 2109 671 2155
rect 625 2003 671 2049
rect 625 1897 671 1943
rect 849 2321 895 2367
rect 849 2215 895 2261
rect 849 2109 895 2155
rect 849 2003 895 2049
rect 849 1897 895 1943
rect 1073 2321 1119 2367
rect 1073 2215 1119 2261
rect 1073 2109 1119 2155
rect 1073 2003 1119 2049
rect 1073 1897 1119 1943
rect 1297 2321 1343 2367
rect 1297 2215 1343 2261
rect 1297 2109 1343 2155
rect 1297 2003 1343 2049
rect 1297 1897 1343 1943
rect 1521 2321 1567 2367
rect 1948 2333 1994 2379
rect 1521 2215 1567 2261
rect 1521 2109 1567 2155
rect 1521 2003 1567 2049
rect 1948 2224 1994 2270
rect 1948 2115 1994 2161
rect 1948 2006 1994 2052
rect 1521 1897 1567 1943
rect 1948 1897 1994 1943
rect 2172 2769 2218 2815
rect 2172 2660 2218 2706
rect 2172 2551 2218 2597
rect 2172 2442 2218 2488
rect 2172 2333 2218 2379
rect 2172 2224 2218 2270
rect 2172 2115 2218 2161
rect 2172 2006 2218 2052
rect 2172 1897 2218 1943
rect 2396 2769 2442 2815
rect 2396 2660 2442 2706
rect 2396 2551 2442 2597
rect 2396 2442 2442 2488
rect 2396 2333 2442 2379
rect 2396 2224 2442 2270
rect 2396 2115 2442 2161
rect 2396 2006 2442 2052
rect 2396 1897 2442 1943
rect 2620 2769 2666 2815
rect 2620 2660 2666 2706
rect 2620 2551 2666 2597
rect 2620 2442 2666 2488
rect 2620 2333 2666 2379
rect 2620 2224 2666 2270
rect 2620 2115 2666 2161
rect 2620 2006 2666 2052
rect 2620 1897 2666 1943
rect 2844 2769 2890 2815
rect 2844 2660 2890 2706
rect 2844 2551 2890 2597
rect 2844 2442 2890 2488
rect 2844 2333 2890 2379
rect 2844 2224 2890 2270
rect 2844 2115 2890 2161
rect 2844 2006 2890 2052
rect 2844 1897 2890 1943
rect 3068 2769 3114 2815
rect 3068 2660 3114 2706
rect 3068 2551 3114 2597
rect 3068 2442 3114 2488
rect 3068 2333 3114 2379
rect 3068 2224 3114 2270
rect 3068 2115 3114 2161
rect 3068 2006 3114 2052
rect 3068 1897 3114 1943
rect 3292 2769 3338 2815
rect 3292 2660 3338 2706
rect 3292 2551 3338 2597
rect 3292 2442 3338 2488
rect 3292 2333 3338 2379
rect 3292 2224 3338 2270
rect 3292 2115 3338 2161
rect 3292 2006 3338 2052
rect 3292 1897 3338 1943
rect 3516 2769 3562 2815
rect 3516 2660 3562 2706
rect 3516 2551 3562 2597
rect 3516 2442 3562 2488
rect 3516 2333 3562 2379
rect 3516 2224 3562 2270
rect 3516 2115 3562 2161
rect 3516 2006 3562 2052
rect 3516 1897 3562 1943
rect 3740 2769 3786 2815
rect 3740 2660 3786 2706
rect 3740 2551 3786 2597
rect 3740 2442 3786 2488
rect 3740 2333 3786 2379
rect 3740 2224 3786 2270
rect 3740 2115 3786 2161
rect 3740 2006 3786 2052
rect 3740 1897 3786 1943
rect 3964 2769 4010 2815
rect 3964 2660 4010 2706
rect 3964 2551 4010 2597
rect 3964 2442 4010 2488
rect 3964 2333 4010 2379
rect 3964 2224 4010 2270
rect 3964 2115 4010 2161
rect 3964 2006 4010 2052
rect 3964 1897 4010 1943
rect 4188 2769 4234 2815
rect 4188 2660 4234 2706
rect 4188 2551 4234 2597
rect 4188 2442 4234 2488
rect 4188 2333 4234 2379
rect 4188 2224 4234 2270
rect 4594 2769 4640 2815
rect 4594 2660 4640 2706
rect 4594 2551 4640 2597
rect 4594 2442 4640 2488
rect 4594 2333 4640 2379
rect 4188 2115 4234 2161
rect 4188 2006 4234 2052
rect 4594 2224 4640 2270
rect 4594 2115 4640 2161
rect 4594 2006 4640 2052
rect 4188 1897 4234 1943
rect 4594 1897 4640 1943
rect 4818 2769 4864 2815
rect 4818 2660 4864 2706
rect 4818 2551 4864 2597
rect 4818 2442 4864 2488
rect 4818 2333 4864 2379
rect 4818 2224 4864 2270
rect 4818 2115 4864 2161
rect 4818 2006 4864 2052
rect 4818 1897 4864 1943
rect 5042 2769 5088 2815
rect 5042 2660 5088 2706
rect 5042 2551 5088 2597
rect 5042 2442 5088 2488
rect 5042 2333 5088 2379
rect 5042 2224 5088 2270
rect 5042 2115 5088 2161
rect 5042 2006 5088 2052
rect 5042 1897 5088 1943
rect 5266 2769 5312 2815
rect 5266 2660 5312 2706
rect 5266 2551 5312 2597
rect 5266 2442 5312 2488
rect 5266 2333 5312 2379
rect 5266 2224 5312 2270
rect 5266 2115 5312 2161
rect 5266 2006 5312 2052
rect 5266 1897 5312 1943
rect 5490 2769 5536 2815
rect 5490 2660 5536 2706
rect 5490 2551 5536 2597
rect 5490 2442 5536 2488
rect 5490 2333 5536 2379
rect 5490 2224 5536 2270
rect 5490 2115 5536 2161
rect 5490 2006 5536 2052
rect 5490 1897 5536 1943
rect 5714 2769 5760 2815
rect 5714 2660 5760 2706
rect 5714 2551 5760 2597
rect 5714 2442 5760 2488
rect 5714 2333 5760 2379
rect 5714 2224 5760 2270
rect 5714 2115 5760 2161
rect 5714 2006 5760 2052
rect 5714 1897 5760 1943
rect 5938 2769 5984 2815
rect 5938 2660 5984 2706
rect 5938 2551 5984 2597
rect 5938 2442 5984 2488
rect 5938 2333 5984 2379
rect 5938 2224 5984 2270
rect 5938 2115 5984 2161
rect 5938 2006 5984 2052
rect 5938 1897 5984 1943
rect 6162 2769 6208 2815
rect 6162 2660 6208 2706
rect 6162 2551 6208 2597
rect 6162 2442 6208 2488
rect 6162 2333 6208 2379
rect 6162 2224 6208 2270
rect 6162 2115 6208 2161
rect 6162 2006 6208 2052
rect 6162 1897 6208 1943
rect 6386 2769 6432 2815
rect 6386 2660 6432 2706
rect 6386 2551 6432 2597
rect 6386 2442 6432 2488
rect 6386 2333 6432 2379
rect 6386 2224 6432 2270
rect 6386 2115 6432 2161
rect 6386 2006 6432 2052
rect 6386 1897 6432 1943
rect 6610 2769 6656 2815
rect 6610 2660 6656 2706
rect 6610 2551 6656 2597
rect 6610 2442 6656 2488
rect 6610 2333 6656 2379
rect 6610 2224 6656 2270
rect 6610 2115 6656 2161
rect 6610 2006 6656 2052
rect 6610 1897 6656 1943
rect 6834 2769 6880 2815
rect 6834 2660 6880 2706
rect 6834 2551 6880 2597
rect 6834 2442 6880 2488
rect 6834 2333 6880 2379
rect 6834 2224 6880 2270
rect 6834 2115 6880 2161
rect 6834 2006 6880 2052
rect 6834 1897 6880 1943
rect 434 1238 480 1284
rect 434 1111 480 1157
rect 434 984 480 1030
rect 434 856 480 902
rect 658 1238 704 1284
rect 658 1111 704 1157
rect 658 984 704 1030
rect 658 856 704 902
rect 882 1238 928 1284
rect 882 1111 928 1157
rect 882 984 928 1030
rect 882 856 928 902
rect 1106 1238 1152 1284
rect 1106 1111 1152 1157
rect 1106 984 1152 1030
rect 1106 856 1152 902
rect 1330 1238 1376 1284
rect 1330 1111 1376 1157
rect 1330 984 1376 1030
rect 1330 856 1376 902
rect 1613 1238 1659 1284
rect 1613 1111 1659 1157
rect 1613 984 1659 1030
rect 1613 856 1659 902
rect 1837 1238 1883 1284
rect 1837 1111 1883 1157
rect 3218 1352 3264 1398
rect 2299 1238 2345 1284
rect 2299 1111 2345 1157
rect 1837 984 1883 1030
rect 1961 976 2007 1022
rect 1837 856 1883 902
rect 1961 856 2007 902
rect 2185 976 2231 1022
rect 2299 984 2345 1030
rect 2185 856 2231 902
rect 2299 856 2345 902
rect 2523 1238 2569 1284
rect 2523 1111 2569 1157
rect 2523 984 2569 1030
rect 2523 856 2569 902
rect 2747 1238 2793 1284
rect 2747 1111 2793 1157
rect 2747 984 2793 1030
rect 2747 856 2793 902
rect 2971 1238 3017 1284
rect 2971 1111 3017 1157
rect 2971 984 3017 1030
rect 2971 856 3017 902
rect 3218 1228 3264 1274
rect 3218 1104 3264 1150
rect 3218 980 3264 1026
rect 3218 856 3264 902
rect 3442 1352 3488 1398
rect 3442 1228 3488 1274
rect 3442 1104 3488 1150
rect 3442 980 3488 1026
rect 3442 856 3488 902
rect 3666 1352 3712 1398
rect 3666 1228 3712 1274
rect 3666 1104 3712 1150
rect 3666 980 3712 1026
rect 3666 856 3712 902
rect 3875 1238 3921 1284
rect 3875 1111 3921 1157
rect 3875 984 3921 1030
rect 3875 856 3921 902
rect 4099 1238 4145 1284
rect 4099 1111 4145 1157
rect 4099 984 4145 1030
rect 4099 856 4145 902
rect 4323 1238 4369 1284
rect 4435 1238 4481 1284
rect 4323 1111 4369 1157
rect 4435 1118 4481 1164
rect 4659 1238 4705 1284
rect 4767 1238 4813 1284
rect 4659 1118 4705 1164
rect 4767 1110 4813 1156
rect 4323 984 4369 1030
rect 4323 856 4369 902
rect 4767 983 4813 1029
rect 4767 856 4813 902
rect 4991 1238 5037 1284
rect 4991 1110 5037 1156
rect 4991 983 5037 1029
rect 4991 856 5037 902
rect 5232 1224 5278 1270
rect 5232 1102 5278 1148
rect 5232 979 5278 1025
rect 5232 856 5278 902
rect 5456 1224 5502 1270
rect 5456 1102 5502 1148
rect 5456 979 5502 1025
rect 5456 856 5502 902
rect 5680 1224 5726 1270
rect 5680 1102 5726 1148
rect 5680 979 5726 1025
rect 5680 856 5726 902
rect 5904 1224 5950 1270
rect 5904 1102 5950 1148
rect 5904 979 5950 1025
rect 5904 856 5950 902
rect 6128 1224 6174 1270
rect 6128 1102 6174 1148
rect 6128 979 6174 1025
rect 6128 856 6174 902
rect 6352 1224 6398 1270
rect 6352 1102 6398 1148
rect 6352 979 6398 1025
rect 6352 856 6398 902
rect 6576 1224 6622 1270
rect 6576 1102 6622 1148
rect 6576 979 6622 1025
rect 6576 856 6622 902
rect 6800 1224 6846 1270
rect 6800 1102 6846 1148
rect 6800 979 6846 1025
rect 6800 856 6846 902
<< psubdiff >>
rect 1244 3525 1610 3544
rect 1244 3291 1263 3525
rect 1591 3291 1610 3525
rect 1244 3272 1610 3291
rect 4372 3525 4456 3544
rect 4372 3291 4391 3525
rect 4437 3291 4456 3525
rect 4372 3272 4456 3291
rect 7032 3525 7210 3544
rect 7032 3291 7051 3525
rect 7191 3291 7210 3525
rect 7032 3272 7210 3291
rect 7032 490 7210 509
rect 7032 256 7051 490
rect 7191 256 7210 490
rect 7032 237 7210 256
<< nsubdiff >>
rect 1706 2249 1790 2268
rect 1706 2015 1725 2249
rect 1771 2015 1790 2249
rect 1706 1996 1790 2015
rect 4372 2249 4456 2268
rect 4372 2015 4391 2249
rect 4437 2015 4456 2249
rect 4372 1996 4456 2015
rect 7032 2249 7210 2268
rect 7032 2015 7051 2249
rect 7191 2015 7210 2249
rect 7032 1996 7210 2015
rect 79 1186 233 1243
rect 79 1140 133 1186
rect 179 1140 233 1186
rect 79 1022 233 1140
rect 79 976 133 1022
rect 179 976 233 1022
rect 79 920 233 976
rect 7047 1186 7201 1243
rect 7047 1140 7101 1186
rect 7147 1140 7201 1186
rect 7047 1022 7201 1140
rect 7047 976 7101 1022
rect 7147 976 7201 1022
rect 7047 920 7201 976
<< psubdiffcont >>
rect 1263 3291 1591 3525
rect 4391 3291 4437 3525
rect 7051 3291 7191 3525
rect 7051 256 7191 490
<< nsubdiffcont >>
rect 1725 2015 1771 2249
rect 4391 2015 4437 2249
rect 7051 2015 7191 2249
rect 133 1140 179 1186
rect 133 976 179 1022
rect 7101 1140 7147 1186
rect 7101 976 7147 1022
<< polysilicon >>
rect 252 3614 372 3658
rect 476 3614 596 3658
rect 700 3614 820 3658
rect 2023 3598 2143 3642
rect 2247 3598 2367 3642
rect 2471 3598 2591 3642
rect 2695 3598 2815 3642
rect 2919 3598 3039 3642
rect 3143 3598 3263 3642
rect 3367 3598 3487 3642
rect 3591 3598 3711 3642
rect 3815 3598 3935 3642
rect 4039 3598 4159 3642
rect 4669 3598 4789 3642
rect 4893 3598 5013 3642
rect 5117 3598 5237 3642
rect 5341 3598 5461 3642
rect 5565 3598 5685 3642
rect 5789 3598 5909 3642
rect 6013 3598 6133 3642
rect 6237 3598 6357 3642
rect 6461 3598 6581 3642
rect 6685 3598 6805 3642
rect 252 2380 372 3214
rect 476 2380 596 3214
rect 700 2380 820 3214
rect 2023 3004 2143 3214
rect 2247 3004 2367 3214
rect 2471 3004 2591 3214
rect 2695 3004 2815 3214
rect 2919 3004 3039 3214
rect 3143 3004 3263 3214
rect 3367 3004 3487 3214
rect 3591 3004 3711 3214
rect 3815 3004 3935 3214
rect 4039 3004 4159 3214
rect 1607 2920 4159 3004
rect 1607 2870 1785 2920
rect 1607 2824 1626 2870
rect 1766 2824 1785 2870
rect 2023 2828 2143 2920
rect 2247 2828 2367 2920
rect 2471 2828 2591 2920
rect 2695 2828 2815 2920
rect 2919 2828 3039 2920
rect 3143 2828 3263 2920
rect 3367 2828 3487 2920
rect 3591 2828 3711 2920
rect 3815 2828 3935 2920
rect 4039 2828 4159 2920
rect 4669 2828 4789 3214
rect 4893 2828 5013 3214
rect 5117 2828 5237 3214
rect 5341 2828 5461 3214
rect 5565 2828 5685 3214
rect 5789 2828 5909 3214
rect 6013 2828 6133 3214
rect 6237 2828 6357 3214
rect 6461 2828 6581 3214
rect 6685 2828 6805 3214
rect 1607 2805 1785 2824
rect 924 2380 1044 2490
rect 1148 2380 1268 2490
rect 1372 2380 1492 2490
rect 252 1705 372 1884
rect 476 1705 596 1884
rect 700 1705 820 1884
rect 924 1705 1044 1884
rect 1148 1705 1268 1884
rect 1372 1705 1492 1884
rect 2023 1840 2143 1884
rect 2247 1840 2367 1884
rect 2471 1840 2591 1884
rect 2695 1840 2815 1884
rect 2919 1840 3039 1884
rect 3143 1840 3263 1884
rect 3367 1840 3487 1884
rect 3591 1840 3711 1884
rect 3815 1840 3935 1884
rect 4039 1840 4159 1884
rect 252 1686 1492 1705
rect 252 1640 470 1686
rect 610 1640 1492 1686
rect 252 1621 1492 1640
rect 4669 1698 4789 1884
rect 4893 1698 5013 1884
rect 5117 1698 5237 1884
rect 5341 1698 5461 1884
rect 5565 1698 5685 1884
rect 5789 1698 5909 1884
rect 6013 1698 6133 1884
rect 6237 1698 6357 1884
rect 6461 1698 6581 1884
rect 6685 1698 6805 1884
rect 4669 1679 6805 1698
rect 4669 1633 5407 1679
rect 5547 1633 5849 1679
rect 5989 1633 6303 1679
rect 6443 1633 6646 1679
rect 6786 1633 6805 1679
rect 4669 1614 6805 1633
rect 1181 1459 2156 1520
rect 451 1429 629 1448
rect 451 1383 470 1429
rect 610 1383 629 1429
rect 451 1364 629 1383
rect 509 1297 629 1364
rect 733 1297 853 1370
rect 1181 1297 1301 1459
rect 1688 1297 1808 1370
rect 2036 1035 2156 1459
rect 4510 1480 4767 1499
rect 3293 1411 3413 1455
rect 3517 1411 3637 1455
rect 3950 1430 4426 1449
rect 2374 1341 2493 1370
rect 2374 1297 2494 1341
rect 2822 1297 2942 1341
rect 3950 1384 4267 1430
rect 4407 1384 4426 1430
rect 3950 1365 4426 1384
rect 4510 1434 4608 1480
rect 4748 1434 4767 1480
rect 4510 1415 4767 1434
rect 3950 1297 4070 1365
rect 4174 1297 4294 1365
rect 4510 1297 4630 1415
rect 4842 1297 4962 1614
rect 5307 1327 5426 1370
rect 5531 1327 5650 1370
rect 5755 1327 5874 1370
rect 5979 1327 6098 1370
rect 6203 1327 6322 1370
rect 6427 1327 6546 1370
rect 6651 1327 6770 1370
rect 4510 1061 4630 1105
rect 5307 1283 5427 1327
rect 5531 1283 5651 1327
rect 5755 1283 5875 1327
rect 5979 1283 6099 1327
rect 6203 1283 6323 1327
rect 6427 1283 6547 1327
rect 6651 1283 6771 1327
rect 509 405 629 843
rect 733 405 853 843
rect 1181 677 1301 843
rect 1688 783 1808 843
rect 2036 799 2156 843
rect 1011 658 1301 677
rect 1011 612 1030 658
rect 1170 612 1301 658
rect 1011 593 1301 612
rect 1364 764 1974 783
rect 1364 624 1383 764
rect 1429 722 1974 764
rect 1429 624 1448 722
rect 1883 685 1974 722
rect 2374 753 2494 843
rect 2374 734 2668 753
rect 2374 688 2509 734
rect 2649 688 2668 734
rect 1364 605 1448 624
rect 1181 487 1301 593
rect 1688 563 1808 636
rect 1883 624 2270 685
rect 2150 564 2270 624
rect 2374 669 2668 688
rect 2374 564 2494 669
rect 2822 564 2942 843
rect 3293 564 3413 843
rect 3517 564 3637 843
rect 3950 769 4070 843
rect 4174 769 4294 843
rect 3950 607 4069 636
rect 4174 607 4293 636
rect 509 140 629 213
rect 733 103 853 213
rect 733 84 911 103
rect 733 38 752 84
rect 892 38 911 84
rect 733 19 911 38
rect 1181 32 1301 295
rect 2150 299 2270 372
rect 2374 328 2494 372
rect 2374 299 2493 328
rect 1688 32 1808 109
rect 2822 89 2942 372
rect 3950 563 4070 607
rect 4174 563 4294 607
rect 1181 -73 1808 32
rect 2439 70 2942 89
rect 2439 24 2458 70
rect 2598 24 2942 70
rect 2439 5 2942 24
rect 3293 89 3413 324
rect 3517 89 3637 324
rect 4618 440 4738 484
rect 4842 440 4962 843
rect 5307 751 5427 843
rect 5531 751 5651 843
rect 5755 751 5875 843
rect 5979 751 6099 843
rect 6203 751 6323 843
rect 6427 751 6547 843
rect 6651 751 6771 843
rect 5154 732 6771 751
rect 5154 686 5173 732
rect 5313 686 6771 732
rect 5154 667 6771 686
rect 5307 559 5427 667
rect 5531 559 5651 667
rect 5755 559 5875 667
rect 5979 559 6099 667
rect 6203 559 6323 667
rect 6427 559 6547 667
rect 6651 559 6771 667
rect 5307 337 5427 381
rect 5531 337 5651 381
rect 5755 337 5875 381
rect 5979 337 6099 381
rect 6203 337 6323 381
rect 6427 337 6547 381
rect 6651 337 6771 381
rect 5307 308 5426 337
rect 5531 308 5650 337
rect 5755 308 5874 337
rect 5979 308 6098 337
rect 6203 308 6322 337
rect 3293 70 3637 89
rect 3293 24 3312 70
rect 3452 24 3637 70
rect 3293 5 3637 24
rect 3950 8 4070 109
rect 4174 8 4294 109
rect 4618 83 4738 248
rect 4842 204 4962 248
rect 1688 -182 1808 -73
rect 3950 -18 4294 8
rect 4560 64 4738 83
rect 4560 18 4579 64
rect 4719 18 4738 64
rect 4560 -1 4738 18
rect 3950 -64 3969 -18
rect 4109 -58 4294 -18
rect 4109 -64 4128 -58
rect 3950 -83 4128 -64
rect 1688 -201 1866 -182
rect 1688 -247 1707 -201
rect 1847 -247 1866 -201
rect 1688 -266 1866 -247
<< polycontact >>
rect 1626 2824 1766 2870
rect 470 1640 610 1686
rect 5407 1633 5547 1679
rect 5849 1633 5989 1679
rect 6303 1633 6443 1679
rect 6646 1633 6786 1679
rect 470 1383 610 1429
rect 4267 1384 4407 1430
rect 4608 1434 4748 1480
rect 1030 612 1170 658
rect 1383 624 1429 764
rect 2509 688 2649 734
rect 752 38 892 84
rect 2458 24 2598 70
rect 5173 686 5313 732
rect 3312 24 3452 70
rect 4579 18 4719 64
rect 3969 -64 4109 -18
rect 1707 -247 1847 -201
<< metal1 >>
rect 177 3601 223 3614
rect 401 3601 447 3614
rect 625 3601 671 3614
rect 849 3601 895 3614
rect 1948 3585 1994 3598
rect 162 3543 238 3555
rect 162 3283 174 3543
rect 226 3283 238 3543
rect 162 3273 238 3283
rect 162 3271 177 3273
rect 223 3271 238 3273
rect 401 3492 447 3555
rect 401 3383 447 3446
rect 401 3273 447 3337
rect 177 3214 223 3227
rect 610 3543 686 3555
rect 610 3283 622 3543
rect 674 3283 686 3543
rect 610 3273 686 3283
rect 610 3271 625 3273
rect 401 2881 447 3227
rect 671 3271 686 3273
rect 849 3492 895 3555
rect 1291 3543 1575 3555
rect 1291 3536 1303 3543
rect 849 3383 895 3446
rect 849 3273 895 3337
rect 1252 3525 1303 3536
rect 1563 3536 1575 3543
rect 1933 3543 1948 3555
rect 2172 3585 2218 3598
rect 1994 3543 2009 3555
rect 1563 3525 1602 3536
rect 1252 3291 1263 3525
rect 1591 3291 1602 3525
rect 1252 3283 1303 3291
rect 1563 3283 1602 3291
rect 1252 3280 1602 3283
rect 1933 3283 1945 3543
rect 1997 3283 2009 3543
rect 625 3214 671 3227
rect 1291 3271 1575 3280
rect 1933 3273 2009 3283
rect 1933 3271 1948 3273
rect 849 2881 895 3227
rect 1994 3271 2009 3273
rect 2396 3585 2442 3598
rect 2172 3481 2218 3539
rect 2172 3377 2218 3435
rect 2172 3273 2218 3331
rect 1948 3214 1994 3227
rect 2381 3543 2396 3555
rect 2620 3585 2666 3598
rect 2442 3543 2457 3555
rect 2381 3283 2393 3543
rect 2445 3283 2457 3543
rect 2381 3273 2457 3283
rect 2381 3271 2396 3273
rect 2172 3052 2218 3227
rect 2442 3271 2457 3273
rect 2844 3585 2890 3598
rect 2620 3481 2666 3539
rect 2620 3377 2666 3435
rect 2620 3273 2666 3331
rect 2396 3214 2442 3227
rect 2829 3543 2844 3555
rect 3068 3585 3114 3598
rect 2890 3543 2905 3555
rect 2829 3283 2841 3543
rect 2893 3283 2905 3543
rect 2829 3273 2905 3283
rect 2829 3271 2844 3273
rect 2004 3040 2392 3052
rect 2004 3037 2016 3040
rect 1397 2991 2016 3037
rect 2004 2988 2016 2991
rect 2380 3037 2392 3040
rect 2620 3037 2666 3227
rect 2890 3271 2905 3273
rect 3292 3585 3338 3598
rect 3068 3481 3114 3539
rect 3068 3377 3114 3435
rect 3068 3273 3114 3331
rect 2844 3214 2890 3227
rect 3277 3543 3292 3555
rect 3516 3585 3562 3598
rect 3338 3543 3353 3555
rect 3277 3283 3289 3543
rect 3341 3283 3353 3543
rect 3277 3273 3353 3283
rect 3277 3271 3292 3273
rect 3068 3037 3114 3227
rect 3338 3271 3353 3273
rect 3740 3585 3786 3598
rect 3516 3481 3562 3539
rect 3516 3377 3562 3435
rect 3516 3273 3562 3331
rect 3292 3214 3338 3227
rect 3725 3543 3740 3555
rect 3964 3585 4010 3598
rect 3786 3543 3801 3555
rect 3725 3283 3737 3543
rect 3789 3283 3801 3543
rect 3725 3273 3801 3283
rect 3725 3271 3740 3273
rect 3516 3037 3562 3227
rect 3786 3271 3801 3273
rect 4188 3585 4234 3598
rect 3964 3481 4010 3539
rect 3964 3377 4010 3435
rect 3964 3273 4010 3331
rect 3740 3214 3786 3227
rect 4173 3543 4188 3555
rect 4594 3585 4640 3598
rect 4234 3543 4249 3555
rect 4173 3283 4185 3543
rect 4237 3283 4249 3543
rect 4173 3273 4249 3283
rect 4173 3271 4188 3273
rect 3964 3037 4010 3227
rect 4234 3271 4249 3273
rect 4376 3543 4452 3555
rect 4376 3283 4388 3543
rect 4440 3283 4452 3543
rect 4376 3271 4452 3283
rect 4579 3543 4594 3555
rect 4818 3585 4864 3598
rect 4640 3543 4655 3555
rect 4579 3283 4591 3543
rect 4643 3283 4655 3543
rect 4579 3273 4655 3283
rect 4579 3271 4594 3273
rect 4188 3214 4234 3227
rect 4640 3271 4655 3273
rect 5042 3585 5088 3598
rect 4818 3481 4864 3539
rect 4818 3377 4864 3435
rect 4818 3273 4864 3331
rect 4594 3214 4640 3227
rect 5027 3543 5042 3555
rect 5266 3585 5312 3598
rect 5088 3543 5103 3555
rect 5027 3283 5039 3543
rect 5091 3283 5103 3543
rect 5027 3273 5103 3283
rect 5027 3271 5042 3273
rect 2380 2991 4010 3037
rect 2380 2988 2392 2991
rect 2004 2976 2392 2988
rect 401 2870 1777 2881
rect 401 2824 1626 2870
rect 1766 2824 1777 2870
rect 401 2813 1777 2824
rect 1948 2815 1994 2828
rect 177 2367 223 2380
rect 177 2279 223 2321
rect 401 2367 447 2813
rect 162 2267 238 2279
rect 162 2007 174 2267
rect 226 2007 238 2267
rect 162 2003 177 2007
rect 223 2003 238 2007
rect 162 1995 238 2003
rect 401 2261 447 2321
rect 625 2367 671 2380
rect 625 2279 671 2321
rect 849 2367 895 2813
rect 401 2155 447 2215
rect 401 2049 447 2109
rect 177 1943 223 1995
rect 177 1884 223 1897
rect 401 1943 447 2003
rect 610 2267 686 2279
rect 610 2007 622 2267
rect 674 2007 686 2267
rect 610 2003 625 2007
rect 671 2003 686 2007
rect 610 1995 686 2003
rect 849 2261 895 2321
rect 1073 2367 1119 2380
rect 1073 2279 1119 2321
rect 1297 2367 1343 2813
rect 1948 2706 1994 2769
rect 1948 2597 1994 2660
rect 1948 2488 1994 2551
rect 849 2155 895 2215
rect 849 2049 895 2109
rect 401 1884 447 1897
rect 625 1943 671 1995
rect 625 1884 671 1897
rect 849 1943 895 2003
rect 1058 2267 1134 2279
rect 1058 2007 1070 2267
rect 1122 2007 1134 2267
rect 1058 2003 1073 2007
rect 1119 2003 1134 2007
rect 1058 1995 1134 2003
rect 1297 2261 1343 2321
rect 1521 2367 1567 2380
rect 1521 2279 1567 2321
rect 1948 2379 1994 2442
rect 1948 2279 1994 2333
rect 2172 2815 2218 2976
rect 2172 2706 2218 2769
rect 2172 2597 2218 2660
rect 2172 2488 2218 2551
rect 2172 2379 2218 2442
rect 1297 2155 1343 2215
rect 1297 2049 1343 2109
rect 849 1884 895 1897
rect 1073 1943 1119 1995
rect 1073 1884 1119 1897
rect 1297 1943 1343 2003
rect 1506 2267 1582 2279
rect 1506 2007 1518 2267
rect 1570 2007 1582 2267
rect 1506 2003 1521 2007
rect 1567 2003 1582 2007
rect 1506 1995 1582 2003
rect 1710 2267 1786 2279
rect 1710 2007 1722 2267
rect 1774 2007 1786 2267
rect 1710 1995 1786 2007
rect 1933 2270 2009 2279
rect 1933 2267 1948 2270
rect 1994 2267 2009 2270
rect 1933 2007 1945 2267
rect 1997 2007 2009 2267
rect 1933 2006 1948 2007
rect 1994 2006 2009 2007
rect 1933 1995 2009 2006
rect 2172 2270 2218 2333
rect 2396 2815 2442 2828
rect 2396 2706 2442 2769
rect 2396 2597 2442 2660
rect 2396 2488 2442 2551
rect 2396 2379 2442 2442
rect 2396 2279 2442 2333
rect 2620 2815 2666 2991
rect 2620 2706 2666 2769
rect 2620 2597 2666 2660
rect 2620 2488 2666 2551
rect 2620 2379 2666 2442
rect 2172 2161 2218 2224
rect 2172 2052 2218 2115
rect 1297 1884 1343 1897
rect 1521 1943 1567 1995
rect 1521 1884 1567 1897
rect 1948 1943 1994 1995
rect 1948 1884 1994 1897
rect 2172 1943 2218 2006
rect 2381 2270 2457 2279
rect 2381 2267 2396 2270
rect 2442 2267 2457 2270
rect 2381 2007 2393 2267
rect 2445 2007 2457 2267
rect 2381 2006 2396 2007
rect 2442 2006 2457 2007
rect 2381 1995 2457 2006
rect 2620 2270 2666 2333
rect 2844 2815 2890 2828
rect 2844 2706 2890 2769
rect 2844 2597 2890 2660
rect 2844 2488 2890 2551
rect 2844 2379 2890 2442
rect 2844 2279 2890 2333
rect 3068 2815 3114 2991
rect 3068 2706 3114 2769
rect 3068 2597 3114 2660
rect 3068 2488 3114 2551
rect 3068 2379 3114 2442
rect 2620 2161 2666 2224
rect 2620 2052 2666 2115
rect 2172 1884 2218 1897
rect 2396 1943 2442 1995
rect 2396 1884 2442 1897
rect 2620 1943 2666 2006
rect 2829 2270 2905 2279
rect 2829 2267 2844 2270
rect 2890 2267 2905 2270
rect 2829 2007 2841 2267
rect 2893 2007 2905 2267
rect 2829 2006 2844 2007
rect 2890 2006 2905 2007
rect 2829 1995 2905 2006
rect 3068 2270 3114 2333
rect 3292 2815 3338 2828
rect 3292 2706 3338 2769
rect 3292 2597 3338 2660
rect 3292 2488 3338 2551
rect 3292 2379 3338 2442
rect 3292 2279 3338 2333
rect 3516 2815 3562 2991
rect 3516 2706 3562 2769
rect 3516 2597 3562 2660
rect 3516 2488 3562 2551
rect 3516 2379 3562 2442
rect 3068 2161 3114 2224
rect 3068 2052 3114 2115
rect 2620 1884 2666 1897
rect 2844 1943 2890 1995
rect 2844 1884 2890 1897
rect 3068 1943 3114 2006
rect 3277 2270 3353 2279
rect 3277 2267 3292 2270
rect 3338 2267 3353 2270
rect 3277 2007 3289 2267
rect 3341 2007 3353 2267
rect 3277 2006 3292 2007
rect 3338 2006 3353 2007
rect 3277 1995 3353 2006
rect 3516 2270 3562 2333
rect 3740 2815 3786 2828
rect 3740 2706 3786 2769
rect 3740 2597 3786 2660
rect 3740 2488 3786 2551
rect 3740 2379 3786 2442
rect 3740 2279 3786 2333
rect 3964 2815 4010 2991
rect 4818 3025 4864 3227
rect 5088 3271 5103 3273
rect 5490 3585 5536 3598
rect 5266 3481 5312 3539
rect 5266 3377 5312 3435
rect 5266 3273 5312 3331
rect 5042 3214 5088 3227
rect 5475 3543 5490 3555
rect 5714 3585 5760 3598
rect 5536 3543 5551 3555
rect 5475 3283 5487 3543
rect 5539 3283 5551 3543
rect 5475 3273 5551 3283
rect 5475 3271 5490 3273
rect 5266 3025 5312 3227
rect 5536 3271 5551 3273
rect 5938 3585 5984 3598
rect 5714 3481 5760 3539
rect 5714 3377 5760 3435
rect 5714 3273 5760 3331
rect 5490 3214 5536 3227
rect 5923 3543 5938 3555
rect 6162 3585 6208 3598
rect 5984 3543 5999 3555
rect 5923 3283 5935 3543
rect 5987 3283 5999 3543
rect 5923 3273 5999 3283
rect 5923 3271 5938 3273
rect 5714 3025 5760 3227
rect 5984 3271 5999 3273
rect 6386 3585 6432 3598
rect 6162 3481 6208 3539
rect 6162 3377 6208 3435
rect 6162 3273 6208 3331
rect 5938 3214 5984 3227
rect 6371 3543 6386 3555
rect 6610 3585 6656 3598
rect 6432 3543 6447 3555
rect 6371 3283 6383 3543
rect 6435 3283 6447 3543
rect 6371 3273 6447 3283
rect 6371 3271 6386 3273
rect 6162 3025 6208 3227
rect 6432 3271 6447 3273
rect 6834 3585 6880 3598
rect 6610 3481 6656 3539
rect 6610 3377 6656 3435
rect 6610 3273 6656 3331
rect 6386 3214 6432 3227
rect 6819 3543 6834 3555
rect 6880 3543 6895 3555
rect 6819 3283 6831 3543
rect 6883 3283 6895 3543
rect 6819 3273 6895 3283
rect 6819 3271 6834 3273
rect 6610 3025 6656 3227
rect 6880 3271 6895 3273
rect 7038 3543 7218 3555
rect 7038 3283 7050 3543
rect 7206 3283 7218 3543
rect 7038 3271 7218 3283
rect 6834 3214 6880 3227
rect 4818 2979 6656 3025
rect 3964 2706 4010 2769
rect 3964 2597 4010 2660
rect 3964 2488 4010 2551
rect 3964 2379 4010 2442
rect 3516 2161 3562 2224
rect 3516 2052 3562 2115
rect 3068 1884 3114 1897
rect 3292 1943 3338 1995
rect 3292 1884 3338 1897
rect 3516 1943 3562 2006
rect 3725 2270 3801 2279
rect 3725 2267 3740 2270
rect 3786 2267 3801 2270
rect 3725 2007 3737 2267
rect 3789 2007 3801 2267
rect 3725 2006 3740 2007
rect 3786 2006 3801 2007
rect 3725 1995 3801 2006
rect 3964 2270 4010 2333
rect 4188 2815 4234 2828
rect 4188 2706 4234 2769
rect 4188 2597 4234 2660
rect 4188 2488 4234 2551
rect 4188 2379 4234 2442
rect 4188 2279 4234 2333
rect 4594 2815 4640 2828
rect 4594 2706 4640 2769
rect 4594 2597 4640 2660
rect 4594 2488 4640 2551
rect 4594 2379 4640 2442
rect 4594 2279 4640 2333
rect 4818 2815 4864 2979
rect 4818 2706 4864 2769
rect 4818 2597 4864 2660
rect 4818 2488 4864 2551
rect 4818 2379 4864 2442
rect 3964 2161 4010 2224
rect 3964 2052 4010 2115
rect 3516 1884 3562 1897
rect 3740 1943 3786 1995
rect 3740 1884 3786 1897
rect 3964 1943 4010 2006
rect 4173 2270 4249 2279
rect 4173 2267 4188 2270
rect 4234 2267 4249 2270
rect 4173 2007 4185 2267
rect 4237 2007 4249 2267
rect 4173 2006 4188 2007
rect 4234 2006 4249 2007
rect 4173 1995 4249 2006
rect 4376 2267 4452 2279
rect 4376 2007 4388 2267
rect 4440 2007 4452 2267
rect 4376 1995 4452 2007
rect 4579 2270 4655 2279
rect 4579 2267 4594 2270
rect 4640 2267 4655 2270
rect 4579 2007 4591 2267
rect 4643 2007 4655 2267
rect 4579 2006 4594 2007
rect 4640 2006 4655 2007
rect 4579 1995 4655 2006
rect 4818 2270 4864 2333
rect 5042 2815 5088 2828
rect 5042 2706 5088 2769
rect 5042 2597 5088 2660
rect 5042 2488 5088 2551
rect 5042 2379 5088 2442
rect 5042 2279 5088 2333
rect 5266 2815 5312 2979
rect 5266 2706 5312 2769
rect 5266 2597 5312 2660
rect 5266 2488 5312 2551
rect 5266 2379 5312 2442
rect 4818 2161 4864 2224
rect 4818 2052 4864 2115
rect 3964 1884 4010 1897
rect 4188 1943 4234 1995
rect 4188 1884 4234 1897
rect 4594 1943 4640 1995
rect 4594 1884 4640 1897
rect 4818 1943 4864 2006
rect 5027 2270 5103 2279
rect 5027 2267 5042 2270
rect 5088 2267 5103 2270
rect 5027 2007 5039 2267
rect 5091 2007 5103 2267
rect 5027 2006 5042 2007
rect 5088 2006 5103 2007
rect 5027 1995 5103 2006
rect 5266 2270 5312 2333
rect 5490 2815 5536 2828
rect 5490 2706 5536 2769
rect 5490 2597 5536 2660
rect 5490 2488 5536 2551
rect 5490 2379 5536 2442
rect 5490 2279 5536 2333
rect 5714 2815 5760 2979
rect 5714 2706 5760 2769
rect 5714 2597 5760 2660
rect 5714 2488 5760 2551
rect 5714 2379 5760 2442
rect 5266 2161 5312 2224
rect 5266 2052 5312 2115
rect 4818 1884 4864 1897
rect 5042 1943 5088 1995
rect 5042 1884 5088 1897
rect 5266 1943 5312 2006
rect 5475 2270 5551 2279
rect 5475 2267 5490 2270
rect 5536 2267 5551 2270
rect 5475 2007 5487 2267
rect 5539 2007 5551 2267
rect 5475 2006 5490 2007
rect 5536 2006 5551 2007
rect 5475 1995 5551 2006
rect 5714 2270 5760 2333
rect 5938 2815 5984 2828
rect 5938 2706 5984 2769
rect 5938 2597 5984 2660
rect 5938 2488 5984 2551
rect 5938 2379 5984 2442
rect 5938 2279 5984 2333
rect 6162 2815 6208 2979
rect 6162 2706 6208 2769
rect 6162 2597 6208 2660
rect 6162 2488 6208 2551
rect 6162 2379 6208 2442
rect 5714 2161 5760 2224
rect 5714 2052 5760 2115
rect 5266 1884 5312 1897
rect 5490 1943 5536 1995
rect 5490 1884 5536 1897
rect 5714 1943 5760 2006
rect 5923 2270 5999 2279
rect 5923 2267 5938 2270
rect 5984 2267 5999 2270
rect 5923 2007 5935 2267
rect 5987 2007 5999 2267
rect 5923 2006 5938 2007
rect 5984 2006 5999 2007
rect 5923 1995 5999 2006
rect 6162 2270 6208 2333
rect 6386 2815 6432 2828
rect 6386 2706 6432 2769
rect 6386 2597 6432 2660
rect 6386 2488 6432 2551
rect 6386 2379 6432 2442
rect 6386 2279 6432 2333
rect 6610 2815 6656 2979
rect 6610 2706 6656 2769
rect 6610 2597 6656 2660
rect 6610 2488 6656 2551
rect 6610 2379 6656 2442
rect 6162 2161 6208 2224
rect 6162 2052 6208 2115
rect 5714 1884 5760 1897
rect 5938 1943 5984 1995
rect 5938 1884 5984 1897
rect 6162 1943 6208 2006
rect 6371 2270 6447 2279
rect 6371 2267 6386 2270
rect 6432 2267 6447 2270
rect 6371 2007 6383 2267
rect 6435 2007 6447 2267
rect 6371 2006 6386 2007
rect 6432 2006 6447 2007
rect 6371 1995 6447 2006
rect 6610 2270 6656 2333
rect 6834 2815 6880 2828
rect 6834 2706 6880 2769
rect 6834 2597 6880 2660
rect 6834 2488 6880 2551
rect 6834 2379 6880 2442
rect 6834 2279 6880 2333
rect 6610 2161 6656 2224
rect 6610 2052 6656 2115
rect 6162 1884 6208 1897
rect 6386 1943 6432 1995
rect 6386 1884 6432 1897
rect 6610 1943 6656 2006
rect 6819 2270 6895 2279
rect 6819 2267 6834 2270
rect 6880 2267 6895 2270
rect 6819 2007 6831 2267
rect 6883 2007 6895 2267
rect 6819 2006 6834 2007
rect 6880 2006 6895 2007
rect 6819 1995 6895 2006
rect 7032 2267 7212 2279
rect 7032 2007 7044 2267
rect 7200 2007 7212 2267
rect 7032 1995 7212 2007
rect 6610 1884 6656 1897
rect 6834 1943 6880 1995
rect 6834 1884 6880 1897
rect 459 1686 621 1697
rect 459 1640 470 1686
rect 610 1640 621 1686
rect 459 1429 621 1640
rect 5396 1679 5558 1690
rect 5396 1633 5407 1679
rect 5547 1633 5558 1679
rect 5396 1622 5558 1633
rect 5838 1679 6000 1690
rect 5838 1633 5849 1679
rect 5989 1633 6000 1679
rect 5838 1622 6000 1633
rect 6292 1679 6454 1690
rect 6292 1633 6303 1679
rect 6443 1633 6454 1679
rect 6292 1622 6454 1633
rect 6635 1679 6846 1690
rect 6635 1633 6646 1679
rect 6786 1633 6846 1679
rect 6635 1622 6846 1633
rect 459 1383 470 1429
rect 610 1383 621 1429
rect 459 1372 621 1383
rect 882 1563 4327 1609
rect 434 1284 480 1297
rect 91 1216 221 1257
rect 91 1164 130 1216
rect 182 1164 221 1216
rect 91 1140 133 1164
rect 179 1140 221 1164
rect 91 1022 221 1140
rect 91 998 133 1022
rect 179 998 221 1022
rect 91 946 130 998
rect 182 946 221 998
rect 91 906 221 946
rect 658 1284 704 1297
rect 434 1157 480 1238
rect 434 1030 480 1111
rect 434 902 480 984
rect 616 1238 658 1246
rect 882 1284 928 1563
rect 1262 1487 1442 1499
rect 1262 1435 1274 1487
rect 1430 1435 1442 1487
rect 1262 1423 1442 1435
rect 3442 1457 4145 1512
rect 1329 1416 1376 1423
rect 1106 1289 1152 1297
rect 704 1238 746 1246
rect 616 1205 746 1238
rect 616 1153 655 1205
rect 707 1153 746 1205
rect 616 1111 658 1153
rect 704 1111 746 1153
rect 616 1030 746 1111
rect 616 987 658 1030
rect 704 987 746 1030
rect 616 935 655 987
rect 707 935 746 987
rect 616 902 746 935
rect 616 895 658 902
rect 91 514 221 555
rect 91 462 130 514
rect 182 462 221 514
rect 91 438 133 462
rect 179 438 221 462
rect 91 320 221 438
rect 91 296 133 320
rect 179 296 221 320
rect 91 244 130 296
rect 182 244 221 296
rect 91 204 221 244
rect 434 392 480 856
rect 704 895 746 902
rect 882 1157 928 1238
rect 882 1030 928 1111
rect 882 902 928 984
rect 658 843 704 856
rect 882 669 928 856
rect 1064 1284 1193 1289
rect 1064 1238 1106 1284
rect 1152 1246 1193 1284
rect 1330 1284 1376 1416
rect 3218 1398 3264 1411
rect 1613 1289 1659 1297
rect 1837 1289 1883 1297
rect 1152 1238 1194 1246
rect 1064 1205 1194 1238
rect 1064 1153 1103 1205
rect 1155 1153 1194 1205
rect 1064 1111 1106 1153
rect 1152 1111 1194 1153
rect 1064 1030 1194 1111
rect 1064 987 1106 1030
rect 1152 987 1194 1030
rect 1064 935 1103 987
rect 1155 935 1194 987
rect 1064 902 1194 935
rect 1064 856 1106 902
rect 1152 895 1194 902
rect 1330 1157 1376 1238
rect 1330 1030 1376 1111
rect 1330 902 1376 984
rect 1152 856 1193 895
rect 1064 852 1193 856
rect 1106 843 1152 852
rect 1330 775 1376 856
rect 1572 1284 1700 1289
rect 1572 1238 1613 1284
rect 1659 1238 1700 1284
rect 1572 1164 1700 1238
rect 1572 1112 1610 1164
rect 1662 1112 1700 1164
rect 1572 1111 1613 1112
rect 1659 1111 1700 1112
rect 1572 1030 1700 1111
rect 1572 984 1613 1030
rect 1659 984 1700 1030
rect 1572 947 1700 984
rect 1572 895 1610 947
rect 1662 895 1700 947
rect 1572 856 1613 895
rect 1659 856 1700 895
rect 1330 764 1440 775
rect 882 658 1181 669
rect 882 612 1030 658
rect 1170 612 1181 658
rect 882 601 1181 612
rect 1330 624 1383 764
rect 1429 624 1440 764
rect 1330 613 1440 624
rect 1572 729 1700 856
rect 1572 677 1610 729
rect 1662 677 1700 729
rect 434 272 480 346
rect 434 -85 480 226
rect 616 514 746 555
rect 616 462 655 514
rect 707 462 746 514
rect 616 392 746 462
rect 616 346 658 392
rect 704 346 746 392
rect 616 296 746 346
rect 616 244 655 296
rect 707 244 746 296
rect 616 226 658 244
rect 704 226 746 244
rect 616 204 746 226
rect 882 392 928 601
rect 882 272 928 346
rect 1065 513 1193 554
rect 1065 461 1103 513
rect 1155 461 1193 513
rect 1065 428 1106 461
rect 1152 428 1193 461
rect 1065 354 1193 428
rect 1065 327 1106 354
rect 1152 327 1193 354
rect 1065 275 1103 327
rect 1155 275 1193 327
rect 1065 235 1193 275
rect 1330 474 1376 613
rect 1330 354 1376 428
rect 882 213 928 226
rect 632 84 972 95
rect 632 55 752 84
rect 892 55 972 84
rect 632 3 670 55
rect 722 38 752 55
rect 722 3 882 38
rect 934 3 972 55
rect 632 -38 972 3
rect 1330 -76 1376 308
rect 1572 550 1700 677
rect 1572 511 1613 550
rect 1659 511 1700 550
rect 1572 459 1610 511
rect 1662 459 1700 511
rect 1572 423 1700 459
rect 1572 377 1613 423
rect 1659 377 1700 423
rect 1572 296 1700 377
rect 1572 294 1613 296
rect 1659 294 1700 296
rect 1572 242 1610 294
rect 1662 242 1700 294
rect 1572 201 1700 242
rect 1796 1284 1924 1289
rect 1796 1238 1837 1284
rect 1883 1238 1924 1284
rect 1796 1157 1924 1238
rect 1796 1111 1837 1157
rect 1883 1111 1924 1157
rect 1796 1035 1924 1111
rect 2299 1284 2345 1297
rect 2523 1289 2569 1297
rect 2747 1289 2793 1297
rect 2971 1289 3017 1297
rect 2481 1284 2609 1289
rect 2481 1246 2523 1284
rect 2299 1157 2345 1238
rect 2299 1036 2345 1111
rect 2190 1035 2345 1036
rect 1796 1030 2007 1035
rect 1796 984 1837 1030
rect 1883 1022 2007 1030
rect 1883 984 1961 1022
rect 1796 976 1961 984
rect 1796 902 2007 976
rect 1796 856 1837 902
rect 1883 856 1961 902
rect 1796 843 2007 856
rect 2185 1030 2345 1035
rect 2185 1022 2299 1030
rect 2231 984 2299 1022
rect 2231 976 2345 984
rect 2185 902 2345 976
rect 2231 856 2299 902
rect 2480 1238 2523 1246
rect 2569 1246 2609 1284
rect 2734 1284 2806 1289
rect 2569 1238 2610 1246
rect 2480 1205 2610 1238
rect 2480 1153 2519 1205
rect 2571 1153 2610 1205
rect 2480 1111 2523 1153
rect 2569 1111 2610 1153
rect 2480 1030 2610 1111
rect 2480 987 2523 1030
rect 2569 987 2610 1030
rect 2480 935 2519 987
rect 2571 935 2610 987
rect 2480 902 2610 935
rect 2480 895 2523 902
rect 2185 843 2345 856
rect 2481 856 2523 895
rect 2569 895 2610 902
rect 2734 1238 2747 1284
rect 2793 1238 2806 1284
rect 2929 1284 3057 1289
rect 2929 1246 2971 1284
rect 2734 1157 2806 1238
rect 2734 1111 2747 1157
rect 2793 1111 2806 1157
rect 2734 1030 2806 1111
rect 2734 984 2747 1030
rect 2793 984 2806 1030
rect 2734 902 2806 984
rect 2569 856 2609 895
rect 2481 852 2609 856
rect 2734 856 2747 902
rect 2793 856 2806 902
rect 2928 1238 2971 1246
rect 3017 1246 3057 1284
rect 3218 1274 3264 1352
rect 3017 1238 3058 1246
rect 2928 1205 3058 1238
rect 2928 1153 2967 1205
rect 3019 1153 3058 1205
rect 2928 1111 2971 1153
rect 3017 1111 3058 1153
rect 2928 1030 3058 1111
rect 2928 987 2971 1030
rect 3017 987 3058 1030
rect 2928 935 2967 987
rect 3019 935 3058 987
rect 3203 1228 3218 1231
rect 3442 1398 3488 1457
rect 3442 1274 3488 1352
rect 3264 1228 3279 1231
rect 3203 1219 3279 1228
rect 3203 959 3215 1219
rect 3267 959 3279 1219
rect 3203 947 3279 959
rect 3666 1398 3712 1411
rect 3666 1274 3712 1352
rect 3875 1289 3921 1297
rect 3442 1150 3488 1228
rect 3442 1026 3488 1104
rect 2928 902 3058 935
rect 2928 895 2971 902
rect 2523 843 2569 852
rect 1796 554 1924 843
rect 2075 554 2121 564
rect 1796 551 2155 554
rect 1796 550 2075 551
rect 1796 504 1837 550
rect 1883 505 2075 550
rect 2121 505 2155 551
rect 1883 504 2155 505
rect 1796 431 2155 504
rect 1796 423 2075 431
rect 1796 377 1837 423
rect 1883 385 2075 423
rect 2121 385 2155 431
rect 1883 380 2155 385
rect 2299 551 2345 843
rect 2734 745 2806 856
rect 2929 856 2971 895
rect 3017 895 3058 902
rect 3218 902 3264 947
rect 3017 856 3057 895
rect 2929 852 3057 856
rect 2971 843 3017 852
rect 3218 843 3264 856
rect 3442 902 3488 980
rect 3651 1228 3666 1231
rect 3833 1284 3961 1289
rect 3833 1238 3875 1284
rect 3921 1238 3961 1284
rect 4099 1284 4145 1457
rect 4281 1441 4327 1563
rect 4590 1487 4770 1499
rect 4256 1430 4418 1441
rect 4256 1384 4267 1430
rect 4407 1384 4418 1430
rect 4590 1435 4602 1487
rect 4758 1435 4770 1487
rect 4590 1434 4608 1435
rect 4748 1434 4770 1435
rect 4590 1423 4770 1434
rect 4256 1373 4418 1384
rect 3712 1228 3727 1231
rect 3651 1219 3727 1228
rect 3651 959 3663 1219
rect 3715 959 3727 1219
rect 3651 947 3727 959
rect 3833 1157 3961 1238
rect 3833 1111 3875 1157
rect 3921 1111 3961 1157
rect 3833 1030 3961 1111
rect 3833 984 3875 1030
rect 3921 984 3961 1030
rect 2498 734 2806 745
rect 2498 688 2509 734
rect 2649 688 2806 734
rect 2498 677 2806 688
rect 2523 554 2569 564
rect 2299 431 2345 505
rect 1883 377 1924 380
rect 1796 296 1924 377
rect 2075 372 2121 380
rect 2299 372 2345 385
rect 2481 551 2609 554
rect 2481 513 2523 551
rect 2569 513 2609 551
rect 2481 461 2519 513
rect 2571 461 2609 513
rect 2481 431 2609 461
rect 2481 385 2523 431
rect 2569 385 2609 431
rect 1796 250 1837 296
rect 1883 250 1924 296
rect 1613 168 1659 201
rect 1613 109 1659 122
rect 1796 168 1924 250
rect 2481 327 2609 385
rect 2481 275 2519 327
rect 2571 275 2609 327
rect 2481 235 2609 275
rect 2734 551 2806 677
rect 2971 554 3017 564
rect 2734 505 2747 551
rect 2793 505 2806 551
rect 2734 431 2806 505
rect 2734 385 2747 431
rect 2793 385 2806 431
rect 1796 122 1837 168
rect 1883 122 1924 168
rect 1796 81 1924 122
rect 2734 81 2806 385
rect 2929 551 3057 554
rect 2929 513 2971 551
rect 3017 513 3057 551
rect 2929 461 2967 513
rect 3019 461 3057 513
rect 3218 551 3264 564
rect 3218 502 3264 505
rect 3442 551 3488 856
rect 3666 902 3712 947
rect 3666 843 3712 856
rect 3833 902 3961 984
rect 3833 856 3875 902
rect 3921 856 3961 902
rect 4056 1238 4099 1246
rect 4323 1284 4481 1297
rect 4145 1238 4186 1246
rect 4056 1205 4186 1238
rect 4056 1153 4095 1205
rect 4147 1153 4186 1205
rect 4056 1111 4099 1153
rect 4145 1111 4186 1153
rect 4056 1030 4186 1111
rect 4056 987 4099 1030
rect 4145 987 4186 1030
rect 4056 935 4095 987
rect 4147 935 4186 987
rect 4056 902 4186 935
rect 4056 895 4099 902
rect 3833 763 3961 856
rect 4145 895 4186 902
rect 4369 1238 4435 1284
rect 4323 1164 4481 1238
rect 4323 1157 4435 1164
rect 4369 1118 4435 1157
rect 4369 1111 4481 1118
rect 4323 1105 4481 1111
rect 4659 1284 4855 1298
rect 4991 1289 5037 1297
rect 4705 1238 4767 1284
rect 4813 1238 4855 1284
rect 4950 1284 5078 1289
rect 4950 1246 4991 1284
rect 4659 1205 4855 1238
rect 4659 1164 4764 1205
rect 4705 1153 4764 1164
rect 4816 1153 4855 1205
rect 4705 1118 4767 1153
rect 4659 1110 4767 1118
rect 4813 1110 4855 1153
rect 4659 1105 4855 1110
rect 4323 1030 4409 1105
rect 4369 984 4409 1030
rect 4323 902 4409 984
rect 4099 843 4145 856
rect 4369 856 4409 902
rect 4725 1029 4855 1105
rect 4725 987 4767 1029
rect 4813 987 4855 1029
rect 4725 935 4764 987
rect 4816 935 4855 987
rect 4725 902 4855 935
rect 4725 895 4767 902
rect 4323 763 4409 856
rect 4813 895 4855 902
rect 4949 1238 4991 1246
rect 5037 1246 5078 1284
rect 5191 1270 5319 1289
rect 5191 1254 5232 1270
rect 5037 1238 5079 1246
rect 4949 1205 5079 1238
rect 4949 1153 4988 1205
rect 5040 1153 5079 1205
rect 4949 1110 4991 1153
rect 5037 1110 5079 1153
rect 4949 1029 5079 1110
rect 4949 987 4991 1029
rect 5037 987 5079 1029
rect 4949 935 4988 987
rect 5040 935 5079 987
rect 4949 902 5079 935
rect 5190 1224 5232 1254
rect 5278 1254 5319 1270
rect 5418 1270 5534 1622
rect 5278 1224 5320 1254
rect 5190 1214 5320 1224
rect 5190 1162 5229 1214
rect 5281 1162 5320 1214
rect 5190 1148 5320 1162
rect 5190 1102 5232 1148
rect 5278 1102 5320 1148
rect 5190 1025 5320 1102
rect 5190 996 5232 1025
rect 5278 996 5320 1025
rect 5190 944 5229 996
rect 5281 944 5320 996
rect 5190 903 5320 944
rect 5418 1224 5456 1270
rect 5502 1224 5534 1270
rect 5418 1148 5534 1224
rect 5418 1102 5456 1148
rect 5502 1102 5534 1148
rect 5418 1025 5534 1102
rect 5418 979 5456 1025
rect 5502 979 5534 1025
rect 4949 895 4991 902
rect 4767 843 4813 856
rect 4950 856 4991 895
rect 5037 895 5079 902
rect 5191 902 5319 903
rect 5037 856 5078 895
rect 4950 852 5078 856
rect 5191 856 5232 902
rect 5278 856 5319 902
rect 5191 852 5319 856
rect 5418 902 5534 979
rect 5418 856 5456 902
rect 5502 856 5534 902
rect 4991 843 5037 852
rect 5232 843 5278 852
rect 3833 743 4409 763
rect 5418 763 5534 856
rect 5638 1270 5767 1289
rect 5638 1224 5680 1270
rect 5726 1254 5767 1270
rect 5866 1270 5981 1622
rect 5726 1224 5768 1254
rect 5638 1214 5768 1224
rect 5638 1162 5677 1214
rect 5729 1162 5768 1214
rect 5638 1148 5768 1162
rect 5638 1102 5680 1148
rect 5726 1102 5768 1148
rect 5638 1025 5768 1102
rect 5638 996 5680 1025
rect 5726 996 5768 1025
rect 5638 944 5677 996
rect 5729 944 5768 996
rect 5638 903 5768 944
rect 5866 1224 5904 1270
rect 5950 1224 5981 1270
rect 5866 1148 5981 1224
rect 5866 1102 5904 1148
rect 5950 1102 5981 1148
rect 5866 1025 5981 1102
rect 5866 979 5904 1025
rect 5950 979 5981 1025
rect 5638 902 5767 903
rect 5638 856 5680 902
rect 5726 856 5767 902
rect 5638 852 5767 856
rect 5866 902 5981 979
rect 5866 856 5904 902
rect 5950 856 5981 902
rect 5680 843 5726 852
rect 5866 763 5981 856
rect 6086 1270 6215 1289
rect 6086 1224 6128 1270
rect 6174 1254 6215 1270
rect 6314 1270 6429 1622
rect 6174 1224 6216 1254
rect 6086 1214 6216 1224
rect 6086 1162 6125 1214
rect 6177 1162 6216 1214
rect 6086 1148 6216 1162
rect 6086 1102 6128 1148
rect 6174 1102 6216 1148
rect 6086 1025 6216 1102
rect 6086 996 6128 1025
rect 6174 996 6216 1025
rect 6086 944 6125 996
rect 6177 944 6216 996
rect 6086 903 6216 944
rect 6314 1224 6352 1270
rect 6398 1224 6429 1270
rect 6314 1148 6429 1224
rect 6314 1102 6352 1148
rect 6398 1102 6429 1148
rect 6314 1025 6429 1102
rect 6314 979 6352 1025
rect 6398 979 6429 1025
rect 6086 902 6215 903
rect 6086 856 6128 902
rect 6174 856 6215 902
rect 6086 852 6215 856
rect 6314 902 6429 979
rect 6314 856 6352 902
rect 6398 856 6429 902
rect 6128 843 6174 852
rect 6314 763 6429 856
rect 6534 1270 6663 1289
rect 6534 1224 6576 1270
rect 6622 1254 6663 1270
rect 6762 1270 6846 1622
rect 6622 1224 6664 1254
rect 6534 1214 6664 1224
rect 6534 1162 6573 1214
rect 6625 1162 6664 1214
rect 6534 1148 6664 1162
rect 6534 1102 6576 1148
rect 6622 1102 6664 1148
rect 6534 1025 6664 1102
rect 6534 996 6576 1025
rect 6622 996 6664 1025
rect 6534 944 6573 996
rect 6625 944 6664 996
rect 6534 903 6664 944
rect 6762 1224 6800 1270
rect 6762 1148 6846 1224
rect 6762 1102 6800 1148
rect 6762 1025 6846 1102
rect 6762 979 6800 1025
rect 6534 902 6663 903
rect 6534 856 6576 902
rect 6622 856 6663 902
rect 6534 852 6663 856
rect 6762 902 6846 979
rect 7059 1216 7189 1257
rect 7059 1164 7098 1216
rect 7150 1164 7189 1216
rect 7059 1140 7101 1164
rect 7147 1140 7189 1164
rect 7059 1022 7189 1140
rect 7059 998 7101 1022
rect 7147 998 7189 1022
rect 7059 946 7098 998
rect 7150 946 7189 998
rect 7059 906 7189 946
rect 6762 856 6800 902
rect 6576 843 6622 852
rect 6762 763 6846 856
rect 3833 732 5324 743
rect 3833 686 5173 732
rect 5313 686 5324 732
rect 3833 675 5324 686
rect 3833 667 5275 675
rect 3833 643 4409 667
rect 2929 431 3057 461
rect 2929 385 2971 431
rect 3017 385 3057 431
rect 2929 327 3057 385
rect 2929 275 2967 327
rect 3019 275 3057 327
rect 2929 235 3057 275
rect 3203 490 3279 502
rect 3203 230 3215 490
rect 3267 230 3279 490
rect 3442 383 3488 505
rect 3666 551 3712 564
rect 3666 502 3712 505
rect 3833 550 3961 643
rect 4099 554 4145 563
rect 3833 504 3875 550
rect 3921 504 3961 550
rect 4057 550 4185 554
rect 4057 512 4099 550
rect 3442 324 3488 337
rect 3651 490 3727 502
rect 3203 218 3279 230
rect 3651 230 3663 490
rect 3715 230 3727 490
rect 3651 218 3727 230
rect 3833 423 3961 504
rect 3833 377 3875 423
rect 3921 377 3961 423
rect 3833 296 3961 377
rect 3833 250 3875 296
rect 3921 250 3961 296
rect 3833 168 3961 250
rect 3833 122 3875 168
rect 3921 122 3961 168
rect 4056 504 4099 512
rect 4145 512 4185 550
rect 4281 550 4409 643
rect 4145 504 4186 512
rect 4056 471 4186 504
rect 4056 419 4095 471
rect 4147 419 4186 471
rect 4056 377 4099 419
rect 4145 377 4186 419
rect 4056 296 4186 377
rect 4056 253 4099 296
rect 4145 253 4186 296
rect 4056 201 4095 253
rect 4147 201 4186 253
rect 4056 168 4186 201
rect 4056 161 4099 168
rect 3833 117 3961 122
rect 4057 122 4099 161
rect 4145 161 4186 168
rect 4281 504 4323 550
rect 4369 504 4409 550
rect 4281 423 4409 504
rect 4281 377 4323 423
rect 4369 377 4409 423
rect 4281 296 4409 377
rect 4281 250 4323 296
rect 4369 250 4409 296
rect 4281 168 4409 250
rect 4543 427 4589 667
rect 5418 643 6846 763
rect 5232 555 5278 559
rect 4950 513 5078 554
rect 4543 307 4589 381
rect 4543 248 4589 261
rect 4725 471 4855 512
rect 4725 419 4764 471
rect 4816 419 4855 471
rect 4725 381 4767 419
rect 4813 381 4855 419
rect 4725 307 4855 381
rect 4725 261 4767 307
rect 4813 261 4855 307
rect 4725 253 4855 261
rect 4145 122 4185 161
rect 4057 117 4185 122
rect 4281 122 4323 168
rect 4369 122 4409 168
rect 4725 201 4764 253
rect 4816 201 4855 253
rect 4950 461 4988 513
rect 5040 461 5078 513
rect 4950 427 5078 461
rect 4950 381 4991 427
rect 5037 381 5078 427
rect 4950 327 5078 381
rect 4950 275 4988 327
rect 5040 275 5078 327
rect 4950 261 4991 275
rect 5037 261 5078 275
rect 4950 235 5078 261
rect 5190 546 5320 555
rect 5190 514 5232 546
rect 5278 514 5320 546
rect 5190 462 5229 514
rect 5281 462 5320 514
rect 5190 440 5320 462
rect 5190 394 5232 440
rect 5278 394 5320 440
rect 5190 296 5320 394
rect 5418 546 5534 643
rect 5680 555 5726 559
rect 5418 500 5456 546
rect 5502 500 5534 546
rect 5418 440 5534 500
rect 5418 394 5456 440
rect 5502 394 5534 440
rect 5418 389 5534 394
rect 5638 546 5768 555
rect 5638 514 5680 546
rect 5726 514 5768 546
rect 5638 462 5677 514
rect 5729 462 5768 514
rect 5638 440 5768 462
rect 5638 394 5680 440
rect 5726 394 5768 440
rect 5456 381 5502 389
rect 5190 244 5229 296
rect 5281 244 5320 296
rect 5190 204 5320 244
rect 5638 296 5768 394
rect 5866 546 5981 643
rect 6128 555 6174 559
rect 5866 500 5904 546
rect 5950 500 5981 546
rect 5866 440 5981 500
rect 5866 394 5904 440
rect 5950 394 5981 440
rect 5866 389 5981 394
rect 6086 546 6216 555
rect 6086 514 6128 546
rect 6174 514 6216 546
rect 6086 462 6125 514
rect 6177 462 6216 514
rect 6086 440 6216 462
rect 6086 394 6128 440
rect 6174 394 6216 440
rect 5904 381 5950 389
rect 5638 244 5677 296
rect 5729 244 5768 296
rect 5638 204 5768 244
rect 6086 296 6216 394
rect 6314 546 6429 643
rect 6576 555 6622 559
rect 6314 500 6352 546
rect 6398 500 6429 546
rect 6314 440 6429 500
rect 6314 394 6352 440
rect 6398 394 6429 440
rect 6314 389 6429 394
rect 6534 546 6664 555
rect 6534 514 6576 546
rect 6622 514 6664 546
rect 6534 462 6573 514
rect 6625 462 6664 514
rect 6534 440 6664 462
rect 6534 394 6576 440
rect 6622 394 6664 440
rect 6352 381 6398 389
rect 6086 244 6125 296
rect 6177 244 6216 296
rect 6086 204 6216 244
rect 6534 296 6664 394
rect 6800 546 6846 643
rect 6800 440 6846 500
rect 6800 381 6846 394
rect 7038 508 7218 520
rect 6534 244 6573 296
rect 6625 244 6664 296
rect 6534 204 6664 244
rect 7038 248 7050 508
rect 7206 248 7218 508
rect 7038 236 7218 248
rect 4725 161 4855 201
rect 4281 117 4409 122
rect 3875 109 3921 117
rect 4099 109 4145 117
rect 4323 109 4369 117
rect 1796 70 2609 81
rect 1796 24 2458 70
rect 2598 24 2609 70
rect 1796 13 2609 24
rect 2734 70 3463 81
rect 2734 24 3312 70
rect 3452 24 3463 70
rect 2734 13 3463 24
rect 4568 64 4730 75
rect 4568 18 4579 64
rect 4719 18 4730 64
rect 4568 7 4730 18
rect 3958 -18 4120 -7
rect 3958 -64 3969 -18
rect 4109 -64 4120 -18
rect 3958 -76 4120 -64
rect 366 -97 546 -85
rect 366 -149 378 -97
rect 534 -149 546 -97
rect 1330 -122 4120 -76
rect 366 -161 546 -149
rect 1696 -201 1858 -190
rect 4633 -201 4679 7
rect 1696 -247 1707 -201
rect 1847 -247 4679 -201
rect 1696 -258 1858 -247
<< via1 >>
rect 174 3492 226 3543
rect 174 3446 177 3492
rect 177 3446 223 3492
rect 223 3446 226 3492
rect 174 3383 226 3446
rect 174 3337 177 3383
rect 177 3337 223 3383
rect 223 3337 226 3383
rect 174 3283 226 3337
rect 622 3492 674 3543
rect 622 3446 625 3492
rect 625 3446 671 3492
rect 671 3446 674 3492
rect 622 3383 674 3446
rect 622 3337 625 3383
rect 625 3337 671 3383
rect 671 3337 674 3383
rect 622 3283 674 3337
rect 1303 3525 1563 3543
rect 1303 3291 1563 3525
rect 1303 3283 1563 3291
rect 1945 3539 1948 3543
rect 1948 3539 1994 3543
rect 1994 3539 1997 3543
rect 1945 3481 1997 3539
rect 1945 3435 1948 3481
rect 1948 3435 1994 3481
rect 1994 3435 1997 3481
rect 1945 3377 1997 3435
rect 1945 3331 1948 3377
rect 1948 3331 1994 3377
rect 1994 3331 1997 3377
rect 1945 3283 1997 3331
rect 2393 3539 2396 3543
rect 2396 3539 2442 3543
rect 2442 3539 2445 3543
rect 2393 3481 2445 3539
rect 2393 3435 2396 3481
rect 2396 3435 2442 3481
rect 2442 3435 2445 3481
rect 2393 3377 2445 3435
rect 2393 3331 2396 3377
rect 2396 3331 2442 3377
rect 2442 3331 2445 3377
rect 2393 3283 2445 3331
rect 2841 3539 2844 3543
rect 2844 3539 2890 3543
rect 2890 3539 2893 3543
rect 2841 3481 2893 3539
rect 2841 3435 2844 3481
rect 2844 3435 2890 3481
rect 2890 3435 2893 3481
rect 2841 3377 2893 3435
rect 2841 3331 2844 3377
rect 2844 3331 2890 3377
rect 2890 3331 2893 3377
rect 2841 3283 2893 3331
rect 2016 2988 2380 3040
rect 3289 3539 3292 3543
rect 3292 3539 3338 3543
rect 3338 3539 3341 3543
rect 3289 3481 3341 3539
rect 3289 3435 3292 3481
rect 3292 3435 3338 3481
rect 3338 3435 3341 3481
rect 3289 3377 3341 3435
rect 3289 3331 3292 3377
rect 3292 3331 3338 3377
rect 3338 3331 3341 3377
rect 3289 3283 3341 3331
rect 3737 3539 3740 3543
rect 3740 3539 3786 3543
rect 3786 3539 3789 3543
rect 3737 3481 3789 3539
rect 3737 3435 3740 3481
rect 3740 3435 3786 3481
rect 3786 3435 3789 3481
rect 3737 3377 3789 3435
rect 3737 3331 3740 3377
rect 3740 3331 3786 3377
rect 3786 3331 3789 3377
rect 3737 3283 3789 3331
rect 4185 3539 4188 3543
rect 4188 3539 4234 3543
rect 4234 3539 4237 3543
rect 4185 3481 4237 3539
rect 4185 3435 4188 3481
rect 4188 3435 4234 3481
rect 4234 3435 4237 3481
rect 4185 3377 4237 3435
rect 4185 3331 4188 3377
rect 4188 3331 4234 3377
rect 4234 3331 4237 3377
rect 4185 3283 4237 3331
rect 4388 3525 4440 3543
rect 4388 3291 4391 3525
rect 4391 3291 4437 3525
rect 4437 3291 4440 3525
rect 4388 3283 4440 3291
rect 4591 3539 4594 3543
rect 4594 3539 4640 3543
rect 4640 3539 4643 3543
rect 4591 3481 4643 3539
rect 4591 3435 4594 3481
rect 4594 3435 4640 3481
rect 4640 3435 4643 3481
rect 4591 3377 4643 3435
rect 4591 3331 4594 3377
rect 4594 3331 4640 3377
rect 4640 3331 4643 3377
rect 4591 3283 4643 3331
rect 5039 3539 5042 3543
rect 5042 3539 5088 3543
rect 5088 3539 5091 3543
rect 5039 3481 5091 3539
rect 5039 3435 5042 3481
rect 5042 3435 5088 3481
rect 5088 3435 5091 3481
rect 5039 3377 5091 3435
rect 5039 3331 5042 3377
rect 5042 3331 5088 3377
rect 5088 3331 5091 3377
rect 5039 3283 5091 3331
rect 174 2261 226 2267
rect 174 2215 177 2261
rect 177 2215 223 2261
rect 223 2215 226 2261
rect 174 2155 226 2215
rect 174 2109 177 2155
rect 177 2109 223 2155
rect 223 2109 226 2155
rect 174 2049 226 2109
rect 174 2007 177 2049
rect 177 2007 223 2049
rect 223 2007 226 2049
rect 622 2261 674 2267
rect 622 2215 625 2261
rect 625 2215 671 2261
rect 671 2215 674 2261
rect 622 2155 674 2215
rect 622 2109 625 2155
rect 625 2109 671 2155
rect 671 2109 674 2155
rect 622 2049 674 2109
rect 622 2007 625 2049
rect 625 2007 671 2049
rect 671 2007 674 2049
rect 1070 2261 1122 2267
rect 1070 2215 1073 2261
rect 1073 2215 1119 2261
rect 1119 2215 1122 2261
rect 1070 2155 1122 2215
rect 1070 2109 1073 2155
rect 1073 2109 1119 2155
rect 1119 2109 1122 2155
rect 1070 2049 1122 2109
rect 1070 2007 1073 2049
rect 1073 2007 1119 2049
rect 1119 2007 1122 2049
rect 1518 2261 1570 2267
rect 1518 2215 1521 2261
rect 1521 2215 1567 2261
rect 1567 2215 1570 2261
rect 1518 2155 1570 2215
rect 1518 2109 1521 2155
rect 1521 2109 1567 2155
rect 1567 2109 1570 2155
rect 1518 2049 1570 2109
rect 1518 2007 1521 2049
rect 1521 2007 1567 2049
rect 1567 2007 1570 2049
rect 1722 2249 1774 2267
rect 1722 2015 1725 2249
rect 1725 2015 1771 2249
rect 1771 2015 1774 2249
rect 1722 2007 1774 2015
rect 1945 2224 1948 2267
rect 1948 2224 1994 2267
rect 1994 2224 1997 2267
rect 1945 2161 1997 2224
rect 1945 2115 1948 2161
rect 1948 2115 1994 2161
rect 1994 2115 1997 2161
rect 1945 2052 1997 2115
rect 1945 2007 1948 2052
rect 1948 2007 1994 2052
rect 1994 2007 1997 2052
rect 2393 2224 2396 2267
rect 2396 2224 2442 2267
rect 2442 2224 2445 2267
rect 2393 2161 2445 2224
rect 2393 2115 2396 2161
rect 2396 2115 2442 2161
rect 2442 2115 2445 2161
rect 2393 2052 2445 2115
rect 2393 2007 2396 2052
rect 2396 2007 2442 2052
rect 2442 2007 2445 2052
rect 2841 2224 2844 2267
rect 2844 2224 2890 2267
rect 2890 2224 2893 2267
rect 2841 2161 2893 2224
rect 2841 2115 2844 2161
rect 2844 2115 2890 2161
rect 2890 2115 2893 2161
rect 2841 2052 2893 2115
rect 2841 2007 2844 2052
rect 2844 2007 2890 2052
rect 2890 2007 2893 2052
rect 3289 2224 3292 2267
rect 3292 2224 3338 2267
rect 3338 2224 3341 2267
rect 3289 2161 3341 2224
rect 3289 2115 3292 2161
rect 3292 2115 3338 2161
rect 3338 2115 3341 2161
rect 3289 2052 3341 2115
rect 3289 2007 3292 2052
rect 3292 2007 3338 2052
rect 3338 2007 3341 2052
rect 5487 3539 5490 3543
rect 5490 3539 5536 3543
rect 5536 3539 5539 3543
rect 5487 3481 5539 3539
rect 5487 3435 5490 3481
rect 5490 3435 5536 3481
rect 5536 3435 5539 3481
rect 5487 3377 5539 3435
rect 5487 3331 5490 3377
rect 5490 3331 5536 3377
rect 5536 3331 5539 3377
rect 5487 3283 5539 3331
rect 5935 3539 5938 3543
rect 5938 3539 5984 3543
rect 5984 3539 5987 3543
rect 5935 3481 5987 3539
rect 5935 3435 5938 3481
rect 5938 3435 5984 3481
rect 5984 3435 5987 3481
rect 5935 3377 5987 3435
rect 5935 3331 5938 3377
rect 5938 3331 5984 3377
rect 5984 3331 5987 3377
rect 5935 3283 5987 3331
rect 6383 3539 6386 3543
rect 6386 3539 6432 3543
rect 6432 3539 6435 3543
rect 6383 3481 6435 3539
rect 6383 3435 6386 3481
rect 6386 3435 6432 3481
rect 6432 3435 6435 3481
rect 6383 3377 6435 3435
rect 6383 3331 6386 3377
rect 6386 3331 6432 3377
rect 6432 3331 6435 3377
rect 6383 3283 6435 3331
rect 6831 3539 6834 3543
rect 6834 3539 6880 3543
rect 6880 3539 6883 3543
rect 6831 3481 6883 3539
rect 6831 3435 6834 3481
rect 6834 3435 6880 3481
rect 6880 3435 6883 3481
rect 6831 3377 6883 3435
rect 6831 3331 6834 3377
rect 6834 3331 6880 3377
rect 6880 3331 6883 3377
rect 6831 3283 6883 3331
rect 7050 3525 7206 3543
rect 7050 3291 7051 3525
rect 7051 3291 7191 3525
rect 7191 3291 7206 3525
rect 7050 3283 7206 3291
rect 3737 2224 3740 2267
rect 3740 2224 3786 2267
rect 3786 2224 3789 2267
rect 3737 2161 3789 2224
rect 3737 2115 3740 2161
rect 3740 2115 3786 2161
rect 3786 2115 3789 2161
rect 3737 2052 3789 2115
rect 3737 2007 3740 2052
rect 3740 2007 3786 2052
rect 3786 2007 3789 2052
rect 4185 2224 4188 2267
rect 4188 2224 4234 2267
rect 4234 2224 4237 2267
rect 4185 2161 4237 2224
rect 4185 2115 4188 2161
rect 4188 2115 4234 2161
rect 4234 2115 4237 2161
rect 4185 2052 4237 2115
rect 4185 2007 4188 2052
rect 4188 2007 4234 2052
rect 4234 2007 4237 2052
rect 4388 2249 4440 2267
rect 4388 2015 4391 2249
rect 4391 2015 4437 2249
rect 4437 2015 4440 2249
rect 4388 2007 4440 2015
rect 4591 2224 4594 2267
rect 4594 2224 4640 2267
rect 4640 2224 4643 2267
rect 4591 2161 4643 2224
rect 4591 2115 4594 2161
rect 4594 2115 4640 2161
rect 4640 2115 4643 2161
rect 4591 2052 4643 2115
rect 4591 2007 4594 2052
rect 4594 2007 4640 2052
rect 4640 2007 4643 2052
rect 5039 2224 5042 2267
rect 5042 2224 5088 2267
rect 5088 2224 5091 2267
rect 5039 2161 5091 2224
rect 5039 2115 5042 2161
rect 5042 2115 5088 2161
rect 5088 2115 5091 2161
rect 5039 2052 5091 2115
rect 5039 2007 5042 2052
rect 5042 2007 5088 2052
rect 5088 2007 5091 2052
rect 5487 2224 5490 2267
rect 5490 2224 5536 2267
rect 5536 2224 5539 2267
rect 5487 2161 5539 2224
rect 5487 2115 5490 2161
rect 5490 2115 5536 2161
rect 5536 2115 5539 2161
rect 5487 2052 5539 2115
rect 5487 2007 5490 2052
rect 5490 2007 5536 2052
rect 5536 2007 5539 2052
rect 5935 2224 5938 2267
rect 5938 2224 5984 2267
rect 5984 2224 5987 2267
rect 5935 2161 5987 2224
rect 5935 2115 5938 2161
rect 5938 2115 5984 2161
rect 5984 2115 5987 2161
rect 5935 2052 5987 2115
rect 5935 2007 5938 2052
rect 5938 2007 5984 2052
rect 5984 2007 5987 2052
rect 6383 2224 6386 2267
rect 6386 2224 6432 2267
rect 6432 2224 6435 2267
rect 6383 2161 6435 2224
rect 6383 2115 6386 2161
rect 6386 2115 6432 2161
rect 6432 2115 6435 2161
rect 6383 2052 6435 2115
rect 6383 2007 6386 2052
rect 6386 2007 6432 2052
rect 6432 2007 6435 2052
rect 6831 2224 6834 2267
rect 6834 2224 6880 2267
rect 6880 2224 6883 2267
rect 6831 2161 6883 2224
rect 6831 2115 6834 2161
rect 6834 2115 6880 2161
rect 6880 2115 6883 2161
rect 6831 2052 6883 2115
rect 6831 2007 6834 2052
rect 6834 2007 6880 2052
rect 6880 2007 6883 2052
rect 7044 2249 7200 2267
rect 7044 2015 7051 2249
rect 7051 2015 7191 2249
rect 7191 2015 7200 2249
rect 7044 2007 7200 2015
rect 130 1186 182 1216
rect 130 1164 133 1186
rect 133 1164 179 1186
rect 179 1164 182 1186
rect 130 976 133 998
rect 133 976 179 998
rect 179 976 182 998
rect 130 946 182 976
rect 1274 1435 1430 1487
rect 655 1157 707 1205
rect 655 1153 658 1157
rect 658 1153 704 1157
rect 704 1153 707 1157
rect 655 984 658 987
rect 658 984 704 987
rect 704 984 707 987
rect 655 935 707 984
rect 130 484 182 514
rect 130 462 133 484
rect 133 462 179 484
rect 179 462 182 484
rect 130 274 133 296
rect 133 274 179 296
rect 179 274 182 296
rect 130 244 182 274
rect 1103 1157 1155 1205
rect 1103 1153 1106 1157
rect 1106 1153 1152 1157
rect 1152 1153 1155 1157
rect 1103 984 1106 987
rect 1106 984 1152 987
rect 1152 984 1155 987
rect 1103 935 1155 984
rect 1610 1157 1662 1164
rect 1610 1112 1613 1157
rect 1613 1112 1659 1157
rect 1659 1112 1662 1157
rect 1610 902 1662 947
rect 1610 895 1613 902
rect 1613 895 1659 902
rect 1659 895 1662 902
rect 1610 677 1662 729
rect 655 462 707 514
rect 655 272 707 296
rect 655 244 658 272
rect 658 244 704 272
rect 704 244 707 272
rect 1103 474 1155 513
rect 1103 461 1106 474
rect 1106 461 1152 474
rect 1152 461 1155 474
rect 1103 308 1106 327
rect 1106 308 1152 327
rect 1152 308 1155 327
rect 1103 275 1155 308
rect 670 3 722 55
rect 882 38 892 55
rect 892 38 934 55
rect 882 3 934 38
rect 1610 504 1613 511
rect 1613 504 1659 511
rect 1659 504 1662 511
rect 1610 459 1662 504
rect 1610 250 1613 294
rect 1613 250 1659 294
rect 1659 250 1662 294
rect 1610 242 1662 250
rect 2519 1157 2571 1205
rect 2519 1153 2523 1157
rect 2523 1153 2569 1157
rect 2569 1153 2571 1157
rect 2519 984 2523 987
rect 2523 984 2569 987
rect 2569 984 2571 987
rect 2519 935 2571 984
rect 2967 1157 3019 1205
rect 2967 1153 2971 1157
rect 2971 1153 3017 1157
rect 3017 1153 3019 1157
rect 2967 984 2971 987
rect 2971 984 3017 987
rect 3017 984 3019 987
rect 2967 935 3019 984
rect 3215 1150 3267 1219
rect 3215 1104 3218 1150
rect 3218 1104 3264 1150
rect 3264 1104 3267 1150
rect 3215 1026 3267 1104
rect 3215 980 3218 1026
rect 3218 980 3264 1026
rect 3264 980 3267 1026
rect 3215 959 3267 980
rect 4602 1480 4758 1487
rect 4602 1435 4608 1480
rect 4608 1435 4748 1480
rect 4748 1435 4758 1480
rect 3663 1150 3715 1219
rect 3663 1104 3666 1150
rect 3666 1104 3712 1150
rect 3712 1104 3715 1150
rect 3663 1026 3715 1104
rect 3663 980 3666 1026
rect 3666 980 3712 1026
rect 3712 980 3715 1026
rect 3663 959 3715 980
rect 2519 505 2523 513
rect 2523 505 2569 513
rect 2569 505 2571 513
rect 2519 461 2571 505
rect 2519 275 2571 327
rect 2967 505 2971 513
rect 2971 505 3017 513
rect 3017 505 3019 513
rect 2967 461 3019 505
rect 4095 1157 4147 1205
rect 4095 1153 4099 1157
rect 4099 1153 4145 1157
rect 4145 1153 4147 1157
rect 4095 984 4099 987
rect 4099 984 4145 987
rect 4145 984 4147 987
rect 4095 935 4147 984
rect 4764 1156 4816 1205
rect 4764 1153 4767 1156
rect 4767 1153 4813 1156
rect 4813 1153 4816 1156
rect 4764 983 4767 987
rect 4767 983 4813 987
rect 4813 983 4816 987
rect 4764 935 4816 983
rect 4988 1156 5040 1205
rect 4988 1153 4991 1156
rect 4991 1153 5037 1156
rect 5037 1153 5040 1156
rect 4988 983 4991 987
rect 4991 983 5037 987
rect 5037 983 5040 987
rect 4988 935 5040 983
rect 5229 1162 5281 1214
rect 5229 979 5232 996
rect 5232 979 5278 996
rect 5278 979 5281 996
rect 5229 944 5281 979
rect 5677 1162 5729 1214
rect 5677 979 5680 996
rect 5680 979 5726 996
rect 5726 979 5729 996
rect 5677 944 5729 979
rect 6125 1162 6177 1214
rect 6125 979 6128 996
rect 6128 979 6174 996
rect 6174 979 6177 996
rect 6125 944 6177 979
rect 6573 1162 6625 1214
rect 6573 979 6576 996
rect 6576 979 6622 996
rect 6622 979 6625 996
rect 6573 944 6625 979
rect 7098 1186 7150 1216
rect 7098 1164 7101 1186
rect 7101 1164 7147 1186
rect 7147 1164 7150 1186
rect 7098 976 7101 998
rect 7101 976 7147 998
rect 7147 976 7150 998
rect 7098 946 7150 976
rect 2967 275 3019 327
rect 3215 383 3267 490
rect 3215 337 3218 383
rect 3218 337 3264 383
rect 3264 337 3267 383
rect 3215 230 3267 337
rect 3663 383 3715 490
rect 3663 337 3666 383
rect 3666 337 3712 383
rect 3712 337 3715 383
rect 3663 230 3715 337
rect 4095 423 4147 471
rect 4095 419 4099 423
rect 4099 419 4145 423
rect 4145 419 4147 423
rect 4095 250 4099 253
rect 4099 250 4145 253
rect 4145 250 4147 253
rect 4095 201 4147 250
rect 4764 427 4816 471
rect 4764 419 4767 427
rect 4767 419 4813 427
rect 4813 419 4816 427
rect 4764 201 4816 253
rect 4988 461 5040 513
rect 4988 307 5040 327
rect 4988 275 4991 307
rect 4991 275 5037 307
rect 5037 275 5040 307
rect 5229 500 5232 514
rect 5232 500 5278 514
rect 5278 500 5281 514
rect 5229 462 5281 500
rect 5677 500 5680 514
rect 5680 500 5726 514
rect 5726 500 5729 514
rect 5677 462 5729 500
rect 5229 244 5281 296
rect 6125 500 6128 514
rect 6128 500 6174 514
rect 6174 500 6177 514
rect 6125 462 6177 500
rect 5677 244 5729 296
rect 6573 500 6576 514
rect 6576 500 6622 514
rect 6622 500 6625 514
rect 6573 462 6625 500
rect 6125 244 6177 296
rect 6573 244 6625 296
rect 7050 490 7206 508
rect 7050 256 7051 490
rect 7051 256 7191 490
rect 7191 256 7206 490
rect 7050 248 7206 256
rect 378 -149 534 -97
<< metal2 >>
rect 162 3545 238 3555
rect 162 3281 172 3545
rect 228 3281 238 3545
rect 162 3271 238 3281
rect 610 3545 686 3555
rect 610 3281 620 3545
rect 676 3281 686 3545
rect 610 3271 686 3281
rect 1291 3545 1575 3555
rect 1291 3281 1301 3545
rect 1565 3281 1575 3545
rect 1291 3271 1575 3281
rect 1933 3545 2009 3555
rect 1933 3281 1943 3545
rect 1999 3281 2009 3545
rect 1933 3271 2009 3281
rect 2381 3545 2457 3555
rect 2381 3281 2391 3545
rect 2447 3281 2457 3545
rect 2381 3271 2457 3281
rect 2829 3545 2905 3555
rect 2829 3281 2839 3545
rect 2895 3281 2905 3545
rect 2829 3271 2905 3281
rect 3277 3545 3353 3555
rect 3277 3281 3287 3545
rect 3343 3281 3353 3545
rect 3277 3271 3353 3281
rect 3725 3545 3801 3555
rect 3725 3281 3735 3545
rect 3791 3281 3801 3545
rect 3725 3271 3801 3281
rect 4173 3545 4249 3555
rect 4173 3281 4183 3545
rect 4239 3281 4249 3545
rect 4173 3271 4249 3281
rect 4376 3545 4452 3555
rect 4376 3281 4386 3545
rect 4442 3281 4452 3545
rect 4376 3271 4452 3281
rect 4579 3545 4655 3555
rect 4579 3281 4589 3545
rect 4645 3281 4655 3545
rect 4579 3271 4655 3281
rect 5027 3545 5103 3555
rect 5027 3281 5037 3545
rect 5093 3281 5103 3545
rect 5027 3271 5103 3281
rect 5475 3545 5551 3555
rect 5475 3281 5485 3545
rect 5541 3281 5551 3545
rect 5475 3271 5551 3281
rect 5923 3545 5999 3555
rect 5923 3281 5933 3545
rect 5989 3281 5999 3545
rect 5923 3271 5999 3281
rect 6371 3545 6447 3555
rect 6371 3281 6381 3545
rect 6437 3281 6447 3545
rect 6371 3271 6447 3281
rect 6819 3545 6895 3555
rect 6819 3281 6829 3545
rect 6885 3281 6895 3545
rect 6819 3271 6895 3281
rect 7038 3545 7218 3555
rect 7038 3281 7048 3545
rect 7208 3281 7218 3545
rect 7038 3271 7218 3281
rect 2004 3042 2392 3052
rect 2004 2986 2014 3042
rect 2382 2986 2392 3042
rect 2004 2976 2392 2986
rect 162 2269 238 2279
rect 162 2005 172 2269
rect 228 2005 238 2269
rect 162 1995 238 2005
rect 610 2269 686 2279
rect 610 2005 620 2269
rect 676 2005 686 2269
rect 610 1995 686 2005
rect 1058 2269 1134 2279
rect 1058 2005 1068 2269
rect 1124 2005 1134 2269
rect 1058 1995 1134 2005
rect 1506 2269 1582 2279
rect 1506 2005 1516 2269
rect 1572 2005 1582 2269
rect 1506 1995 1582 2005
rect 1710 2269 1786 2279
rect 1710 2005 1720 2269
rect 1776 2005 1786 2269
rect 1710 1995 1786 2005
rect 1933 2269 2009 2279
rect 1933 2005 1943 2269
rect 1999 2005 2009 2269
rect 1933 1995 2009 2005
rect 2381 2269 2457 2279
rect 2381 2005 2391 2269
rect 2447 2005 2457 2269
rect 2381 1995 2457 2005
rect 2829 2269 2905 2279
rect 2829 2005 2839 2269
rect 2895 2005 2905 2269
rect 2829 1995 2905 2005
rect 3277 2269 3353 2279
rect 3277 2005 3287 2269
rect 3343 2005 3353 2269
rect 3277 1995 3353 2005
rect 3725 2269 3801 2279
rect 3725 2005 3735 2269
rect 3791 2005 3801 2269
rect 3725 1995 3801 2005
rect 4173 2269 4249 2279
rect 4173 2005 4183 2269
rect 4239 2005 4249 2269
rect 4173 1995 4249 2005
rect 4376 2269 4452 2279
rect 4376 2005 4386 2269
rect 4442 2005 4452 2269
rect 4376 1995 4452 2005
rect 4579 2269 4655 2279
rect 4579 2005 4589 2269
rect 4645 2005 4655 2269
rect 4579 1995 4655 2005
rect 5027 2269 5103 2279
rect 5027 2005 5037 2269
rect 5093 2005 5103 2269
rect 5027 1995 5103 2005
rect 5475 2269 5551 2279
rect 5475 2005 5485 2269
rect 5541 2005 5551 2269
rect 5475 1995 5551 2005
rect 5923 2269 5999 2279
rect 5923 2005 5933 2269
rect 5989 2005 5999 2269
rect 5923 1995 5999 2005
rect 6371 2269 6447 2279
rect 6371 2005 6381 2269
rect 6437 2005 6447 2269
rect 6371 1995 6447 2005
rect 6819 2269 6895 2279
rect 6819 2005 6829 2269
rect 6885 2005 6895 2269
rect 6819 1995 6895 2005
rect 7032 2269 7212 2279
rect 7032 2005 7042 2269
rect 7202 2005 7212 2269
rect 7032 1995 7212 2005
rect 1262 1489 1442 1499
rect 1262 1433 1272 1489
rect 1432 1433 1442 1489
rect 1262 1423 1442 1433
rect 4590 1489 4770 1499
rect 4590 1433 4600 1489
rect 4760 1433 4770 1489
rect 4590 1423 4770 1433
rect 91 1218 221 1257
rect 91 1162 128 1218
rect 184 1162 221 1218
rect 91 1000 221 1162
rect 91 944 128 1000
rect 184 944 221 1000
rect 91 906 221 944
rect 616 1207 746 1246
rect 616 1151 653 1207
rect 709 1151 746 1207
rect 616 989 746 1151
rect 616 933 653 989
rect 709 933 746 989
rect 616 895 746 933
rect 1064 1207 1194 1246
rect 1064 1151 1101 1207
rect 1157 1151 1194 1207
rect 1064 989 1194 1151
rect 1064 933 1101 989
rect 1157 933 1194 989
rect 1064 895 1194 933
rect 1572 1164 1700 1289
rect 4057 1246 4185 1289
rect 4726 1246 4854 1289
rect 1572 1112 1610 1164
rect 1662 1112 1700 1164
rect 1572 947 1700 1112
rect 1572 895 1610 947
rect 1662 895 1700 947
rect 2480 1207 2610 1246
rect 2480 1151 2517 1207
rect 2573 1151 2610 1207
rect 2480 989 2610 1151
rect 2480 933 2517 989
rect 2573 933 2610 989
rect 2480 895 2610 933
rect 2928 1207 3058 1246
rect 2928 1151 2965 1207
rect 3021 1151 3058 1207
rect 2928 989 3058 1151
rect 2928 933 2965 989
rect 3021 933 3058 989
rect 3203 1221 3279 1231
rect 3203 957 3213 1221
rect 3269 957 3279 1221
rect 3203 947 3279 957
rect 3651 1221 3727 1231
rect 3651 957 3661 1221
rect 3717 957 3727 1221
rect 3651 947 3727 957
rect 4056 1205 4186 1246
rect 4056 1153 4095 1205
rect 4147 1153 4186 1205
rect 4056 987 4186 1153
rect 2928 895 3058 933
rect 4056 935 4095 987
rect 4147 935 4186 987
rect 4056 895 4186 935
rect 4725 1205 4855 1246
rect 4725 1153 4764 1205
rect 4816 1153 4855 1205
rect 4725 987 4855 1153
rect 4725 935 4764 987
rect 4816 935 4855 987
rect 4725 895 4855 935
rect 4949 1207 5079 1246
rect 4949 1151 4986 1207
rect 5042 1151 5079 1207
rect 4949 989 5079 1151
rect 4949 933 4986 989
rect 5042 933 5079 989
rect 4949 895 5079 933
rect 5190 1216 5320 1254
rect 5190 1160 5227 1216
rect 5283 1160 5320 1216
rect 5190 998 5320 1160
rect 5190 942 5227 998
rect 5283 942 5320 998
rect 5190 903 5320 942
rect 5638 1216 5768 1254
rect 5638 1160 5675 1216
rect 5731 1160 5768 1216
rect 5638 998 5768 1160
rect 5638 942 5675 998
rect 5731 942 5768 998
rect 5638 903 5768 942
rect 6086 1216 6216 1254
rect 6086 1160 6123 1216
rect 6179 1160 6216 1216
rect 6086 998 6216 1160
rect 6086 942 6123 998
rect 6179 942 6216 998
rect 6086 903 6216 942
rect 6534 1216 6664 1254
rect 6534 1160 6571 1216
rect 6627 1160 6664 1216
rect 6534 998 6664 1160
rect 6534 942 6571 998
rect 6627 942 6664 998
rect 6534 903 6664 942
rect 7059 1218 7189 1257
rect 7059 1162 7096 1218
rect 7152 1162 7189 1218
rect 7059 1000 7189 1162
rect 7059 944 7096 1000
rect 7152 944 7189 1000
rect 7059 906 7189 944
rect 1572 729 1700 895
rect 1572 677 1610 729
rect 1662 677 1700 729
rect 91 516 221 555
rect 91 460 128 516
rect 184 460 221 516
rect 91 298 221 460
rect 91 242 128 298
rect 184 242 221 298
rect 91 204 221 242
rect 616 516 746 555
rect 616 460 653 516
rect 709 460 746 516
rect 616 298 746 460
rect 616 242 653 298
rect 709 242 746 298
rect 616 204 746 242
rect 1065 515 1193 554
rect 1065 459 1101 515
rect 1157 459 1193 515
rect 1065 329 1193 459
rect 1065 273 1101 329
rect 1157 273 1193 329
rect 1065 235 1193 273
rect 1572 511 1700 677
rect 1572 459 1610 511
rect 1662 459 1700 511
rect 1572 294 1700 459
rect 1572 242 1610 294
rect 1662 242 1700 294
rect 1572 201 1700 242
rect 2481 515 2609 554
rect 2481 459 2517 515
rect 2573 459 2609 515
rect 2481 329 2609 459
rect 2481 273 2517 329
rect 2573 273 2609 329
rect 2481 235 2609 273
rect 2929 515 3057 554
rect 2929 459 2965 515
rect 3021 459 3057 515
rect 4057 512 4185 895
rect 4726 512 4854 895
rect 4950 515 5078 554
rect 2929 329 3057 459
rect 2929 273 2965 329
rect 3021 273 3057 329
rect 2929 235 3057 273
rect 3203 492 3279 502
rect 3203 228 3213 492
rect 3269 228 3279 492
rect 3203 218 3279 228
rect 3651 492 3727 502
rect 3651 228 3661 492
rect 3717 228 3727 492
rect 3651 218 3727 228
rect 4056 471 4186 512
rect 4056 419 4095 471
rect 4147 419 4186 471
rect 4056 253 4186 419
rect 4056 201 4095 253
rect 4147 201 4186 253
rect 632 56 972 96
rect 632 0 668 56
rect 724 0 880 56
rect 936 0 972 56
rect 632 -38 972 0
rect 366 -94 546 -85
rect 1608 -94 1664 201
rect 4056 161 4186 201
rect 4725 471 4855 512
rect 4725 419 4764 471
rect 4816 419 4855 471
rect 4725 253 4855 419
rect 4725 201 4764 253
rect 4816 201 4855 253
rect 4950 459 4986 515
rect 5042 459 5078 515
rect 4950 329 5078 459
rect 4950 273 4986 329
rect 5042 273 5078 329
rect 4950 235 5078 273
rect 5190 516 5320 555
rect 5190 460 5227 516
rect 5283 460 5320 516
rect 5190 298 5320 460
rect 5190 242 5227 298
rect 5283 242 5320 298
rect 5190 204 5320 242
rect 5638 516 5768 555
rect 5638 460 5675 516
rect 5731 460 5768 516
rect 5638 298 5768 460
rect 5638 242 5675 298
rect 5731 242 5768 298
rect 5638 204 5768 242
rect 6086 516 6216 555
rect 6086 460 6123 516
rect 6179 460 6216 516
rect 6086 298 6216 460
rect 6086 242 6123 298
rect 6179 242 6216 298
rect 6086 204 6216 242
rect 6534 516 6664 555
rect 6534 460 6571 516
rect 6627 460 6664 516
rect 6534 298 6664 460
rect 6534 242 6571 298
rect 6627 242 6664 298
rect 6534 204 6664 242
rect 7038 510 7218 520
rect 7038 246 7048 510
rect 7208 246 7218 510
rect 7038 236 7218 246
rect 4725 161 4855 201
rect 4057 117 4185 161
rect 4726 117 4854 161
rect 366 -97 1664 -94
rect 366 -149 378 -97
rect 534 -149 1664 -97
rect 366 -150 1664 -149
rect 366 -161 546 -150
<< via2 >>
rect 172 3543 228 3545
rect 172 3283 174 3543
rect 174 3283 226 3543
rect 226 3283 228 3543
rect 172 3281 228 3283
rect 620 3543 676 3545
rect 620 3283 622 3543
rect 622 3283 674 3543
rect 674 3283 676 3543
rect 620 3281 676 3283
rect 1301 3543 1565 3545
rect 1301 3283 1303 3543
rect 1303 3283 1563 3543
rect 1563 3283 1565 3543
rect 1301 3281 1565 3283
rect 1943 3543 1999 3545
rect 1943 3283 1945 3543
rect 1945 3283 1997 3543
rect 1997 3283 1999 3543
rect 1943 3281 1999 3283
rect 2391 3543 2447 3545
rect 2391 3283 2393 3543
rect 2393 3283 2445 3543
rect 2445 3283 2447 3543
rect 2391 3281 2447 3283
rect 2839 3543 2895 3545
rect 2839 3283 2841 3543
rect 2841 3283 2893 3543
rect 2893 3283 2895 3543
rect 2839 3281 2895 3283
rect 3287 3543 3343 3545
rect 3287 3283 3289 3543
rect 3289 3283 3341 3543
rect 3341 3283 3343 3543
rect 3287 3281 3343 3283
rect 3735 3543 3791 3545
rect 3735 3283 3737 3543
rect 3737 3283 3789 3543
rect 3789 3283 3791 3543
rect 3735 3281 3791 3283
rect 4183 3543 4239 3545
rect 4183 3283 4185 3543
rect 4185 3283 4237 3543
rect 4237 3283 4239 3543
rect 4183 3281 4239 3283
rect 4386 3543 4442 3545
rect 4386 3283 4388 3543
rect 4388 3283 4440 3543
rect 4440 3283 4442 3543
rect 4386 3281 4442 3283
rect 4589 3543 4645 3545
rect 4589 3283 4591 3543
rect 4591 3283 4643 3543
rect 4643 3283 4645 3543
rect 4589 3281 4645 3283
rect 5037 3543 5093 3545
rect 5037 3283 5039 3543
rect 5039 3283 5091 3543
rect 5091 3283 5093 3543
rect 5037 3281 5093 3283
rect 5485 3543 5541 3545
rect 5485 3283 5487 3543
rect 5487 3283 5539 3543
rect 5539 3283 5541 3543
rect 5485 3281 5541 3283
rect 5933 3543 5989 3545
rect 5933 3283 5935 3543
rect 5935 3283 5987 3543
rect 5987 3283 5989 3543
rect 5933 3281 5989 3283
rect 6381 3543 6437 3545
rect 6381 3283 6383 3543
rect 6383 3283 6435 3543
rect 6435 3283 6437 3543
rect 6381 3281 6437 3283
rect 6829 3543 6885 3545
rect 6829 3283 6831 3543
rect 6831 3283 6883 3543
rect 6883 3283 6885 3543
rect 6829 3281 6885 3283
rect 7048 3543 7208 3545
rect 7048 3283 7050 3543
rect 7050 3283 7206 3543
rect 7206 3283 7208 3543
rect 7048 3281 7208 3283
rect 2014 3040 2382 3042
rect 2014 2988 2016 3040
rect 2016 2988 2380 3040
rect 2380 2988 2382 3040
rect 2014 2986 2382 2988
rect 172 2267 228 2269
rect 172 2007 174 2267
rect 174 2007 226 2267
rect 226 2007 228 2267
rect 172 2005 228 2007
rect 620 2267 676 2269
rect 620 2007 622 2267
rect 622 2007 674 2267
rect 674 2007 676 2267
rect 620 2005 676 2007
rect 1068 2267 1124 2269
rect 1068 2007 1070 2267
rect 1070 2007 1122 2267
rect 1122 2007 1124 2267
rect 1068 2005 1124 2007
rect 1516 2267 1572 2269
rect 1516 2007 1518 2267
rect 1518 2007 1570 2267
rect 1570 2007 1572 2267
rect 1516 2005 1572 2007
rect 1720 2267 1776 2269
rect 1720 2007 1722 2267
rect 1722 2007 1774 2267
rect 1774 2007 1776 2267
rect 1720 2005 1776 2007
rect 1943 2267 1999 2269
rect 1943 2007 1945 2267
rect 1945 2007 1997 2267
rect 1997 2007 1999 2267
rect 1943 2005 1999 2007
rect 2391 2267 2447 2269
rect 2391 2007 2393 2267
rect 2393 2007 2445 2267
rect 2445 2007 2447 2267
rect 2391 2005 2447 2007
rect 2839 2267 2895 2269
rect 2839 2007 2841 2267
rect 2841 2007 2893 2267
rect 2893 2007 2895 2267
rect 2839 2005 2895 2007
rect 3287 2267 3343 2269
rect 3287 2007 3289 2267
rect 3289 2007 3341 2267
rect 3341 2007 3343 2267
rect 3287 2005 3343 2007
rect 3735 2267 3791 2269
rect 3735 2007 3737 2267
rect 3737 2007 3789 2267
rect 3789 2007 3791 2267
rect 3735 2005 3791 2007
rect 4183 2267 4239 2269
rect 4183 2007 4185 2267
rect 4185 2007 4237 2267
rect 4237 2007 4239 2267
rect 4183 2005 4239 2007
rect 4386 2267 4442 2269
rect 4386 2007 4388 2267
rect 4388 2007 4440 2267
rect 4440 2007 4442 2267
rect 4386 2005 4442 2007
rect 4589 2267 4645 2269
rect 4589 2007 4591 2267
rect 4591 2007 4643 2267
rect 4643 2007 4645 2267
rect 4589 2005 4645 2007
rect 5037 2267 5093 2269
rect 5037 2007 5039 2267
rect 5039 2007 5091 2267
rect 5091 2007 5093 2267
rect 5037 2005 5093 2007
rect 5485 2267 5541 2269
rect 5485 2007 5487 2267
rect 5487 2007 5539 2267
rect 5539 2007 5541 2267
rect 5485 2005 5541 2007
rect 5933 2267 5989 2269
rect 5933 2007 5935 2267
rect 5935 2007 5987 2267
rect 5987 2007 5989 2267
rect 5933 2005 5989 2007
rect 6381 2267 6437 2269
rect 6381 2007 6383 2267
rect 6383 2007 6435 2267
rect 6435 2007 6437 2267
rect 6381 2005 6437 2007
rect 6829 2267 6885 2269
rect 6829 2007 6831 2267
rect 6831 2007 6883 2267
rect 6883 2007 6885 2267
rect 6829 2005 6885 2007
rect 7042 2267 7202 2269
rect 7042 2007 7044 2267
rect 7044 2007 7200 2267
rect 7200 2007 7202 2267
rect 7042 2005 7202 2007
rect 1272 1487 1432 1489
rect 1272 1435 1274 1487
rect 1274 1435 1430 1487
rect 1430 1435 1432 1487
rect 1272 1433 1432 1435
rect 4600 1487 4760 1489
rect 4600 1435 4602 1487
rect 4602 1435 4758 1487
rect 4758 1435 4760 1487
rect 4600 1433 4760 1435
rect 128 1216 184 1218
rect 128 1164 130 1216
rect 130 1164 182 1216
rect 182 1164 184 1216
rect 128 1162 184 1164
rect 128 998 184 1000
rect 128 946 130 998
rect 130 946 182 998
rect 182 946 184 998
rect 128 944 184 946
rect 653 1205 709 1207
rect 653 1153 655 1205
rect 655 1153 707 1205
rect 707 1153 709 1205
rect 653 1151 709 1153
rect 653 987 709 989
rect 653 935 655 987
rect 655 935 707 987
rect 707 935 709 987
rect 653 933 709 935
rect 1101 1205 1157 1207
rect 1101 1153 1103 1205
rect 1103 1153 1155 1205
rect 1155 1153 1157 1205
rect 1101 1151 1157 1153
rect 1101 987 1157 989
rect 1101 935 1103 987
rect 1103 935 1155 987
rect 1155 935 1157 987
rect 1101 933 1157 935
rect 2517 1205 2573 1207
rect 2517 1153 2519 1205
rect 2519 1153 2571 1205
rect 2571 1153 2573 1205
rect 2517 1151 2573 1153
rect 2517 987 2573 989
rect 2517 935 2519 987
rect 2519 935 2571 987
rect 2571 935 2573 987
rect 2517 933 2573 935
rect 2965 1205 3021 1207
rect 2965 1153 2967 1205
rect 2967 1153 3019 1205
rect 3019 1153 3021 1205
rect 2965 1151 3021 1153
rect 2965 987 3021 989
rect 2965 935 2967 987
rect 2967 935 3019 987
rect 3019 935 3021 987
rect 2965 933 3021 935
rect 3213 1219 3269 1221
rect 3213 959 3215 1219
rect 3215 959 3267 1219
rect 3267 959 3269 1219
rect 3213 957 3269 959
rect 3661 1219 3717 1221
rect 3661 959 3663 1219
rect 3663 959 3715 1219
rect 3715 959 3717 1219
rect 3661 957 3717 959
rect 4986 1205 5042 1207
rect 4986 1153 4988 1205
rect 4988 1153 5040 1205
rect 5040 1153 5042 1205
rect 4986 1151 5042 1153
rect 4986 987 5042 989
rect 4986 935 4988 987
rect 4988 935 5040 987
rect 5040 935 5042 987
rect 4986 933 5042 935
rect 5227 1214 5283 1216
rect 5227 1162 5229 1214
rect 5229 1162 5281 1214
rect 5281 1162 5283 1214
rect 5227 1160 5283 1162
rect 5227 996 5283 998
rect 5227 944 5229 996
rect 5229 944 5281 996
rect 5281 944 5283 996
rect 5227 942 5283 944
rect 5675 1214 5731 1216
rect 5675 1162 5677 1214
rect 5677 1162 5729 1214
rect 5729 1162 5731 1214
rect 5675 1160 5731 1162
rect 5675 996 5731 998
rect 5675 944 5677 996
rect 5677 944 5729 996
rect 5729 944 5731 996
rect 5675 942 5731 944
rect 6123 1214 6179 1216
rect 6123 1162 6125 1214
rect 6125 1162 6177 1214
rect 6177 1162 6179 1214
rect 6123 1160 6179 1162
rect 6123 996 6179 998
rect 6123 944 6125 996
rect 6125 944 6177 996
rect 6177 944 6179 996
rect 6123 942 6179 944
rect 6571 1214 6627 1216
rect 6571 1162 6573 1214
rect 6573 1162 6625 1214
rect 6625 1162 6627 1214
rect 6571 1160 6627 1162
rect 6571 996 6627 998
rect 6571 944 6573 996
rect 6573 944 6625 996
rect 6625 944 6627 996
rect 6571 942 6627 944
rect 7096 1216 7152 1218
rect 7096 1164 7098 1216
rect 7098 1164 7150 1216
rect 7150 1164 7152 1216
rect 7096 1162 7152 1164
rect 7096 998 7152 1000
rect 7096 946 7098 998
rect 7098 946 7150 998
rect 7150 946 7152 998
rect 7096 944 7152 946
rect 128 514 184 516
rect 128 462 130 514
rect 130 462 182 514
rect 182 462 184 514
rect 128 460 184 462
rect 128 296 184 298
rect 128 244 130 296
rect 130 244 182 296
rect 182 244 184 296
rect 128 242 184 244
rect 653 514 709 516
rect 653 462 655 514
rect 655 462 707 514
rect 707 462 709 514
rect 653 460 709 462
rect 653 296 709 298
rect 653 244 655 296
rect 655 244 707 296
rect 707 244 709 296
rect 653 242 709 244
rect 1101 513 1157 515
rect 1101 461 1103 513
rect 1103 461 1155 513
rect 1155 461 1157 513
rect 1101 459 1157 461
rect 1101 327 1157 329
rect 1101 275 1103 327
rect 1103 275 1155 327
rect 1155 275 1157 327
rect 1101 273 1157 275
rect 2517 513 2573 515
rect 2517 461 2519 513
rect 2519 461 2571 513
rect 2571 461 2573 513
rect 2517 459 2573 461
rect 2517 327 2573 329
rect 2517 275 2519 327
rect 2519 275 2571 327
rect 2571 275 2573 327
rect 2517 273 2573 275
rect 2965 513 3021 515
rect 2965 461 2967 513
rect 2967 461 3019 513
rect 3019 461 3021 513
rect 2965 459 3021 461
rect 2965 327 3021 329
rect 2965 275 2967 327
rect 2967 275 3019 327
rect 3019 275 3021 327
rect 2965 273 3021 275
rect 3213 490 3269 492
rect 3213 230 3215 490
rect 3215 230 3267 490
rect 3267 230 3269 490
rect 3213 228 3269 230
rect 3661 490 3717 492
rect 3661 230 3663 490
rect 3663 230 3715 490
rect 3715 230 3717 490
rect 3661 228 3717 230
rect 668 55 724 56
rect 668 3 670 55
rect 670 3 722 55
rect 722 3 724 55
rect 668 0 724 3
rect 880 55 936 56
rect 880 3 882 55
rect 882 3 934 55
rect 934 3 936 55
rect 880 0 936 3
rect 4986 513 5042 515
rect 4986 461 4988 513
rect 4988 461 5040 513
rect 5040 461 5042 513
rect 4986 459 5042 461
rect 4986 327 5042 329
rect 4986 275 4988 327
rect 4988 275 5040 327
rect 5040 275 5042 327
rect 4986 273 5042 275
rect 5227 514 5283 516
rect 5227 462 5229 514
rect 5229 462 5281 514
rect 5281 462 5283 514
rect 5227 460 5283 462
rect 5227 296 5283 298
rect 5227 244 5229 296
rect 5229 244 5281 296
rect 5281 244 5283 296
rect 5227 242 5283 244
rect 5675 514 5731 516
rect 5675 462 5677 514
rect 5677 462 5729 514
rect 5729 462 5731 514
rect 5675 460 5731 462
rect 5675 296 5731 298
rect 5675 244 5677 296
rect 5677 244 5729 296
rect 5729 244 5731 296
rect 5675 242 5731 244
rect 6123 514 6179 516
rect 6123 462 6125 514
rect 6125 462 6177 514
rect 6177 462 6179 514
rect 6123 460 6179 462
rect 6123 296 6179 298
rect 6123 244 6125 296
rect 6125 244 6177 296
rect 6177 244 6179 296
rect 6123 242 6179 244
rect 6571 514 6627 516
rect 6571 462 6573 514
rect 6573 462 6625 514
rect 6625 462 6627 514
rect 6571 460 6627 462
rect 6571 296 6627 298
rect 6571 244 6573 296
rect 6573 244 6625 296
rect 6625 244 6627 296
rect 6571 242 6627 244
rect 7048 508 7208 510
rect 7048 248 7050 508
rect 7050 248 7206 508
rect 7206 248 7208 508
rect 7048 246 7208 248
<< metal3 >>
rect 91 3545 7407 3555
rect 91 3281 172 3545
rect 228 3281 620 3545
rect 676 3281 1301 3545
rect 1565 3281 1943 3545
rect 1999 3281 2391 3545
rect 2447 3281 2839 3545
rect 2895 3281 3287 3545
rect 3343 3281 3735 3545
rect 3791 3281 4183 3545
rect 4239 3281 4386 3545
rect 4442 3281 4589 3545
rect 4645 3281 5037 3545
rect 5093 3281 5485 3545
rect 5541 3281 5933 3545
rect 5989 3281 6381 3545
rect 6437 3281 6829 3545
rect 6885 3281 7048 3545
rect 7208 3281 7407 3545
rect 91 3271 7407 3281
rect 2004 3042 2392 3058
rect 2004 2986 2014 3042
rect 2382 2986 2392 3042
rect 2004 2970 2392 2986
rect 91 2269 7407 2279
rect 91 2005 172 2269
rect 228 2005 620 2269
rect 676 2005 1068 2269
rect 1124 2005 1516 2269
rect 1572 2005 1720 2269
rect 1776 2005 1943 2269
rect 1999 2005 2391 2269
rect 2447 2005 2839 2269
rect 2895 2005 3287 2269
rect 3343 2005 3735 2269
rect 3791 2005 4183 2269
rect 4239 2005 4386 2269
rect 4442 2005 4589 2269
rect 4645 2005 5037 2269
rect 5093 2005 5485 2269
rect 5541 2005 5933 2269
rect 5989 2005 6381 2269
rect 6437 2005 6829 2269
rect 6885 2005 7042 2269
rect 7202 2005 7407 2269
rect 91 1995 7407 2005
rect 1262 1489 4770 1505
rect 1262 1433 1272 1489
rect 1432 1433 4600 1489
rect 4760 1433 4770 1489
rect 1262 1417 4770 1433
rect 91 1221 7407 1298
rect 91 1218 3213 1221
rect 91 1162 128 1218
rect 184 1207 3213 1218
rect 184 1162 653 1207
rect 91 1151 653 1162
rect 709 1151 1101 1207
rect 1157 1151 2517 1207
rect 2573 1151 2965 1207
rect 3021 1151 3213 1207
rect 91 1000 3213 1151
rect 91 944 128 1000
rect 184 989 3213 1000
rect 184 944 653 989
rect 91 933 653 944
rect 709 933 1101 989
rect 1157 933 2517 989
rect 2573 933 2965 989
rect 3021 957 3213 989
rect 3269 957 3661 1221
rect 3717 1218 7407 1221
rect 3717 1216 7096 1218
rect 3717 1207 5227 1216
rect 3717 1151 4986 1207
rect 5042 1160 5227 1207
rect 5283 1160 5675 1216
rect 5731 1160 6123 1216
rect 6179 1160 6571 1216
rect 6627 1162 7096 1216
rect 7152 1162 7407 1218
rect 6627 1160 7407 1162
rect 5042 1151 7407 1160
rect 3717 1000 7407 1151
rect 3717 998 7096 1000
rect 3717 989 5227 998
rect 3717 957 4986 989
rect 3021 933 4986 957
rect 5042 942 5227 989
rect 5283 942 5675 998
rect 5731 942 6123 998
rect 6179 942 6571 998
rect 6627 944 7096 998
rect 7152 944 7407 1000
rect 6627 942 7407 944
rect 5042 933 7407 942
rect 91 843 7407 933
rect 91 554 221 555
rect 616 554 746 555
rect 5190 554 5320 555
rect 5638 554 5768 555
rect 6086 554 6216 555
rect 6534 554 6664 555
rect 91 516 7407 554
rect 91 460 128 516
rect 184 460 653 516
rect 709 515 5227 516
rect 709 460 1101 515
rect 91 459 1101 460
rect 1157 459 2517 515
rect 2573 459 2965 515
rect 3021 492 4986 515
rect 3021 459 3213 492
rect 91 329 3213 459
rect 91 298 1101 329
rect 91 242 128 298
rect 184 242 653 298
rect 709 273 1101 298
rect 1157 273 2517 329
rect 2573 273 2965 329
rect 3021 273 3213 329
rect 709 242 3213 273
rect 91 228 3213 242
rect 3269 228 3661 492
rect 3717 459 4986 492
rect 5042 460 5227 515
rect 5283 460 5675 516
rect 5731 460 6123 516
rect 6179 460 6571 516
rect 6627 510 7407 516
rect 6627 460 7048 510
rect 5042 459 7048 460
rect 3717 329 7048 459
rect 3717 273 4986 329
rect 5042 298 7048 329
rect 5042 273 5227 298
rect 3717 242 5227 273
rect 5283 242 5675 298
rect 5731 242 6123 298
rect 6179 242 6571 298
rect 6627 246 7048 298
rect 7208 246 7407 510
rect 6627 242 7407 246
rect 3717 228 7407 242
rect 91 203 7407 228
rect 632 56 972 95
rect 632 0 668 56
rect 724 0 880 56
rect 936 0 972 56
rect 632 -38 972 0
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_0
timestamp 1749760379
transform 1 0 1748 0 1 2132
box 0 0 1 1
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_1
timestamp 1749760379
transform 1 0 4414 0 1 2132
box 0 0 1 1
use M1_NACTIVE4310591302070_512x8m81  M1_NACTIVE4310591302070_512x8m81_0
timestamp 1749760379
transform 1 0 7121 0 1 2132
box 0 0 1 1
use M1_NACTIVE_01_512x8m81  M1_NACTIVE_01_512x8m81_0
timestamp 1749760379
transform 1 0 7124 0 1 1081
box 0 0 1 1
use M1_NACTIVE_01_512x8m81  M1_NACTIVE_01_512x8m81_1
timestamp 1749760379
transform 1 0 156 0 1 379
box 0 0 1 1
use M1_NACTIVE_01_512x8m81  M1_NACTIVE_01_512x8m81_2
timestamp 1749760379
transform 1 0 156 0 1 1081
box 0 0 1 1
use M1_PACTIVE4310591302039_512x8m81  M1_PACTIVE4310591302039_512x8m81_0
timestamp 1749760379
transform 1 0 4414 0 1 3408
box 0 0 1 1
use M1_PACTIVE4310591302069_512x8m81  M1_PACTIVE4310591302069_512x8m81_0
timestamp 1749760379
transform 1 0 7121 0 1 373
box 0 0 1 1
use M1_PACTIVE4310591302069_512x8m81  M1_PACTIVE4310591302069_512x8m81_1
timestamp 1749760379
transform 1 0 7121 0 1 3408
box 0 0 1 1
use M1_PACTIVE4310591302071_512x8m81  M1_PACTIVE4310591302071_512x8m81_0
timestamp 1749760379
transform 1 0 1427 0 1 3408
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_0
timestamp 1749760379
transform 1 0 4039 0 1 -41
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_1
timestamp 1749760379
transform 1 0 4337 0 1 1407
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_2
timestamp 1749760379
transform 1 0 5243 0 1 709
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_3
timestamp 1749760379
transform 1 0 5477 0 1 1656
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_4
timestamp 1749760379
transform 1 0 4649 0 1 41
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_5
timestamp 1749760379
transform 1 0 4678 0 1 1457
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_6
timestamp 1749760379
transform 1 0 5919 0 1 1656
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_7
timestamp 1749760379
transform 1 0 6373 0 1 1656
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_8
timestamp 1749760379
transform 1 0 6716 0 1 1656
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_9
timestamp 1749760379
transform 0 -1 1406 1 0 694
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_10
timestamp 1749760379
transform 1 0 822 0 1 61
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_11
timestamp 1749760379
transform 1 0 1100 0 1 635
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_12
timestamp 1749760379
transform 1 0 2579 0 1 711
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_13
timestamp 1749760379
transform 1 0 2528 0 1 47
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_14
timestamp 1749760379
transform 1 0 3382 0 1 47
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_15
timestamp 1749760379
transform 1 0 1777 0 1 -224
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_16
timestamp 1749760379
transform 1 0 540 0 1 1663
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_17
timestamp 1749760379
transform 1 0 540 0 1 1406
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_18
timestamp 1749760379
transform 1 0 1696 0 1 2847
box 0 0 1 1
use M2_M1$$201262124_512x8m81  M2_M1$$201262124_512x8m81_0
timestamp 1749760379
transform 1 0 802 0 1 29
box 0 0 1 1
use M2_M1$$202395692_512x8m81  M2_M1$$202395692_512x8m81_0
timestamp 1749760379
transform 1 0 5014 0 1 394
box 0 0 1 1
use M2_M1$$202395692_512x8m81  M2_M1$$202395692_512x8m81_1
timestamp 1749760379
transform 1 0 1129 0 1 394
box 0 0 1 1
use M2_M1$$202395692_512x8m81  M2_M1$$202395692_512x8m81_2
timestamp 1749760379
transform 1 0 2545 0 1 394
box 0 0 1 1
use M2_M1$$202395692_512x8m81  M2_M1$$202395692_512x8m81_3
timestamp 1749760379
transform 1 0 2993 0 1 394
box 0 0 1 1
use M2_M1$$202396716_512x8m81  M2_M1$$202396716_512x8m81_0
timestamp 1749760379
transform 1 0 1636 0 1 703
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_0
timestamp 1749760379
transform 1 0 5255 0 -1 1079
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_1
timestamp 1749760379
transform 1 0 4121 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_2
timestamp 1749760379
transform 1 0 7124 0 1 1081
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_3
timestamp 1749760379
transform 1 0 6599 0 1 379
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_4
timestamp 1749760379
transform 1 0 6151 0 1 379
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_5
timestamp 1749760379
transform 1 0 5703 0 1 379
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_6
timestamp 1749760379
transform 1 0 5255 0 1 379
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_7
timestamp 1749760379
transform 1 0 5014 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_8
timestamp 1749760379
transform 1 0 4790 0 1 336
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_9
timestamp 1749760379
transform 1 0 4790 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_10
timestamp 1749760379
transform 1 0 4121 0 1 336
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_11
timestamp 1749760379
transform 1 0 5703 0 -1 1079
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_12
timestamp 1749760379
transform 1 0 6151 0 -1 1079
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_13
timestamp 1749760379
transform 1 0 6599 0 -1 1079
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_14
timestamp 1749760379
transform 1 0 2545 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_15
timestamp 1749760379
transform 1 0 2993 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_16
timestamp 1749760379
transform 1 0 156 0 1 1081
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_17
timestamp 1749760379
transform 1 0 156 0 1 379
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_18
timestamp 1749760379
transform 1 0 681 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_19
timestamp 1749760379
transform 1 0 681 0 1 379
box 0 0 1 1
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_20
timestamp 1749760379
transform 1 0 1129 0 1 1070
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1749760379
transform 0 -1 4680 1 0 1461
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_1
timestamp 1749760379
transform 0 -1 456 1 0 -123
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_2
timestamp 1749760379
transform 0 -1 1352 1 0 1461
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_0
timestamp 1749760379
transform 1 0 3689 0 1 1089
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_1
timestamp 1749760379
transform 1 0 3689 0 1 360
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_2
timestamp 1749760379
transform 1 0 3241 0 1 1089
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_3
timestamp 1749760379
transform 1 0 3241 0 1 360
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_4
timestamp 1749760379
transform 1 0 3315 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_5
timestamp 1749760379
transform 1 0 1971 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_6
timestamp 1749760379
transform 1 0 2419 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_7
timestamp 1749760379
transform 1 0 2867 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_8
timestamp 1749760379
transform 1 0 3315 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_9
timestamp 1749760379
transform 1 0 1748 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_10
timestamp 1749760379
transform 1 0 200 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_11
timestamp 1749760379
transform 1 0 648 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_12
timestamp 1749760379
transform 1 0 648 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_13
timestamp 1749760379
transform 1 0 200 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_14
timestamp 1749760379
transform 1 0 1544 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_15
timestamp 1749760379
transform 1 0 1096 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_16
timestamp 1749760379
transform 1 0 2867 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_17
timestamp 1749760379
transform 1 0 2419 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_18
timestamp 1749760379
transform 1 0 1971 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_19
timestamp 1749760379
transform 1 0 6409 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_20
timestamp 1749760379
transform 1 0 4414 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_21
timestamp 1749760379
transform 1 0 4414 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_22
timestamp 1749760379
transform 1 0 4211 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_23
timestamp 1749760379
transform 1 0 3763 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_24
timestamp 1749760379
transform 1 0 4211 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_25
timestamp 1749760379
transform 1 0 3763 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_26
timestamp 1749760379
transform 1 0 5513 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_27
timestamp 1749760379
transform 1 0 5065 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_28
timestamp 1749760379
transform 1 0 4617 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_29
timestamp 1749760379
transform 1 0 5961 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_30
timestamp 1749760379
transform 1 0 6857 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_31
timestamp 1749760379
transform 1 0 6409 0 1 2137
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_32
timestamp 1749760379
transform 1 0 4617 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_33
timestamp 1749760379
transform 1 0 5065 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_34
timestamp 1749760379
transform 1 0 5513 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_35
timestamp 1749760379
transform 1 0 5961 0 1 3413
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_36
timestamp 1749760379
transform 1 0 6857 0 1 3413
box 0 0 1 1
use M2_M14310591302025_512x8m81  M2_M14310591302025_512x8m81_0
timestamp 1749760379
transform 0 -1 2198 1 0 3014
box 0 0 1 1
use M2_M14310591302073_512x8m81  M2_M14310591302073_512x8m81_0
timestamp 1749760379
transform 1 0 7128 0 1 378
box 0 0 1 1
use M2_M14310591302073_512x8m81  M2_M14310591302073_512x8m81_1
timestamp 1749760379
transform 1 0 7128 0 1 3413
box 0 0 1 1
use M2_M14310591302073_512x8m81  M2_M14310591302073_512x8m81_2
timestamp 1749760379
transform 1 0 7122 0 1 2137
box 0 0 1 1
use M2_M14310591302074_512x8m81  M2_M14310591302074_512x8m81_0
timestamp 1749760379
transform 1 0 1433 0 1 3413
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_0
timestamp 1749760379
transform 1 0 5255 0 -1 1079
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_1
timestamp 1749760379
transform 1 0 6599 0 1 379
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_2
timestamp 1749760379
transform 1 0 7124 0 1 1081
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_3
timestamp 1749760379
transform 1 0 5255 0 1 379
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_4
timestamp 1749760379
transform 1 0 5703 0 1 379
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_5
timestamp 1749760379
transform 1 0 6151 0 1 379
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_6
timestamp 1749760379
transform 1 0 5014 0 1 1070
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_7
timestamp 1749760379
transform 1 0 5703 0 -1 1079
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_8
timestamp 1749760379
transform 1 0 6599 0 -1 1079
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_9
timestamp 1749760379
transform 1 0 6151 0 -1 1079
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_10
timestamp 1749760379
transform 1 0 2545 0 1 1070
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_11
timestamp 1749760379
transform 1 0 2993 0 1 1070
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_12
timestamp 1749760379
transform 1 0 156 0 1 1081
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_13
timestamp 1749760379
transform 1 0 156 0 1 379
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_14
timestamp 1749760379
transform 1 0 681 0 1 1070
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_15
timestamp 1749760379
transform 1 0 681 0 1 379
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_16
timestamp 1749760379
transform 1 0 1129 0 1 1070
box 0 0 1 1
use M3_M2$$201255980_512x8m81  M3_M2$$201255980_512x8m81_0
timestamp 1749760379
transform 1 0 802 0 1 28
box 0 0 1 1
use M3_M2$$202397740_512x8m81  M3_M2$$202397740_512x8m81_0
timestamp 1749760379
transform 1 0 5014 0 1 394
box 0 0 1 1
use M3_M2$$202397740_512x8m81  M3_M2$$202397740_512x8m81_1
timestamp 1749760379
transform 1 0 2545 0 1 394
box 0 0 1 1
use M3_M2$$202397740_512x8m81  M3_M2$$202397740_512x8m81_2
timestamp 1749760379
transform 1 0 2993 0 1 394
box 0 0 1 1
use M3_M2$$202397740_512x8m81  M3_M2$$202397740_512x8m81_3
timestamp 1749760379
transform 1 0 1129 0 1 394
box 0 0 1 1
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_0
timestamp 1749760379
transform 1 0 4680 0 1 1461
box 0 0 1 1
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_1
timestamp 1749760379
transform 1 0 1352 0 1 1461
box 0 0 1 1
use M3_M24310591302026_512x8m81  M3_M24310591302026_512x8m81_0
timestamp 1749760379
transform 0 -1 2198 1 0 3014
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_0
timestamp 1749760379
transform 1 0 3689 0 1 1089
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_1
timestamp 1749760379
transform 1 0 3689 0 1 360
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_2
timestamp 1749760379
transform 1 0 3241 0 1 1089
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_3
timestamp 1749760379
transform 1 0 3241 0 1 360
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_4
timestamp 1749760379
transform 1 0 1544 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_5
timestamp 1749760379
transform 1 0 1096 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_6
timestamp 1749760379
transform 1 0 1748 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_7
timestamp 1749760379
transform 1 0 648 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_8
timestamp 1749760379
transform 1 0 1971 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_9
timestamp 1749760379
transform 1 0 2419 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_10
timestamp 1749760379
transform 1 0 2867 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_11
timestamp 1749760379
transform 1 0 3315 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_12
timestamp 1749760379
transform 1 0 200 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_13
timestamp 1749760379
transform 1 0 200 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_14
timestamp 1749760379
transform 1 0 648 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_15
timestamp 1749760379
transform 1 0 1971 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_16
timestamp 1749760379
transform 1 0 2419 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_17
timestamp 1749760379
transform 1 0 2867 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_18
timestamp 1749760379
transform 1 0 3315 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_19
timestamp 1749760379
transform 1 0 4211 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_20
timestamp 1749760379
transform 1 0 3763 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_21
timestamp 1749760379
transform 1 0 4617 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_22
timestamp 1749760379
transform 1 0 5065 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_23
timestamp 1749760379
transform 1 0 5513 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_24
timestamp 1749760379
transform 1 0 5961 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_25
timestamp 1749760379
transform 1 0 6857 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_26
timestamp 1749760379
transform 1 0 6409 0 1 3413
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_27
timestamp 1749760379
transform 1 0 4211 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_28
timestamp 1749760379
transform 1 0 3763 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_29
timestamp 1749760379
transform 1 0 4617 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_30
timestamp 1749760379
transform 1 0 5065 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_31
timestamp 1749760379
transform 1 0 5513 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_32
timestamp 1749760379
transform 1 0 5961 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_33
timestamp 1749760379
transform 1 0 6857 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_34
timestamp 1749760379
transform 1 0 6409 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_35
timestamp 1749760379
transform 1 0 4414 0 1 2137
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_36
timestamp 1749760379
transform 1 0 4414 0 1 3413
box 0 0 1 1
use M3_M24310591302050_512x8m81  M3_M24310591302050_512x8m81_0
timestamp 1749760379
transform 1 0 1433 0 1 3413
box 0 0 1 1
use M3_M24310591302072_512x8m81  M3_M24310591302072_512x8m81_0
timestamp 1749760379
transform 1 0 7128 0 1 378
box 0 0 1 1
use M3_M24310591302072_512x8m81  M3_M24310591302072_512x8m81_1
timestamp 1749760379
transform 1 0 7128 0 1 3413
box 0 0 1 1
use M3_M24310591302072_512x8m81  M3_M24310591302072_512x8m81_2
timestamp 1749760379
transform 1 0 7122 0 1 2137
box 0 0 1 1
use nmos_1p2$$202595372_512x8m81  nmos_1p2$$202595372_512x8m81_0
timestamp 1749760379
transform 1 0 2853 0 1 372
box -31 0 -30 1
use nmos_1p2$$202595372_512x8m81  nmos_1p2$$202595372_512x8m81_1
timestamp 1749760379
transform 1 0 2181 0 1 372
box -31 0 -30 1
use nmos_1p2$$202596396_512x8m81  nmos_1p2$$202596396_512x8m81_0
timestamp 1749760379
transform 1 0 2405 0 1 372
box -31 0 -30 1
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_0
timestamp 1749760379
transform 1 0 4842 0 -1 440
box 0 0 1 1
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_1
timestamp 1749760379
transform 1 0 4618 0 -1 440
box 0 0 1 1
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_2
timestamp 1749760379
transform 1 0 509 0 1 213
box 0 0 1 1
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_3
timestamp 1749760379
transform 1 0 733 0 1 213
box 0 0 1 1
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_4
timestamp 1749760379
transform 1 0 1181 0 1 295
box 0 0 1 1
use nmos_5p04310591302010_512x8m81  nmos_5p04310591302010_512x8m81_0
timestamp 1749760379
transform 1 0 1688 0 1 109
box 0 0 1 1
use nmos_5p04310591302039_512x8m81  nmos_5p04310591302039_512x8m81_0
timestamp 1749760379
transform 1 0 3950 0 1 109
box 0 0 1 1
use nmos_5p04310591302075_512x8m81  nmos_5p04310591302075_512x8m81_0
timestamp 1749760379
transform 1 0 4669 0 1 3214
box 0 0 1 1
use nmos_5p04310591302075_512x8m81  nmos_5p04310591302075_512x8m81_1
timestamp 1749760379
transform 1 0 2023 0 1 3214
box 0 0 1 1
use nmos_5p04310591302076_512x8m81  nmos_5p04310591302076_512x8m81_0
timestamp 1749760379
transform 1 0 3293 0 1 324
box 0 0 1 1
use nmos_5p04310591302078_512x8m81  nmos_5p04310591302078_512x8m81_0
timestamp 1749760379
transform 1 0 252 0 1 3214
box 0 0 1 1
use nmos_5p04310591302081_512x8m81  nmos_5p04310591302081_512x8m81_0
timestamp 1749760379
transform 1 0 5307 0 1 381
box 0 0 1 1
use pmos_1p2$$202586156_512x8m81  pmos_1p2$$202586156_512x8m81_0
timestamp 1749760379
transform 1 0 2405 0 1 843
box -31 0 -30 1
use pmos_1p2$$202587180_512x8m81  pmos_1p2$$202587180_512x8m81_0
timestamp 1749760379
transform 1 0 1719 0 1 843
box -31 0 -30 1
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_0
timestamp 1749760379
transform 1 0 4842 0 -1 1297
box 0 0 1 1
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_1
timestamp 1749760379
transform 1 0 733 0 1 843
box 0 0 1 1
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_2
timestamp 1749760379
transform 1 0 2822 0 1 843
box 0 0 1 1
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_3
timestamp 1749760379
transform 1 0 509 0 1 843
box 0 0 1 1
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_4
timestamp 1749760379
transform 1 0 1181 0 1 843
box 0 0 1 1
use pmos_5p04310591302020_512x8m81  pmos_5p04310591302020_512x8m81_0
timestamp 1749760379
transform 1 0 3950 0 1 843
box 0 0 1 1
use pmos_5p04310591302041_512x8m81  pmos_5p04310591302041_512x8m81_0
timestamp 1749760379
transform 1 0 4510 0 -1 1297
box 0 0 1 1
use pmos_5p04310591302041_512x8m81  pmos_5p04310591302041_512x8m81_1
timestamp 1749760379
transform 1 0 2036 0 1 843
box 0 0 1 1
use pmos_5p04310591302077_512x8m81  pmos_5p04310591302077_512x8m81_0
timestamp 1749760379
transform 1 0 4669 0 1 1884
box 0 0 1 1
use pmos_5p04310591302077_512x8m81  pmos_5p04310591302077_512x8m81_1
timestamp 1749760379
transform 1 0 2023 0 1 1884
box 0 0 1 1
use pmos_5p04310591302079_512x8m81  pmos_5p04310591302079_512x8m81_0
timestamp 1749760379
transform 1 0 5307 0 1 843
box 0 0 1 1
use pmos_5p04310591302080_512x8m81  pmos_5p04310591302080_512x8m81_0
timestamp 1749760379
transform 1 0 3293 0 1 843
box 0 0 1 1
use pmos_5p04310591302082_512x8m81  pmos_5p04310591302082_512x8m81_0
timestamp 1749760379
transform 1 0 252 0 1 1884
box 0 0 1 1
<< labels >>
rlabel metal3 s 252 3479 252 3479 4 vss
port 1 nsew
flabel metal3 s 2197 3015 2197 3015 0 FreeSans 1000 0 0 0 IGWEN
port 2 nsew
rlabel metal3 s 252 2175 252 2175 4 vdd
port 3 nsew
rlabel metal3 s 252 379 252 379 4 vss
port 1 nsew
rlabel metal3 s 252 1070 252 1070 4 vdd
port 3 nsew
rlabel metal3 s 865 61 865 61 4 clk
port 4 nsew
rlabel metal1 s 481 1428 481 1428 4 wen
port 5 nsew
rlabel metal1 s 6626 3004 6626 3004 4 GWE
port 6 nsew
<< properties >>
string GDS_END 992554
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 969586
string path 6.310 7.305 23.850 7.305 
<< end >>
