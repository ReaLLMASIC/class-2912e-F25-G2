magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< metal3 >>
rect 430 28230 21970 28590
rect 430 27210 21970 27570
rect 430 26430 21970 26790
rect 430 25410 21970 25770
rect 430 24630 21970 24990
rect 430 23610 21970 23970
rect 430 22830 21970 23190
rect 430 21810 21970 22170
rect 430 21030 21970 21390
rect 430 20010 21970 20370
rect 430 19230 21970 19590
rect 430 18210 21970 18570
rect 430 17430 21970 17790
rect 430 16410 21970 16770
rect 430 15630 21970 15990
rect 430 14610 21970 14970
rect 430 13830 21970 14190
rect 430 12810 21970 13170
rect 430 12030 21970 12390
rect 430 11010 21970 11370
rect 430 10230 21970 10590
rect 430 9210 21970 9570
rect 430 8430 21970 8790
rect 430 7410 21970 7770
rect 430 6630 21970 6990
rect 430 5610 21970 5970
rect 430 4830 21970 5190
rect 430 3810 21970 4170
rect 430 3030 21970 3390
rect 430 2010 21970 2370
rect 430 1230 21970 1590
rect 430 210 21970 570
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_0
timestamp 1749760379
transform -1 0 16800 0 1 2700
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_1
timestamp 1749760379
transform -1 0 16800 0 1 4500
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_2
timestamp 1749760379
transform -1 0 16800 0 1 6300
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_3
timestamp 1749760379
transform -1 0 16800 0 1 8100
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_4
timestamp 1749760379
transform -1 0 16800 0 1 9900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_5
timestamp 1749760379
transform -1 0 16800 0 1 11700
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_6
timestamp 1749760379
transform -1 0 16800 0 1 900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_7
timestamp 1749760379
transform -1 0 6000 0 1 2700
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_8
timestamp 1749760379
transform -1 0 6000 0 1 4500
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_9
timestamp 1749760379
transform -1 0 6000 0 1 6300
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_10
timestamp 1749760379
transform -1 0 6000 0 1 11700
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_11
timestamp 1749760379
transform -1 0 6000 0 1 9900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_12
timestamp 1749760379
transform -1 0 6000 0 1 8100
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_13
timestamp 1749760379
transform -1 0 6000 0 1 900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_14
timestamp 1749760379
transform -1 0 6000 0 1 26100
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_15
timestamp 1749760379
transform -1 0 6000 0 1 27900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_16
timestamp 1749760379
transform -1 0 6000 0 1 18900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_17
timestamp 1749760379
transform -1 0 6000 0 1 17100
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_18
timestamp 1749760379
transform -1 0 6000 0 1 22500
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_19
timestamp 1749760379
transform -1 0 6000 0 1 20700
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_20
timestamp 1749760379
transform -1 0 6000 0 1 24300
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_21
timestamp 1749760379
transform -1 0 16800 0 1 17100
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_22
timestamp 1749760379
transform -1 0 16800 0 1 18900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_23
timestamp 1749760379
transform -1 0 16800 0 1 20700
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_24
timestamp 1749760379
transform -1 0 16800 0 1 22500
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_25
timestamp 1749760379
transform -1 0 16800 0 1 24300
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_26
timestamp 1749760379
transform -1 0 16800 0 1 26100
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_27
timestamp 1749760379
transform -1 0 16800 0 1 27900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_28
timestamp 1749760379
transform -1 0 6000 0 1 13500
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_29
timestamp 1749760379
transform -1 0 6000 0 1 15300
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_30
timestamp 1749760379
transform -1 0 11400 0 1 4500
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_31
timestamp 1749760379
transform -1 0 11400 0 1 6300
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_32
timestamp 1749760379
transform -1 0 11400 0 1 8100
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_33
timestamp 1749760379
transform -1 0 11400 0 1 9900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_34
timestamp 1749760379
transform -1 0 11400 0 1 11700
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_35
timestamp 1749760379
transform -1 0 11400 0 1 13500
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_36
timestamp 1749760379
transform -1 0 11400 0 1 15300
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_37
timestamp 1749760379
transform -1 0 11400 0 1 17100
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_38
timestamp 1749760379
transform -1 0 11400 0 1 18900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_39
timestamp 1749760379
transform -1 0 11400 0 1 20700
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_40
timestamp 1749760379
transform -1 0 11400 0 1 22500
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_41
timestamp 1749760379
transform -1 0 11400 0 1 24300
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_42
timestamp 1749760379
transform -1 0 11400 0 1 26100
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_43
timestamp 1749760379
transform -1 0 11400 0 1 27900
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_44
timestamp 1749760379
transform -1 0 11400 0 1 2700
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_45
timestamp 1749760379
transform -1 0 16800 0 1 13500
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_46
timestamp 1749760379
transform -1 0 16800 0 1 15300
box -68 -968 668 968
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_47
timestamp 1749760379
transform -1 0 11400 0 1 900
box -68 -968 668 968
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_0
timestamp 1749760379
transform -1 0 18000 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_1
timestamp 1749760379
transform -1 0 18600 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_2
timestamp 1749760379
transform -1 0 19200 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_3
timestamp 1749760379
transform -1 0 19800 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_4
timestamp 1749760379
transform -1 0 20400 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_5
timestamp 1749760379
transform -1 0 21000 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_6
timestamp 1749760379
transform -1 0 21600 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_7
timestamp 1749760379
transform -1 0 6600 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_8
timestamp 1749760379
transform -1 0 7200 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_9
timestamp 1749760379
transform -1 0 7800 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_10
timestamp 1749760379
transform -1 0 8400 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_11
timestamp 1749760379
transform -1 0 9000 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_12
timestamp 1749760379
transform -1 0 9600 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_13
timestamp 1749760379
transform -1 0 10200 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_14
timestamp 1749760379
transform -1 0 10800 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_15
timestamp 1749760379
transform -1 0 17400 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_16
timestamp 1749760379
transform 1 0 12600 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_17
timestamp 1749760379
transform 1 0 12000 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_18
timestamp 1749760379
transform 1 0 11400 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_19
timestamp 1749760379
transform 1 0 13800 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_20
timestamp 1749760379
transform 1 0 600 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_21
timestamp 1749760379
transform 1 0 1200 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_22
timestamp 1749760379
transform 1 0 1800 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_23
timestamp 1749760379
transform 1 0 2400 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_24
timestamp 1749760379
transform 1 0 3000 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_25
timestamp 1749760379
transform 1 0 3600 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_26
timestamp 1749760379
transform 1 0 4200 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_27
timestamp 1749760379
transform 1 0 4800 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_28
timestamp 1749760379
transform 1 0 14400 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_29
timestamp 1749760379
transform 1 0 15000 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_30
timestamp 1749760379
transform 1 0 15600 0 1 0
box -68 -68 668 28868
use Cell_array32x1_256x8m81  Cell_array32x1_256x8m81_31
timestamp 1749760379
transform 1 0 13200 0 1 0
box -68 -68 668 28868
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_0
timestamp 1749760379
transform 1 0 21600 0 1 1780
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_1
timestamp 1749760379
transform 1 0 21600 0 1 3580
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_2
timestamp 1749760379
transform 1 0 21600 0 1 5380
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_3
timestamp 1749760379
transform 1 0 21600 0 1 7180
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_4
timestamp 1749760379
transform 1 0 21600 0 1 8980
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_5
timestamp 1749760379
transform 1 0 21600 0 1 -20
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_6
timestamp 1749760379
transform 1 0 21600 0 1 10780
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_7
timestamp 1749760379
transform 1 0 21600 0 1 23380
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_8
timestamp 1749760379
transform 1 0 21600 0 1 21580
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_9
timestamp 1749760379
transform 1 0 21600 0 1 19780
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_10
timestamp 1749760379
transform 1 0 21600 0 1 17980
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_11
timestamp 1749760379
transform 1 0 21600 0 1 16180
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_12
timestamp 1749760379
transform 1 0 21600 0 1 25180
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_13
timestamp 1749760379
transform 1 0 21600 0 1 26980
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_14
timestamp 1749760379
transform 1 0 21600 0 1 12580
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_15
timestamp 1749760379
transform 1 0 21600 0 1 14380
box -68 -48 668 1888
<< labels >>
rlabel metal3 20377 26560 20377 26560 4 WL[29]
rlabel metal3 20377 25660 20377 25660 4 WL[28]
rlabel metal3 21577 25660 21577 25660 4 WL[28]
rlabel metal3 21577 26560 21577 26560 4 WL[29]
rlabel metal3 21577 27460 21577 27460 4 WL[30]
rlabel metal3 21577 28360 21577 28360 4 WL[31]
rlabel metal3 20377 27460 20377 27460 4 WL[30]
rlabel metal3 20377 28360 20377 28360 4 WL[31]
rlabel metal3 21519 28360 21519 28360 4 WL[31]
rlabel metal3 21519 25660 21519 25660 4 WL[28]
rlabel metal3 21519 26560 21519 26560 4 WL[29]
rlabel metal3 21519 27460 21519 27460 4 WL[30]
rlabel metal3 19279 25660 19279 25660 4 WL[28]
rlabel metal3 19279 26560 19279 26560 4 WL[29]
rlabel metal3 19279 27460 19279 27460 4 WL[30]
rlabel metal3 19279 28360 19279 28360 4 WL[31]
rlabel metal3 20479 25660 20479 25660 4 WL[28]
rlabel metal3 20479 26560 20479 26560 4 WL[29]
rlabel metal3 20479 27460 20479 27460 4 WL[30]
rlabel metal3 20479 28360 20479 28360 4 WL[31]
rlabel metal3 20977 28360 20977 28360 4 WL[31]
rlabel metal3 20977 27460 20977 27460 4 WL[30]
rlabel metal3 20977 26560 20977 26560 4 WL[29]
rlabel metal3 20977 25660 20977 25660 4 WL[28]
rlabel metal3 19777 26560 19777 26560 4 WL[29]
rlabel metal3 19777 25660 19777 25660 4 WL[28]
rlabel metal3 19777 28360 19777 28360 4 WL[31]
rlabel metal3 19777 27460 19777 27460 4 WL[30]
rlabel metal3 19177 25660 19177 25660 4 WL[28]
rlabel metal3 19177 28360 19177 28360 4 WL[31]
rlabel metal3 19177 27460 19177 27460 4 WL[30]
rlabel metal3 19177 26560 19177 26560 4 WL[29]
rlabel metal3 17977 28360 17977 28360 4 WL[31]
rlabel metal3 17977 27460 17977 27460 4 WL[30]
rlabel metal3 17977 26560 17977 26560 4 WL[29]
rlabel metal3 17977 25660 17977 25660 4 WL[28]
rlabel metal3 16879 25660 16879 25660 4 WL[28]
rlabel metal3 16879 26560 16879 26560 4 WL[29]
rlabel metal3 16879 27460 16879 27460 4 WL[30]
rlabel metal3 16879 28360 16879 28360 4 WL[31]
rlabel metal3 18079 25660 18079 25660 4 WL[28]
rlabel metal3 18079 26560 18079 26560 4 WL[29]
rlabel metal3 18079 27460 18079 27460 4 WL[30]
rlabel metal3 18079 28360 18079 28360 4 WL[31]
rlabel metal3 17377 26560 17377 26560 4 WL[29]
rlabel metal3 17377 25660 17377 25660 4 WL[28]
rlabel metal3 17377 28360 17377 28360 4 WL[31]
rlabel metal3 17377 27460 17377 27460 4 WL[30]
rlabel metal3 18577 28360 18577 28360 4 WL[31]
rlabel metal3 18577 27460 18577 27460 4 WL[30]
rlabel metal3 18577 26560 18577 26560 4 WL[29]
rlabel metal3 18577 25660 18577 25660 4 WL[28]
rlabel metal3 17977 24760 17977 24760 4 WL[27]
rlabel metal3 17977 23860 17977 23860 4 WL[26]
rlabel metal3 16879 22060 16879 22060 4 WL[24]
rlabel metal3 16879 22960 16879 22960 4 WL[25]
rlabel metal3 18079 23860 18079 23860 4 WL[26]
rlabel metal3 18079 24760 18079 24760 4 WL[27]
rlabel metal3 16879 23860 16879 23860 4 WL[26]
rlabel metal3 16879 24760 16879 24760 4 WL[27]
rlabel metal3 17377 24760 17377 24760 4 WL[27]
rlabel metal3 17377 23860 17377 23860 4 WL[26]
rlabel metal3 18079 22060 18079 22060 4 WL[24]
rlabel metal3 18079 22960 18079 22960 4 WL[25]
rlabel metal3 18577 24760 18577 24760 4 WL[27]
rlabel metal3 18577 23860 18577 23860 4 WL[26]
rlabel metal3 18577 22960 18577 22960 4 WL[25]
rlabel metal3 18577 22060 18577 22060 4 WL[24]
rlabel metal3 17977 22960 17977 22960 4 WL[25]
rlabel metal3 17977 22060 17977 22060 4 WL[24]
rlabel metal3 17377 22960 17377 22960 4 WL[25]
rlabel metal3 17377 22060 17377 22060 4 WL[24]
rlabel metal3 21577 23860 21577 23860 4 WL[26]
rlabel metal3 21519 23860 21519 23860 4 WL[26]
rlabel metal3 21519 24760 21519 24760 4 WL[27]
rlabel metal3 21577 24760 21577 24760 4 WL[27]
rlabel metal3 20977 24760 20977 24760 4 WL[27]
rlabel metal3 20977 23860 20977 23860 4 WL[26]
rlabel metal3 20377 22960 20377 22960 4 WL[25]
rlabel metal3 20377 22060 20377 22060 4 WL[24]
rlabel metal3 21519 22960 21519 22960 4 WL[25]
rlabel metal3 20977 22960 20977 22960 4 WL[25]
rlabel metal3 19777 24760 19777 24760 4 WL[27]
rlabel metal3 19777 23860 19777 23860 4 WL[26]
rlabel metal3 19279 23860 19279 23860 4 WL[26]
rlabel metal3 19279 24760 19279 24760 4 WL[27]
rlabel metal3 20977 22060 20977 22060 4 WL[24]
rlabel metal3 19177 24760 19177 24760 4 WL[27]
rlabel metal3 19177 23860 19177 23860 4 WL[26]
rlabel metal3 21519 22060 21519 22060 4 WL[24]
rlabel metal3 19177 22960 19177 22960 4 WL[25]
rlabel metal3 19177 22060 19177 22060 4 WL[24]
rlabel metal3 19279 22060 19279 22060 4 WL[24]
rlabel metal3 19279 22960 19279 22960 4 WL[25]
rlabel metal3 20479 23860 20479 23860 4 WL[26]
rlabel metal3 20479 24760 20479 24760 4 WL[27]
rlabel metal3 19777 22960 19777 22960 4 WL[25]
rlabel metal3 19777 22060 19777 22060 4 WL[24]
rlabel metal3 20377 24760 20377 24760 4 WL[27]
rlabel metal3 20377 23860 20377 23860 4 WL[26]
rlabel metal3 20479 22060 20479 22060 4 WL[24]
rlabel metal3 20479 22960 20479 22960 4 WL[25]
rlabel metal3 21577 22960 21577 22960 4 WL[25]
rlabel metal3 21577 22060 21577 22060 4 WL[24]
rlabel metal3 13721 27460 13721 27460 4 WL[30]
rlabel metal3 13721 28360 13721 28360 4 WL[31]
rlabel metal3 13223 22060 13223 22060 4 WL[24]
rlabel metal3 13823 22060 13823 22060 4 WL[24]
rlabel metal3 13823 26560 13823 26560 4 WL[29]
rlabel metal3 12023 23860 12023 23860 4 WL[26]
rlabel metal3 14921 22060 14921 22060 4 WL[24]
rlabel metal3 14921 22960 14921 22960 4 WL[25]
rlabel metal3 13223 25660 13223 25660 4 WL[28]
rlabel metal3 13223 22960 13223 22960 4 WL[25]
rlabel metal3 12023 25660 12023 25660 4 WL[28]
rlabel metal3 12023 28360 12023 28360 4 WL[31]
rlabel metal3 12623 26560 12623 26560 4 WL[29]
rlabel metal3 12521 23860 12521 23860 4 WL[26]
rlabel metal3 12521 24760 12521 24760 4 WL[27]
rlabel metal3 13823 27460 13823 27460 4 WL[30]
rlabel metal3 12521 25660 12521 25660 4 WL[28]
rlabel metal3 12521 26560 12521 26560 4 WL[29]
rlabel metal3 14921 23860 14921 23860 4 WL[26]
rlabel metal3 14921 24760 14921 24760 4 WL[27]
rlabel metal3 14921 25660 14921 25660 4 WL[28]
rlabel metal3 14921 26560 14921 26560 4 WL[29]
rlabel metal3 14921 27460 14921 27460 4 WL[30]
rlabel metal3 14921 28360 14921 28360 4 WL[31]
rlabel metal3 13823 23860 13823 23860 4 WL[26]
rlabel metal3 15623 28360 15623 28360 4 WL[31]
rlabel metal3 15623 27460 15623 27460 4 WL[30]
rlabel metal3 15623 26560 15623 26560 4 WL[29]
rlabel metal3 15623 25660 15623 25660 4 WL[28]
rlabel metal3 15623 24760 15623 24760 4 WL[27]
rlabel metal3 15623 23860 15623 23860 4 WL[26]
rlabel metal3 15623 22960 15623 22960 4 WL[25]
rlabel metal3 15623 22060 15623 22060 4 WL[24]
rlabel metal3 15023 22960 15023 22960 4 WL[25]
rlabel metal3 15023 22060 15023 22060 4 WL[24]
rlabel metal3 14423 28360 14423 28360 4 WL[31]
rlabel metal3 14423 27460 14423 27460 4 WL[30]
rlabel metal3 14423 26560 14423 26560 4 WL[29]
rlabel metal3 14423 25660 14423 25660 4 WL[28]
rlabel metal3 14423 24760 14423 24760 4 WL[27]
rlabel metal3 14423 23860 14423 23860 4 WL[26]
rlabel metal3 12023 24760 12023 24760 4 WL[27]
rlabel metal3 13721 22060 13721 22060 4 WL[24]
rlabel metal3 13721 22960 13721 22960 4 WL[25]
rlabel metal3 13823 25660 13823 25660 4 WL[28]
rlabel metal3 14423 22960 14423 22960 4 WL[25]
rlabel metal3 13223 26560 13223 26560 4 WL[29]
rlabel metal3 13823 22960 13823 22960 4 WL[25]
rlabel metal3 12623 22960 12623 22960 4 WL[25]
rlabel metal3 13223 28360 13223 28360 4 WL[31]
rlabel metal3 12521 27460 12521 27460 4 WL[30]
rlabel metal3 12623 24760 12623 24760 4 WL[27]
rlabel metal3 12623 23860 12623 23860 4 WL[26]
rlabel metal3 13823 24760 13823 24760 4 WL[27]
rlabel metal3 12521 28360 12521 28360 4 WL[31]
rlabel metal3 12521 22060 12521 22060 4 WL[24]
rlabel metal3 12521 22960 12521 22960 4 WL[25]
rlabel metal3 14423 22060 14423 22060 4 WL[24]
rlabel metal3 16121 22060 16121 22060 4 WL[24]
rlabel metal3 16121 22960 16121 22960 4 WL[25]
rlabel metal3 12023 26560 12023 26560 4 WL[29]
rlabel metal3 13223 24760 13223 24760 4 WL[27]
rlabel metal3 15023 28360 15023 28360 4 WL[31]
rlabel metal3 12023 27460 12023 27460 4 WL[30]
rlabel metal3 15023 27460 15023 27460 4 WL[30]
rlabel metal3 12623 25660 12623 25660 4 WL[28]
rlabel metal3 13823 28360 13823 28360 4 WL[31]
rlabel metal3 15023 26560 15023 26560 4 WL[29]
rlabel metal3 15023 25660 15023 25660 4 WL[28]
rlabel metal3 13223 27460 13223 27460 4 WL[30]
rlabel metal3 15023 24760 15023 24760 4 WL[27]
rlabel metal3 15023 23860 15023 23860 4 WL[26]
rlabel metal3 13721 23860 13721 23860 4 WL[26]
rlabel metal3 16121 23860 16121 23860 4 WL[26]
rlabel metal3 16121 24760 16121 24760 4 WL[27]
rlabel metal3 16121 25660 16121 25660 4 WL[28]
rlabel metal3 12023 22060 12023 22060 4 WL[24]
rlabel metal3 12623 27460 12623 27460 4 WL[30]
rlabel metal3 16121 26560 16121 26560 4 WL[29]
rlabel metal3 16121 27460 16121 27460 4 WL[30]
rlabel metal3 12023 22960 12023 22960 4 WL[25]
rlabel metal3 12623 28360 12623 28360 4 WL[31]
rlabel metal3 16121 28360 16121 28360 4 WL[31]
rlabel metal3 13721 24760 13721 24760 4 WL[27]
rlabel metal3 12623 22060 12623 22060 4 WL[24]
rlabel metal3 13223 23860 13223 23860 4 WL[26]
rlabel metal3 13721 25660 13721 25660 4 WL[28]
rlabel metal3 13721 26560 13721 26560 4 WL[29]
rlabel metal3 13721 16660 13721 16660 4 WL[18]
rlabel metal3 13721 17560 13721 17560 4 WL[19]
rlabel metal3 12023 16660 12023 16660 4 WL[18]
rlabel metal3 14423 19360 14423 19360 4 WL[21]
rlabel metal3 12521 14860 12521 14860 4 WL[16]
rlabel metal3 15623 21160 15623 21160 4 WL[23]
rlabel metal3 15623 20260 15623 20260 4 WL[22]
rlabel metal3 15623 19360 15623 19360 4 WL[21]
rlabel metal3 15623 18460 15623 18460 4 WL[20]
rlabel metal3 15623 17560 15623 17560 4 WL[19]
rlabel metal3 15623 16660 15623 16660 4 WL[18]
rlabel metal3 15623 15760 15623 15760 4 WL[17]
rlabel metal3 15623 14860 15623 14860 4 WL[16]
rlabel metal3 13223 18460 13223 18460 4 WL[20]
rlabel metal3 13223 20260 13223 20260 4 WL[22]
rlabel metal3 15023 21160 15023 21160 4 WL[23]
rlabel metal3 15023 20260 15023 20260 4 WL[22]
rlabel metal3 15023 19360 15023 19360 4 WL[21]
rlabel metal3 15023 18460 15023 18460 4 WL[20]
rlabel metal3 15023 17560 15023 17560 4 WL[19]
rlabel metal3 15023 16660 15023 16660 4 WL[18]
rlabel metal3 15023 15760 15023 15760 4 WL[17]
rlabel metal3 15023 14860 15023 14860 4 WL[16]
rlabel metal3 12521 15760 12521 15760 4 WL[17]
rlabel metal3 14423 15760 14423 15760 4 WL[17]
rlabel metal3 13223 19360 13223 19360 4 WL[21]
rlabel metal3 13223 21160 13223 21160 4 WL[23]
rlabel metal3 13823 15760 13823 15760 4 WL[17]
rlabel metal3 12023 18460 12023 18460 4 WL[20]
rlabel metal3 12521 16660 12521 16660 4 WL[18]
rlabel metal3 12623 15760 12623 15760 4 WL[17]
rlabel metal3 12521 17560 12521 17560 4 WL[19]
rlabel metal3 12023 21160 12023 21160 4 WL[23]
rlabel metal3 12521 18460 12521 18460 4 WL[20]
rlabel metal3 12521 19360 12521 19360 4 WL[21]
rlabel metal3 12623 19360 12623 19360 4 WL[21]
rlabel metal3 12023 17560 12023 17560 4 WL[19]
rlabel metal3 12521 20260 12521 20260 4 WL[22]
rlabel metal3 13721 18460 13721 18460 4 WL[20]
rlabel metal3 13223 15760 13223 15760 4 WL[17]
rlabel metal3 12521 21160 12521 21160 4 WL[23]
rlabel metal3 13823 18460 13823 18460 4 WL[20]
rlabel metal3 13223 17560 13223 17560 4 WL[19]
rlabel metal3 13721 19360 13721 19360 4 WL[21]
rlabel metal3 13721 20260 13721 20260 4 WL[22]
rlabel metal3 14423 14860 14423 14860 4 WL[16]
rlabel metal3 14921 14860 14921 14860 4 WL[16]
rlabel metal3 14921 15760 14921 15760 4 WL[17]
rlabel metal3 14921 16660 14921 16660 4 WL[18]
rlabel metal3 13823 20260 13823 20260 4 WL[22]
rlabel metal3 14921 17560 14921 17560 4 WL[19]
rlabel metal3 12023 19360 12023 19360 4 WL[21]
rlabel metal3 14921 18460 14921 18460 4 WL[20]
rlabel metal3 14921 19360 14921 19360 4 WL[21]
rlabel metal3 12623 17560 12623 17560 4 WL[19]
rlabel metal3 13823 21160 13823 21160 4 WL[23]
rlabel metal3 14921 20260 14921 20260 4 WL[22]
rlabel metal3 14921 21160 14921 21160 4 WL[23]
rlabel metal3 12023 20260 12023 20260 4 WL[22]
rlabel metal3 12623 16660 12623 16660 4 WL[18]
rlabel metal3 14423 16660 14423 16660 4 WL[18]
rlabel metal3 12623 18460 12623 18460 4 WL[20]
rlabel metal3 13721 21160 13721 21160 4 WL[23]
rlabel metal3 12623 14860 12623 14860 4 WL[16]
rlabel metal3 13823 14860 13823 14860 4 WL[16]
rlabel metal3 12023 15760 12023 15760 4 WL[17]
rlabel metal3 13823 19360 13823 19360 4 WL[21]
rlabel metal3 14423 21160 14423 21160 4 WL[23]
rlabel metal3 13823 17560 13823 17560 4 WL[19]
rlabel metal3 13223 14860 13223 14860 4 WL[16]
rlabel metal3 13223 16660 13223 16660 4 WL[18]
rlabel metal3 14423 18460 14423 18460 4 WL[20]
rlabel metal3 14423 20260 14423 20260 4 WL[22]
rlabel metal3 14423 17560 14423 17560 4 WL[19]
rlabel metal3 12623 20260 12623 20260 4 WL[22]
rlabel metal3 13721 14860 13721 14860 4 WL[16]
rlabel metal3 16121 14860 16121 14860 4 WL[16]
rlabel metal3 16121 15760 16121 15760 4 WL[17]
rlabel metal3 16121 16660 16121 16660 4 WL[18]
rlabel metal3 12623 21160 12623 21160 4 WL[23]
rlabel metal3 16121 17560 16121 17560 4 WL[19]
rlabel metal3 16121 18460 16121 18460 4 WL[20]
rlabel metal3 16121 19360 16121 19360 4 WL[21]
rlabel metal3 12023 14860 12023 14860 4 WL[16]
rlabel metal3 13823 16660 13823 16660 4 WL[18]
rlabel metal3 16121 20260 16121 20260 4 WL[22]
rlabel metal3 16121 21160 16121 21160 4 WL[23]
rlabel metal3 13721 15760 13721 15760 4 WL[17]
rlabel metal3 21577 21160 21577 21160 4 WL[23]
rlabel metal3 21577 20260 21577 20260 4 WL[22]
rlabel metal3 21577 19360 21577 19360 4 WL[21]
rlabel metal3 21577 18460 21577 18460 4 WL[20]
rlabel metal3 20479 18460 20479 18460 4 WL[20]
rlabel metal3 20479 19360 20479 19360 4 WL[21]
rlabel metal3 20479 20260 20479 20260 4 WL[22]
rlabel metal3 20479 21160 20479 21160 4 WL[23]
rlabel metal3 20377 21160 20377 21160 4 WL[23]
rlabel metal3 20377 20260 20377 20260 4 WL[22]
rlabel metal3 20377 19360 20377 19360 4 WL[21]
rlabel metal3 20377 18460 20377 18460 4 WL[20]
rlabel metal3 21519 21160 21519 21160 4 WL[23]
rlabel metal3 20977 18460 20977 18460 4 WL[20]
rlabel metal3 19177 21160 19177 21160 4 WL[23]
rlabel metal3 20977 20260 20977 20260 4 WL[22]
rlabel metal3 19777 21160 19777 21160 4 WL[23]
rlabel metal3 19177 20260 19177 20260 4 WL[22]
rlabel metal3 19177 19360 19177 19360 4 WL[21]
rlabel metal3 19177 18460 19177 18460 4 WL[20]
rlabel metal3 19279 18460 19279 18460 4 WL[20]
rlabel metal3 19279 19360 19279 19360 4 WL[21]
rlabel metal3 19279 20260 19279 20260 4 WL[22]
rlabel metal3 19279 21160 19279 21160 4 WL[23]
rlabel metal3 19777 20260 19777 20260 4 WL[22]
rlabel metal3 19777 19360 19777 19360 4 WL[21]
rlabel metal3 19777 18460 19777 18460 4 WL[20]
rlabel metal3 21519 18460 21519 18460 4 WL[20]
rlabel metal3 20977 19360 20977 19360 4 WL[21]
rlabel metal3 21519 20260 21519 20260 4 WL[22]
rlabel metal3 20977 21160 20977 21160 4 WL[23]
rlabel metal3 21519 19360 21519 19360 4 WL[21]
rlabel metal3 18079 18460 18079 18460 4 WL[20]
rlabel metal3 18079 19360 18079 19360 4 WL[21]
rlabel metal3 18079 20260 18079 20260 4 WL[22]
rlabel metal3 18079 21160 18079 21160 4 WL[23]
rlabel metal3 18577 21160 18577 21160 4 WL[23]
rlabel metal3 18577 20260 18577 20260 4 WL[22]
rlabel metal3 18577 19360 18577 19360 4 WL[21]
rlabel metal3 18577 18460 18577 18460 4 WL[20]
rlabel metal3 16879 18460 16879 18460 4 WL[20]
rlabel metal3 17977 21160 17977 21160 4 WL[23]
rlabel metal3 17977 20260 17977 20260 4 WL[22]
rlabel metal3 17977 19360 17977 19360 4 WL[21]
rlabel metal3 17977 18460 17977 18460 4 WL[20]
rlabel metal3 16879 19360 16879 19360 4 WL[21]
rlabel metal3 16879 20260 16879 20260 4 WL[22]
rlabel metal3 16879 21160 16879 21160 4 WL[23]
rlabel metal3 17377 21160 17377 21160 4 WL[23]
rlabel metal3 17377 20260 17377 20260 4 WL[22]
rlabel metal3 17377 19360 17377 19360 4 WL[21]
rlabel metal3 17377 18460 17377 18460 4 WL[20]
rlabel metal3 18079 15760 18079 15760 4 WL[17]
rlabel metal3 18079 16660 18079 16660 4 WL[18]
rlabel metal3 18079 17560 18079 17560 4 WL[19]
rlabel metal3 16879 14860 16879 14860 4 WL[16]
rlabel metal3 16879 15760 16879 15760 4 WL[17]
rlabel metal3 17977 17560 17977 17560 4 WL[19]
rlabel metal3 17977 16660 17977 16660 4 WL[18]
rlabel metal3 17977 15760 17977 15760 4 WL[17]
rlabel metal3 17977 14860 17977 14860 4 WL[16]
rlabel metal3 16879 16660 16879 16660 4 WL[18]
rlabel metal3 16879 17560 16879 17560 4 WL[19]
rlabel metal3 18079 14860 18079 14860 4 WL[16]
rlabel metal3 18577 16660 18577 16660 4 WL[18]
rlabel metal3 18577 15760 18577 15760 4 WL[17]
rlabel metal3 18577 14860 18577 14860 4 WL[16]
rlabel metal3 18577 17560 18577 17560 4 WL[19]
rlabel metal3 17377 17560 17377 17560 4 WL[19]
rlabel metal3 17377 16660 17377 16660 4 WL[18]
rlabel metal3 17377 15760 17377 15760 4 WL[17]
rlabel metal3 17377 14860 17377 14860 4 WL[16]
rlabel metal3 19777 14860 19777 14860 4 WL[16]
rlabel metal3 19279 14860 19279 14860 4 WL[16]
rlabel metal3 19177 17560 19177 17560 4 WL[19]
rlabel metal3 19177 16660 19177 16660 4 WL[18]
rlabel metal3 21519 14860 21519 14860 4 WL[16]
rlabel metal3 19177 15760 19177 15760 4 WL[17]
rlabel metal3 21519 15760 21519 15760 4 WL[17]
rlabel metal3 20977 15760 20977 15760 4 WL[17]
rlabel metal3 20977 16660 20977 16660 4 WL[18]
rlabel metal3 19177 14860 19177 14860 4 WL[16]
rlabel metal3 21519 17560 21519 17560 4 WL[19]
rlabel metal3 20479 15760 20479 15760 4 WL[17]
rlabel metal3 20479 16660 20479 16660 4 WL[18]
rlabel metal3 19279 15760 19279 15760 4 WL[17]
rlabel metal3 19279 16660 19279 16660 4 WL[18]
rlabel metal3 19279 17560 19279 17560 4 WL[19]
rlabel metal3 20479 17560 20479 17560 4 WL[19]
rlabel metal3 21577 15760 21577 15760 4 WL[17]
rlabel metal3 21577 14860 21577 14860 4 WL[16]
rlabel metal3 20377 17560 20377 17560 4 WL[19]
rlabel metal3 20377 16660 20377 16660 4 WL[18]
rlabel metal3 20977 14860 20977 14860 4 WL[16]
rlabel metal3 20377 15760 20377 15760 4 WL[17]
rlabel metal3 20977 17560 20977 17560 4 WL[19]
rlabel metal3 20377 14860 20377 14860 4 WL[16]
rlabel metal3 21577 17560 21577 17560 4 WL[19]
rlabel metal3 21577 16660 21577 16660 4 WL[18]
rlabel metal3 21519 16660 21519 16660 4 WL[18]
rlabel metal3 19777 17560 19777 17560 4 WL[19]
rlabel metal3 20479 14860 20479 14860 4 WL[16]
rlabel metal3 19777 16660 19777 16660 4 WL[18]
rlabel metal3 19777 15760 19777 15760 4 WL[17]
rlabel metal3 10719 26560 10719 26560 4 WL[29]
rlabel metal3 10719 27460 10719 27460 4 WL[30]
rlabel metal3 10719 28360 10719 28360 4 WL[31]
rlabel metal3 9679 25660 9679 25660 4 WL[28]
rlabel metal3 9679 26560 9679 26560 4 WL[29]
rlabel metal3 9679 27460 9679 27460 4 WL[30]
rlabel metal3 9679 28360 9679 28360 4 WL[31]
rlabel metal3 11423 26560 11423 26560 4 WL[29]
rlabel metal3 11481 28360 11481 28360 4 WL[31]
rlabel metal3 11481 27460 11481 27460 4 WL[30]
rlabel metal3 11481 26560 11481 26560 4 WL[29]
rlabel metal3 11481 25660 11481 25660 4 WL[28]
rlabel metal3 11423 27460 11423 27460 4 WL[30]
rlabel metal3 11423 28360 11423 28360 4 WL[31]
rlabel metal3 11423 25660 11423 25660 4 WL[28]
rlabel metal3 9577 28360 9577 28360 4 WL[31]
rlabel metal3 9577 27460 9577 27460 4 WL[30]
rlabel metal3 9577 26560 9577 26560 4 WL[29]
rlabel metal3 9577 25660 9577 25660 4 WL[28]
rlabel metal3 10719 25660 10719 25660 4 WL[28]
rlabel metal3 10177 28360 10177 28360 4 WL[31]
rlabel metal3 10177 27460 10177 27460 4 WL[30]
rlabel metal3 10177 26560 10177 26560 4 WL[29]
rlabel metal3 10177 25660 10177 25660 4 WL[28]
rlabel metal3 10777 28360 10777 28360 4 WL[31]
rlabel metal3 10777 27460 10777 27460 4 WL[30]
rlabel metal3 10777 26560 10777 26560 4 WL[29]
rlabel metal3 10777 25660 10777 25660 4 WL[28]
rlabel metal3 8377 28360 8377 28360 4 WL[31]
rlabel metal3 8377 27460 8377 27460 4 WL[30]
rlabel metal3 8377 26560 8377 26560 4 WL[29]
rlabel metal3 8377 25660 8377 25660 4 WL[28]
rlabel metal3 7279 28360 7279 28360 4 WL[31]
rlabel metal3 8977 28360 8977 28360 4 WL[31]
rlabel metal3 8977 27460 8977 27460 4 WL[30]
rlabel metal3 8977 26560 8977 26560 4 WL[29]
rlabel metal3 8977 25660 8977 25660 4 WL[28]
rlabel metal3 8479 28360 8479 28360 4 WL[31]
rlabel metal3 8479 27460 8479 27460 4 WL[30]
rlabel metal3 7279 25660 7279 25660 4 WL[28]
rlabel metal3 7279 26560 7279 26560 4 WL[29]
rlabel metal3 7279 27460 7279 27460 4 WL[30]
rlabel metal3 7177 28360 7177 28360 4 WL[31]
rlabel metal3 7177 27460 7177 27460 4 WL[30]
rlabel metal3 7177 26560 7177 26560 4 WL[29]
rlabel metal3 7177 25660 7177 25660 4 WL[28]
rlabel metal3 8479 25660 8479 25660 4 WL[28]
rlabel metal3 8479 26560 8479 26560 4 WL[29]
rlabel metal3 7777 28360 7777 28360 4 WL[31]
rlabel metal3 7777 27460 7777 27460 4 WL[30]
rlabel metal3 7777 26560 7777 26560 4 WL[29]
rlabel metal3 7777 25660 7777 25660 4 WL[28]
rlabel metal3 8977 22060 8977 22060 4 WL[24]
rlabel metal3 7177 23860 7177 23860 4 WL[26]
rlabel metal3 7777 22960 7777 22960 4 WL[25]
rlabel metal3 7777 22060 7777 22060 4 WL[24]
rlabel metal3 7279 24760 7279 24760 4 WL[27]
rlabel metal3 8977 24760 8977 24760 4 WL[27]
rlabel metal3 8977 23860 8977 23860 4 WL[26]
rlabel metal3 7279 22060 7279 22060 4 WL[24]
rlabel metal3 7177 22960 7177 22960 4 WL[25]
rlabel metal3 7177 22060 7177 22060 4 WL[24]
rlabel metal3 7777 24760 7777 24760 4 WL[27]
rlabel metal3 7777 23860 7777 23860 4 WL[26]
rlabel metal3 8377 22960 8377 22960 4 WL[25]
rlabel metal3 8377 22060 8377 22060 4 WL[24]
rlabel metal3 7279 22960 7279 22960 4 WL[25]
rlabel metal3 8479 22960 8479 22960 4 WL[25]
rlabel metal3 8479 23860 8479 23860 4 WL[26]
rlabel metal3 8479 24760 8479 24760 4 WL[27]
rlabel metal3 8479 22060 8479 22060 4 WL[24]
rlabel metal3 7279 23860 7279 23860 4 WL[26]
rlabel metal3 8377 24760 8377 24760 4 WL[27]
rlabel metal3 8377 23860 8377 23860 4 WL[26]
rlabel metal3 7177 24760 7177 24760 4 WL[27]
rlabel metal3 8977 22960 8977 22960 4 WL[25]
rlabel metal3 11423 22060 11423 22060 4 WL[24]
rlabel metal3 11481 24760 11481 24760 4 WL[27]
rlabel metal3 11481 23860 11481 23860 4 WL[26]
rlabel metal3 9577 24760 9577 24760 4 WL[27]
rlabel metal3 9577 23860 9577 23860 4 WL[26]
rlabel metal3 10177 22960 10177 22960 4 WL[25]
rlabel metal3 10177 22060 10177 22060 4 WL[24]
rlabel metal3 10719 23860 10719 23860 4 WL[26]
rlabel metal3 10719 24760 10719 24760 4 WL[27]
rlabel metal3 10719 22060 10719 22060 4 WL[24]
rlabel metal3 11423 24760 11423 24760 4 WL[27]
rlabel metal3 11423 23860 11423 23860 4 WL[26]
rlabel metal3 11481 22960 11481 22960 4 WL[25]
rlabel metal3 11481 22060 11481 22060 4 WL[24]
rlabel metal3 10177 24760 10177 24760 4 WL[27]
rlabel metal3 10177 23860 10177 23860 4 WL[26]
rlabel metal3 9679 23860 9679 23860 4 WL[26]
rlabel metal3 10777 22960 10777 22960 4 WL[25]
rlabel metal3 10777 22060 10777 22060 4 WL[24]
rlabel metal3 10719 22960 10719 22960 4 WL[25]
rlabel metal3 9679 24760 9679 24760 4 WL[27]
rlabel metal3 11423 22960 11423 22960 4 WL[25]
rlabel metal3 9679 22060 9679 22060 4 WL[24]
rlabel metal3 9577 22960 9577 22960 4 WL[25]
rlabel metal3 9577 22060 9577 22060 4 WL[24]
rlabel metal3 9679 22960 9679 22960 4 WL[25]
rlabel metal3 10777 24760 10777 24760 4 WL[27]
rlabel metal3 10777 23860 10777 23860 4 WL[26]
rlabel metal3 2423 27460 2423 27460 4 WL[30]
rlabel metal3 2423 26560 2423 26560 4 WL[29]
rlabel metal3 2423 25660 2423 25660 4 WL[28]
rlabel metal3 2423 24760 2423 24760 4 WL[27]
rlabel metal3 5321 27460 5321 27460 4 WL[30]
rlabel metal3 2423 23860 2423 23860 4 WL[26]
rlabel metal3 4121 23860 4121 23860 4 WL[26]
rlabel metal3 4121 28360 4121 28360 4 WL[31]
rlabel metal3 4121 26560 4121 26560 4 WL[29]
rlabel metal3 4121 24760 4121 24760 4 WL[27]
rlabel metal3 1721 26560 1721 26560 4 WL[29]
rlabel metal3 5321 25660 5321 25660 4 WL[28]
rlabel metal3 5321 28360 5321 28360 4 WL[31]
rlabel metal3 1823 22960 1823 22960 4 WL[25]
rlabel metal3 5321 26560 5321 26560 4 WL[29]
rlabel metal3 5321 24760 5321 24760 4 WL[27]
rlabel metal3 5321 23860 5321 23860 4 WL[26]
rlabel metal3 3023 22960 3023 22960 4 WL[25]
rlabel metal3 3023 22060 3023 22060 4 WL[24]
rlabel metal3 3023 28360 3023 28360 4 WL[31]
rlabel metal3 3023 27460 3023 27460 4 WL[30]
rlabel metal3 3023 26560 3023 26560 4 WL[29]
rlabel metal3 3023 25660 3023 25660 4 WL[28]
rlabel metal3 3023 24760 3023 24760 4 WL[27]
rlabel metal3 3023 23860 3023 23860 4 WL[26]
rlabel metal3 2921 24760 2921 24760 4 WL[27]
rlabel metal3 2921 23860 2921 23860 4 WL[26]
rlabel metal3 2921 25660 2921 25660 4 WL[28]
rlabel metal3 1823 22060 1823 22060 4 WL[24]
rlabel metal3 1823 28360 1823 28360 4 WL[31]
rlabel metal3 3623 22960 3623 22960 4 WL[25]
rlabel metal3 2921 26560 2921 26560 4 WL[29]
rlabel metal3 3623 22060 3623 22060 4 WL[24]
rlabel metal3 3623 28360 3623 28360 4 WL[31]
rlabel metal3 3623 27460 3623 27460 4 WL[30]
rlabel metal3 3623 26560 3623 26560 4 WL[29]
rlabel metal3 3623 25660 3623 25660 4 WL[28]
rlabel metal3 3623 24760 3623 24760 4 WL[27]
rlabel metal3 2921 27460 2921 27460 4 WL[30]
rlabel metal3 2921 28360 2921 28360 4 WL[31]
rlabel metal3 3623 23860 3623 23860 4 WL[26]
rlabel metal3 1823 27460 1823 27460 4 WL[30]
rlabel metal3 4121 22060 4121 22060 4 WL[24]
rlabel metal3 1721 22960 1721 22960 4 WL[25]
rlabel metal3 6079 22060 6079 22060 4 WL[24]
rlabel metal3 4121 22960 4121 22960 4 WL[25]
rlabel metal3 1823 26560 1823 26560 4 WL[29]
rlabel metal3 4223 22960 4223 22960 4 WL[25]
rlabel metal3 4223 22060 4223 22060 4 WL[24]
rlabel metal3 1823 25660 1823 25660 4 WL[28]
rlabel metal3 5321 22960 5321 22960 4 WL[25]
rlabel metal3 4223 28360 4223 28360 4 WL[31]
rlabel metal3 4223 27460 4223 27460 4 WL[30]
rlabel metal3 5321 22060 5321 22060 4 WL[24]
rlabel metal3 4223 26560 4223 26560 4 WL[29]
rlabel metal3 4223 25660 4223 25660 4 WL[28]
rlabel metal3 4223 24760 4223 24760 4 WL[27]
rlabel metal3 4223 23860 4223 23860 4 WL[26]
rlabel metal3 1823 24760 1823 24760 4 WL[27]
rlabel metal3 1823 23860 1823 23860 4 WL[26]
rlabel metal3 2921 22060 2921 22060 4 WL[24]
rlabel metal3 2921 22960 2921 22960 4 WL[25]
rlabel metal3 1721 28360 1721 28360 4 WL[31]
rlabel metal3 4823 22960 4823 22960 4 WL[25]
rlabel metal3 4823 22060 4823 22060 4 WL[24]
rlabel metal3 1721 27460 1721 27460 4 WL[30]
rlabel metal3 4121 27460 4121 27460 4 WL[30]
rlabel metal3 4823 28360 4823 28360 4 WL[31]
rlabel metal3 6079 27460 6079 27460 4 WL[30]
rlabel metal3 4823 27460 4823 27460 4 WL[30]
rlabel metal3 4823 26560 4823 26560 4 WL[29]
rlabel metal3 4823 25660 4823 25660 4 WL[28]
rlabel metal3 4823 24760 4823 24760 4 WL[27]
rlabel metal3 4823 23860 4823 23860 4 WL[26]
rlabel metal3 4121 25660 4121 25660 4 WL[28]
rlabel metal3 1721 24760 1721 24760 4 WL[27]
rlabel metal3 6079 28360 6079 28360 4 WL[31]
rlabel metal3 1721 23860 1721 23860 4 WL[26]
rlabel metal3 6079 26560 6079 26560 4 WL[29]
rlabel metal3 6079 25660 6079 25660 4 WL[28]
rlabel metal3 6079 24760 6079 24760 4 WL[27]
rlabel metal3 1721 25660 1721 25660 4 WL[28]
rlabel metal3 6079 23860 6079 23860 4 WL[26]
rlabel metal3 1721 22060 1721 22060 4 WL[24]
rlabel metal3 2423 22960 2423 22960 4 WL[25]
rlabel metal3 2423 22060 2423 22060 4 WL[24]
rlabel metal3 6079 22960 6079 22960 4 WL[25]
rlabel metal3 2423 28360 2423 28360 4 WL[31]
rlabel metal3 6577 22960 6577 22960 4 WL[25]
rlabel metal3 6577 22060 6577 22060 4 WL[24]
rlabel metal3 6577 28360 6577 28360 4 WL[31]
rlabel metal3 6577 27460 6577 27460 4 WL[30]
rlabel metal3 6577 26560 6577 26560 4 WL[29]
rlabel metal3 6577 25660 6577 25660 4 WL[28]
rlabel metal3 6577 24760 6577 24760 4 WL[27]
rlabel metal3 6577 23860 6577 23860 4 WL[26]
rlabel metal3 2423 17560 2423 17560 4 WL[19]
rlabel metal3 2423 16660 2423 16660 4 WL[18]
rlabel metal3 2423 15760 2423 15760 4 WL[17]
rlabel metal3 2423 14860 2423 14860 4 WL[16]
rlabel metal3 6079 20260 6079 20260 4 WL[22]
rlabel metal3 6079 15760 6079 15760 4 WL[17]
rlabel metal3 1721 14860 1721 14860 4 WL[16]
rlabel metal3 5321 17560 5321 17560 4 WL[19]
rlabel metal3 4823 21160 4823 21160 4 WL[23]
rlabel metal3 4823 20260 4823 20260 4 WL[22]
rlabel metal3 4823 19360 4823 19360 4 WL[21]
rlabel metal3 4823 18460 4823 18460 4 WL[20]
rlabel metal3 4823 17560 4823 17560 4 WL[19]
rlabel metal3 4823 16660 4823 16660 4 WL[18]
rlabel metal3 6079 19360 6079 19360 4 WL[21]
rlabel metal3 4823 15760 4823 15760 4 WL[17]
rlabel metal3 4823 14860 4823 14860 4 WL[16]
rlabel metal3 1823 21160 1823 21160 4 WL[23]
rlabel metal3 1823 20260 1823 20260 4 WL[22]
rlabel metal3 1823 19360 1823 19360 4 WL[21]
rlabel metal3 1823 18460 1823 18460 4 WL[20]
rlabel metal3 3623 21160 3623 21160 4 WL[23]
rlabel metal3 3623 20260 3623 20260 4 WL[22]
rlabel metal3 2921 15760 2921 15760 4 WL[17]
rlabel metal3 2921 16660 2921 16660 4 WL[18]
rlabel metal3 3623 19360 3623 19360 4 WL[21]
rlabel metal3 3623 18460 3623 18460 4 WL[20]
rlabel metal3 3623 17560 3623 17560 4 WL[19]
rlabel metal3 2921 14860 2921 14860 4 WL[16]
rlabel metal3 2921 18460 2921 18460 4 WL[20]
rlabel metal3 3623 16660 3623 16660 4 WL[18]
rlabel metal3 3623 15760 3623 15760 4 WL[17]
rlabel metal3 3623 14860 3623 14860 4 WL[16]
rlabel metal3 1823 17560 1823 17560 4 WL[19]
rlabel metal3 1721 21160 1721 21160 4 WL[23]
rlabel metal3 1721 16660 1721 16660 4 WL[18]
rlabel metal3 1721 15760 1721 15760 4 WL[17]
rlabel metal3 2921 17560 2921 17560 4 WL[19]
rlabel metal3 1823 16660 1823 16660 4 WL[18]
rlabel metal3 2921 19360 2921 19360 4 WL[21]
rlabel metal3 2921 20260 2921 20260 4 WL[22]
rlabel metal3 1823 15760 1823 15760 4 WL[17]
rlabel metal3 6577 21160 6577 21160 4 WL[23]
rlabel metal3 6577 20260 6577 20260 4 WL[22]
rlabel metal3 5321 21160 5321 21160 4 WL[23]
rlabel metal3 5321 20260 5321 20260 4 WL[22]
rlabel metal3 5321 19360 5321 19360 4 WL[21]
rlabel metal3 6577 19360 6577 19360 4 WL[21]
rlabel metal3 6577 18460 6577 18460 4 WL[20]
rlabel metal3 6577 17560 6577 17560 4 WL[19]
rlabel metal3 6577 16660 6577 16660 4 WL[18]
rlabel metal3 6577 15760 6577 15760 4 WL[17]
rlabel metal3 6577 14860 6577 14860 4 WL[16]
rlabel metal3 2921 21160 2921 21160 4 WL[23]
rlabel metal3 6079 21160 6079 21160 4 WL[23]
rlabel metal3 1823 14860 1823 14860 4 WL[16]
rlabel metal3 1721 17560 1721 17560 4 WL[19]
rlabel metal3 5321 18460 5321 18460 4 WL[20]
rlabel metal3 6079 17560 6079 17560 4 WL[19]
rlabel metal3 6079 16660 6079 16660 4 WL[18]
rlabel metal3 6079 14860 6079 14860 4 WL[16]
rlabel metal3 2423 21160 2423 21160 4 WL[23]
rlabel metal3 2423 20260 2423 20260 4 WL[22]
rlabel metal3 2423 19360 2423 19360 4 WL[21]
rlabel metal3 4121 18460 4121 18460 4 WL[20]
rlabel metal3 4121 17560 4121 17560 4 WL[19]
rlabel metal3 4121 15760 4121 15760 4 WL[17]
rlabel metal3 1721 18460 1721 18460 4 WL[20]
rlabel metal3 1721 20260 1721 20260 4 WL[22]
rlabel metal3 2423 18460 2423 18460 4 WL[20]
rlabel metal3 5321 16660 5321 16660 4 WL[18]
rlabel metal3 4121 21160 4121 21160 4 WL[23]
rlabel metal3 5321 14860 5321 14860 4 WL[16]
rlabel metal3 4121 20260 4121 20260 4 WL[22]
rlabel metal3 4121 19360 4121 19360 4 WL[21]
rlabel metal3 6079 18460 6079 18460 4 WL[20]
rlabel metal3 3023 21160 3023 21160 4 WL[23]
rlabel metal3 3023 20260 3023 20260 4 WL[22]
rlabel metal3 3023 19360 3023 19360 4 WL[21]
rlabel metal3 4223 21160 4223 21160 4 WL[23]
rlabel metal3 4223 20260 4223 20260 4 WL[22]
rlabel metal3 4223 19360 4223 19360 4 WL[21]
rlabel metal3 4223 18460 4223 18460 4 WL[20]
rlabel metal3 4121 16660 4121 16660 4 WL[18]
rlabel metal3 4223 17560 4223 17560 4 WL[19]
rlabel metal3 4223 16660 4223 16660 4 WL[18]
rlabel metal3 4223 15760 4223 15760 4 WL[17]
rlabel metal3 4223 14860 4223 14860 4 WL[16]
rlabel metal3 3023 18460 3023 18460 4 WL[20]
rlabel metal3 3023 17560 3023 17560 4 WL[19]
rlabel metal3 1721 19360 1721 19360 4 WL[21]
rlabel metal3 3023 16660 3023 16660 4 WL[18]
rlabel metal3 3023 15760 3023 15760 4 WL[17]
rlabel metal3 4121 14860 4121 14860 4 WL[16]
rlabel metal3 5321 15760 5321 15760 4 WL[17]
rlabel metal3 3023 14860 3023 14860 4 WL[16]
rlabel metal3 10719 21160 10719 21160 4 WL[23]
rlabel metal3 10719 20260 10719 20260 4 WL[22]
rlabel metal3 9577 21160 9577 21160 4 WL[23]
rlabel metal3 9577 20260 9577 20260 4 WL[22]
rlabel metal3 9577 19360 9577 19360 4 WL[21]
rlabel metal3 9577 18460 9577 18460 4 WL[20]
rlabel metal3 11423 18460 11423 18460 4 WL[20]
rlabel metal3 11481 21160 11481 21160 4 WL[23]
rlabel metal3 11481 20260 11481 20260 4 WL[22]
rlabel metal3 11481 19360 11481 19360 4 WL[21]
rlabel metal3 11481 18460 11481 18460 4 WL[20]
rlabel metal3 11423 20260 11423 20260 4 WL[22]
rlabel metal3 10177 21160 10177 21160 4 WL[23]
rlabel metal3 10177 20260 10177 20260 4 WL[22]
rlabel metal3 10177 19360 10177 19360 4 WL[21]
rlabel metal3 10177 18460 10177 18460 4 WL[20]
rlabel metal3 10719 18460 10719 18460 4 WL[20]
rlabel metal3 9679 18460 9679 18460 4 WL[20]
rlabel metal3 9679 19360 9679 19360 4 WL[21]
rlabel metal3 9679 20260 9679 20260 4 WL[22]
rlabel metal3 9679 21160 9679 21160 4 WL[23]
rlabel metal3 11423 19360 11423 19360 4 WL[21]
rlabel metal3 11423 21160 11423 21160 4 WL[23]
rlabel metal3 10719 19360 10719 19360 4 WL[21]
rlabel metal3 10777 21160 10777 21160 4 WL[23]
rlabel metal3 10777 20260 10777 20260 4 WL[22]
rlabel metal3 10777 19360 10777 19360 4 WL[21]
rlabel metal3 10777 18460 10777 18460 4 WL[20]
rlabel metal3 8479 18460 8479 18460 4 WL[20]
rlabel metal3 8479 19360 8479 19360 4 WL[21]
rlabel metal3 7279 19360 7279 19360 4 WL[21]
rlabel metal3 7279 20260 7279 20260 4 WL[22]
rlabel metal3 7777 21160 7777 21160 4 WL[23]
rlabel metal3 7777 20260 7777 20260 4 WL[22]
rlabel metal3 7777 19360 7777 19360 4 WL[21]
rlabel metal3 8377 21160 8377 21160 4 WL[23]
rlabel metal3 8377 20260 8377 20260 4 WL[22]
rlabel metal3 8377 19360 8377 19360 4 WL[21]
rlabel metal3 8377 18460 8377 18460 4 WL[20]
rlabel metal3 7777 18460 7777 18460 4 WL[20]
rlabel metal3 7279 21160 7279 21160 4 WL[23]
rlabel metal3 8479 20260 8479 20260 4 WL[22]
rlabel metal3 8977 18460 8977 18460 4 WL[20]
rlabel metal3 8479 21160 8479 21160 4 WL[23]
rlabel metal3 8977 19360 8977 19360 4 WL[21]
rlabel metal3 7279 18460 7279 18460 4 WL[20]
rlabel metal3 7177 21160 7177 21160 4 WL[23]
rlabel metal3 7177 20260 7177 20260 4 WL[22]
rlabel metal3 7177 19360 7177 19360 4 WL[21]
rlabel metal3 7177 18460 7177 18460 4 WL[20]
rlabel metal3 8977 21160 8977 21160 4 WL[23]
rlabel metal3 8977 20260 8977 20260 4 WL[22]
rlabel metal3 8479 15760 8479 15760 4 WL[17]
rlabel metal3 8977 14860 8977 14860 4 WL[16]
rlabel metal3 8479 16660 8479 16660 4 WL[18]
rlabel metal3 8377 17560 8377 17560 4 WL[19]
rlabel metal3 8377 16660 8377 16660 4 WL[18]
rlabel metal3 8377 15760 8377 15760 4 WL[17]
rlabel metal3 8377 14860 8377 14860 4 WL[16]
rlabel metal3 7177 14860 7177 14860 4 WL[16]
rlabel metal3 7279 16660 7279 16660 4 WL[18]
rlabel metal3 8977 17560 8977 17560 4 WL[19]
rlabel metal3 7279 17560 7279 17560 4 WL[19]
rlabel metal3 8977 16660 8977 16660 4 WL[18]
rlabel metal3 8479 17560 8479 17560 4 WL[19]
rlabel metal3 7777 17560 7777 17560 4 WL[19]
rlabel metal3 7279 14860 7279 14860 4 WL[16]
rlabel metal3 7777 16660 7777 16660 4 WL[18]
rlabel metal3 7777 15760 7777 15760 4 WL[17]
rlabel metal3 7777 14860 7777 14860 4 WL[16]
rlabel metal3 8479 14860 8479 14860 4 WL[16]
rlabel metal3 7177 17560 7177 17560 4 WL[19]
rlabel metal3 7177 16660 7177 16660 4 WL[18]
rlabel metal3 7177 15760 7177 15760 4 WL[17]
rlabel metal3 7279 15760 7279 15760 4 WL[17]
rlabel metal3 8977 15760 8977 15760 4 WL[17]
rlabel metal3 11423 17560 11423 17560 4 WL[19]
rlabel metal3 10177 17560 10177 17560 4 WL[19]
rlabel metal3 10177 16660 10177 16660 4 WL[18]
rlabel metal3 10177 15760 10177 15760 4 WL[17]
rlabel metal3 10177 14860 10177 14860 4 WL[16]
rlabel metal3 10719 14860 10719 14860 4 WL[16]
rlabel metal3 9679 14860 9679 14860 4 WL[16]
rlabel metal3 9679 15760 9679 15760 4 WL[17]
rlabel metal3 10719 16660 10719 16660 4 WL[18]
rlabel metal3 9679 16660 9679 16660 4 WL[18]
rlabel metal3 9679 17560 9679 17560 4 WL[19]
rlabel metal3 11423 14860 11423 14860 4 WL[16]
rlabel metal3 11423 15760 11423 15760 4 WL[17]
rlabel metal3 11423 16660 11423 16660 4 WL[18]
rlabel metal3 10719 15760 10719 15760 4 WL[17]
rlabel metal3 10777 17560 10777 17560 4 WL[19]
rlabel metal3 10777 16660 10777 16660 4 WL[18]
rlabel metal3 10777 15760 10777 15760 4 WL[17]
rlabel metal3 10777 14860 10777 14860 4 WL[16]
rlabel metal3 11481 17560 11481 17560 4 WL[19]
rlabel metal3 11481 16660 11481 16660 4 WL[18]
rlabel metal3 11481 15760 11481 15760 4 WL[17]
rlabel metal3 10719 17560 10719 17560 4 WL[19]
rlabel metal3 11481 14860 11481 14860 4 WL[16]
rlabel metal3 9577 17560 9577 17560 4 WL[19]
rlabel metal3 9577 16660 9577 16660 4 WL[18]
rlabel metal3 9577 15760 9577 15760 4 WL[17]
rlabel metal3 9577 14860 9577 14860 4 WL[16]
rlabel metal3 11423 11260 11423 11260 4 WL[12]
rlabel metal3 11423 13960 11423 13960 4 WL[15]
rlabel metal3 11423 12160 11423 12160 4 WL[13]
rlabel metal3 9679 11260 9679 11260 4 WL[12]
rlabel metal3 9679 12160 9679 12160 4 WL[13]
rlabel metal3 9679 13060 9679 13060 4 WL[14]
rlabel metal3 11423 13060 11423 13060 4 WL[14]
rlabel metal3 9679 13960 9679 13960 4 WL[15]
rlabel metal3 10719 11260 10719 11260 4 WL[12]
rlabel metal3 10719 12160 10719 12160 4 WL[13]
rlabel metal3 10719 13060 10719 13060 4 WL[14]
rlabel metal3 10719 13960 10719 13960 4 WL[15]
rlabel metal3 11481 13960 11481 13960 4 WL[15]
rlabel metal3 11481 13060 11481 13060 4 WL[14]
rlabel metal3 11481 12160 11481 12160 4 WL[13]
rlabel metal3 11481 11260 11481 11260 4 WL[12]
rlabel metal3 9577 13960 9577 13960 4 WL[15]
rlabel metal3 9577 13060 9577 13060 4 WL[14]
rlabel metal3 9577 12160 9577 12160 4 WL[13]
rlabel metal3 9577 11260 9577 11260 4 WL[12]
rlabel metal3 10177 13960 10177 13960 4 WL[15]
rlabel metal3 10177 13060 10177 13060 4 WL[14]
rlabel metal3 10177 12160 10177 12160 4 WL[13]
rlabel metal3 10177 11260 10177 11260 4 WL[12]
rlabel metal3 10777 13960 10777 13960 4 WL[15]
rlabel metal3 10777 13060 10777 13060 4 WL[14]
rlabel metal3 10777 12160 10777 12160 4 WL[13]
rlabel metal3 10777 11260 10777 11260 4 WL[12]
rlabel metal3 8377 13060 8377 13060 4 WL[14]
rlabel metal3 8377 12160 8377 12160 4 WL[13]
rlabel metal3 8377 11260 8377 11260 4 WL[12]
rlabel metal3 7177 13960 7177 13960 4 WL[15]
rlabel metal3 8977 13960 8977 13960 4 WL[15]
rlabel metal3 8977 13060 8977 13060 4 WL[14]
rlabel metal3 8977 12160 8977 12160 4 WL[13]
rlabel metal3 8977 11260 8977 11260 4 WL[12]
rlabel metal3 7177 13060 7177 13060 4 WL[14]
rlabel metal3 7177 12160 7177 12160 4 WL[13]
rlabel metal3 7177 11260 7177 11260 4 WL[12]
rlabel metal3 8479 13960 8479 13960 4 WL[15]
rlabel metal3 8479 11260 8479 11260 4 WL[12]
rlabel metal3 8479 12160 8479 12160 4 WL[13]
rlabel metal3 7279 11260 7279 11260 4 WL[12]
rlabel metal3 7279 12160 7279 12160 4 WL[13]
rlabel metal3 7777 13960 7777 13960 4 WL[15]
rlabel metal3 7777 13060 7777 13060 4 WL[14]
rlabel metal3 7777 12160 7777 12160 4 WL[13]
rlabel metal3 7777 11260 7777 11260 4 WL[12]
rlabel metal3 7279 13060 7279 13060 4 WL[14]
rlabel metal3 7279 13960 7279 13960 4 WL[15]
rlabel metal3 8479 13060 8479 13060 4 WL[14]
rlabel metal3 8377 13960 8377 13960 4 WL[15]
rlabel metal3 7177 10360 7177 10360 4 WL[11]
rlabel metal3 7177 9460 7177 9460 4 WL[10]
rlabel metal3 7777 10360 7777 10360 4 WL[11]
rlabel metal3 8977 10360 8977 10360 4 WL[11]
rlabel metal3 8977 9460 8977 9460 4 WL[10]
rlabel metal3 8977 8560 8977 8560 4 WL[9]
rlabel metal3 8977 7660 8977 7660 4 WL[8]
rlabel metal3 7777 9460 7777 9460 4 WL[10]
rlabel metal3 7777 8560 7777 8560 4 WL[9]
rlabel metal3 7777 7660 7777 7660 4 WL[8]
rlabel metal3 7177 8560 7177 8560 4 WL[9]
rlabel metal3 7177 7660 7177 7660 4 WL[8]
rlabel metal3 8479 10360 8479 10360 4 WL[11]
rlabel metal3 7279 7660 7279 7660 4 WL[8]
rlabel metal3 7279 8560 7279 8560 4 WL[9]
rlabel metal3 7279 9460 7279 9460 4 WL[10]
rlabel metal3 7279 10360 7279 10360 4 WL[11]
rlabel metal3 8377 10360 8377 10360 4 WL[11]
rlabel metal3 8377 9460 8377 9460 4 WL[10]
rlabel metal3 8377 8560 8377 8560 4 WL[9]
rlabel metal3 8377 7660 8377 7660 4 WL[8]
rlabel metal3 8479 8560 8479 8560 4 WL[9]
rlabel metal3 8479 9460 8479 9460 4 WL[10]
rlabel metal3 8479 7660 8479 7660 4 WL[8]
rlabel metal3 11481 9460 11481 9460 4 WL[10]
rlabel metal3 11481 8560 11481 8560 4 WL[9]
rlabel metal3 11481 7660 11481 7660 4 WL[8]
rlabel metal3 9679 8560 9679 8560 4 WL[9]
rlabel metal3 11423 7660 11423 7660 4 WL[8]
rlabel metal3 9679 9460 9679 9460 4 WL[10]
rlabel metal3 9679 10360 9679 10360 4 WL[11]
rlabel metal3 9577 10360 9577 10360 4 WL[11]
rlabel metal3 9577 9460 9577 9460 4 WL[10]
rlabel metal3 9577 8560 9577 8560 4 WL[9]
rlabel metal3 9577 7660 9577 7660 4 WL[8]
rlabel metal3 11423 10360 11423 10360 4 WL[11]
rlabel metal3 10719 7660 10719 7660 4 WL[8]
rlabel metal3 10719 8560 10719 8560 4 WL[9]
rlabel metal3 10719 9460 10719 9460 4 WL[10]
rlabel metal3 10177 10360 10177 10360 4 WL[11]
rlabel metal3 10177 9460 10177 9460 4 WL[10]
rlabel metal3 10177 8560 10177 8560 4 WL[9]
rlabel metal3 10177 7660 10177 7660 4 WL[8]
rlabel metal3 10719 10360 10719 10360 4 WL[11]
rlabel metal3 11423 9460 11423 9460 4 WL[10]
rlabel metal3 11423 8560 11423 8560 4 WL[9]
rlabel metal3 9679 7660 9679 7660 4 WL[8]
rlabel metal3 10777 10360 10777 10360 4 WL[11]
rlabel metal3 10777 9460 10777 9460 4 WL[10]
rlabel metal3 10777 8560 10777 8560 4 WL[9]
rlabel metal3 10777 7660 10777 7660 4 WL[8]
rlabel metal3 11481 10360 11481 10360 4 WL[11]
rlabel metal3 6079 7660 6079 7660 4 WL[8]
rlabel metal3 4823 13960 4823 13960 4 WL[15]
rlabel metal3 2921 12160 2921 12160 4 WL[13]
rlabel metal3 4823 13060 4823 13060 4 WL[14]
rlabel metal3 4823 12160 4823 12160 4 WL[13]
rlabel metal3 4823 11260 4823 11260 4 WL[12]
rlabel metal3 4823 10360 4823 10360 4 WL[11]
rlabel metal3 4823 9460 4823 9460 4 WL[10]
rlabel metal3 2423 13960 2423 13960 4 WL[15]
rlabel metal3 2423 13060 2423 13060 4 WL[14]
rlabel metal3 2423 12160 2423 12160 4 WL[13]
rlabel metal3 2423 11260 2423 11260 4 WL[12]
rlabel metal3 2423 10360 2423 10360 4 WL[11]
rlabel metal3 2423 9460 2423 9460 4 WL[10]
rlabel metal3 2423 8560 2423 8560 4 WL[9]
rlabel metal3 2423 7660 2423 7660 4 WL[8]
rlabel metal3 4823 8560 4823 8560 4 WL[9]
rlabel metal3 4823 7660 4823 7660 4 WL[8]
rlabel metal3 2921 9460 2921 9460 4 WL[10]
rlabel metal3 2921 8560 2921 8560 4 WL[9]
rlabel metal3 2921 7660 2921 7660 4 WL[8]
rlabel metal3 5321 13060 5321 13060 4 WL[14]
rlabel metal3 4223 12160 4223 12160 4 WL[13]
rlabel metal3 6079 13960 6079 13960 4 WL[15]
rlabel metal3 6079 13060 6079 13060 4 WL[14]
rlabel metal3 6079 11260 6079 11260 4 WL[12]
rlabel metal3 6079 10360 6079 10360 4 WL[11]
rlabel metal3 4223 11260 4223 11260 4 WL[12]
rlabel metal3 4223 10360 4223 10360 4 WL[11]
rlabel metal3 2921 11260 2921 11260 4 WL[12]
rlabel metal3 2921 10360 2921 10360 4 WL[11]
rlabel metal3 5321 13960 5321 13960 4 WL[15]
rlabel metal3 5321 12160 5321 12160 4 WL[13]
rlabel metal3 5321 11260 5321 11260 4 WL[12]
rlabel metal3 5321 9460 5321 9460 4 WL[10]
rlabel metal3 1823 13960 1823 13960 4 WL[15]
rlabel metal3 1823 13060 1823 13060 4 WL[14]
rlabel metal3 1823 12160 1823 12160 4 WL[13]
rlabel metal3 4223 9460 4223 9460 4 WL[10]
rlabel metal3 1823 11260 1823 11260 4 WL[12]
rlabel metal3 1823 10360 1823 10360 4 WL[11]
rlabel metal3 1823 9460 1823 9460 4 WL[10]
rlabel metal3 1823 8560 1823 8560 4 WL[9]
rlabel metal3 3023 13960 3023 13960 4 WL[15]
rlabel metal3 3023 13060 3023 13060 4 WL[14]
rlabel metal3 3023 12160 3023 12160 4 WL[13]
rlabel metal3 1823 7660 1823 7660 4 WL[8]
rlabel metal3 4223 8560 4223 8560 4 WL[9]
rlabel metal3 4223 7660 4223 7660 4 WL[8]
rlabel metal3 4223 13960 4223 13960 4 WL[15]
rlabel metal3 4223 13060 4223 13060 4 WL[14]
rlabel metal3 4121 12160 4121 12160 4 WL[13]
rlabel metal3 6079 9460 6079 9460 4 WL[10]
rlabel metal3 1721 13960 1721 13960 4 WL[15]
rlabel metal3 3023 11260 3023 11260 4 WL[12]
rlabel metal3 3023 10360 3023 10360 4 WL[11]
rlabel metal3 3023 9460 3023 9460 4 WL[10]
rlabel metal3 3023 8560 3023 8560 4 WL[9]
rlabel metal3 3023 7660 3023 7660 4 WL[8]
rlabel metal3 1721 12160 1721 12160 4 WL[13]
rlabel metal3 1721 11260 1721 11260 4 WL[12]
rlabel metal3 1721 10360 1721 10360 4 WL[11]
rlabel metal3 1721 9460 1721 9460 4 WL[10]
rlabel metal3 1721 8560 1721 8560 4 WL[9]
rlabel metal3 5321 8560 5321 8560 4 WL[9]
rlabel metal3 5321 7660 5321 7660 4 WL[8]
rlabel metal3 1721 7660 1721 7660 4 WL[8]
rlabel metal3 6079 8560 6079 8560 4 WL[9]
rlabel metal3 1721 13060 1721 13060 4 WL[14]
rlabel metal3 2921 13060 2921 13060 4 WL[14]
rlabel metal3 2921 13960 2921 13960 4 WL[15]
rlabel metal3 6577 13960 6577 13960 4 WL[15]
rlabel metal3 6577 13060 6577 13060 4 WL[14]
rlabel metal3 6577 12160 6577 12160 4 WL[13]
rlabel metal3 6577 11260 6577 11260 4 WL[12]
rlabel metal3 3623 13960 3623 13960 4 WL[15]
rlabel metal3 3623 13060 3623 13060 4 WL[14]
rlabel metal3 3623 12160 3623 12160 4 WL[13]
rlabel metal3 3623 11260 3623 11260 4 WL[12]
rlabel metal3 3623 10360 3623 10360 4 WL[11]
rlabel metal3 3623 9460 3623 9460 4 WL[10]
rlabel metal3 3623 8560 3623 8560 4 WL[9]
rlabel metal3 3623 7660 3623 7660 4 WL[8]
rlabel metal3 4121 11260 4121 11260 4 WL[12]
rlabel metal3 4121 10360 4121 10360 4 WL[11]
rlabel metal3 4121 8560 4121 8560 4 WL[9]
rlabel metal3 4121 7660 4121 7660 4 WL[8]
rlabel metal3 6577 10360 6577 10360 4 WL[11]
rlabel metal3 6577 9460 6577 9460 4 WL[10]
rlabel metal3 6577 8560 6577 8560 4 WL[9]
rlabel metal3 4121 9460 4121 9460 4 WL[10]
rlabel metal3 4121 13960 4121 13960 4 WL[15]
rlabel metal3 5321 10360 5321 10360 4 WL[11]
rlabel metal3 4121 13060 4121 13060 4 WL[14]
rlabel metal3 6577 7660 6577 7660 4 WL[8]
rlabel metal3 6079 12160 6079 12160 4 WL[13]
rlabel metal3 4223 6760 4223 6760 4 WL[7]
rlabel metal3 4223 5860 4223 5860 4 WL[6]
rlabel metal3 4223 4960 4223 4960 4 WL[5]
rlabel metal3 4223 4060 4223 4060 4 WL[4]
rlabel metal3 6577 6760 6577 6760 4 WL[7]
rlabel metal3 6577 5860 6577 5860 4 WL[6]
rlabel metal3 6577 4960 6577 4960 4 WL[5]
rlabel metal3 6577 4060 6577 4060 4 WL[4]
rlabel metal3 5321 6760 5321 6760 4 WL[7]
rlabel metal3 5321 5860 5321 5860 4 WL[6]
rlabel metal3 6079 6760 6079 6760 4 WL[7]
rlabel metal3 6079 5860 6079 5860 4 WL[6]
rlabel metal3 6079 4960 6079 4960 4 WL[5]
rlabel metal3 6079 4060 6079 4060 4 WL[4]
rlabel metal3 5321 4960 5321 4960 4 WL[5]
rlabel metal3 5321 4060 5321 4060 4 WL[4]
rlabel metal3 4823 6760 4823 6760 4 WL[7]
rlabel metal3 4823 5860 4823 5860 4 WL[6]
rlabel metal3 4823 4960 4823 4960 4 WL[5]
rlabel metal3 4823 4060 4823 4060 4 WL[4]
rlabel metal3 1721 4960 1721 4960 4 WL[5]
rlabel metal3 2921 4960 2921 4960 4 WL[5]
rlabel metal3 2921 5860 2921 5860 4 WL[6]
rlabel metal3 1721 5860 1721 5860 4 WL[6]
rlabel metal3 1823 6760 1823 6760 4 WL[7]
rlabel metal3 1721 6760 1721 6760 4 WL[7]
rlabel metal3 1823 5860 1823 5860 4 WL[6]
rlabel metal3 1823 4960 1823 4960 4 WL[5]
rlabel metal3 1823 4060 1823 4060 4 WL[4]
rlabel metal3 2921 4060 2921 4060 4 WL[4]
rlabel metal3 1721 4060 1721 4060 4 WL[4]
rlabel metal3 2921 6760 2921 6760 4 WL[7]
rlabel metal3 3023 6760 3023 6760 4 WL[7]
rlabel metal3 3623 6760 3623 6760 4 WL[7]
rlabel metal3 3623 5860 3623 5860 4 WL[6]
rlabel metal3 3623 4960 3623 4960 4 WL[5]
rlabel metal3 3623 4060 3623 4060 4 WL[4]
rlabel metal3 3023 5860 3023 5860 4 WL[6]
rlabel metal3 3023 4960 3023 4960 4 WL[5]
rlabel metal3 4121 6760 4121 6760 4 WL[7]
rlabel metal3 4121 5860 4121 5860 4 WL[6]
rlabel metal3 4121 4960 4121 4960 4 WL[5]
rlabel metal3 3023 4060 3023 4060 4 WL[4]
rlabel metal3 4121 4060 4121 4060 4 WL[4]
rlabel metal3 2423 6760 2423 6760 4 WL[7]
rlabel metal3 2423 5860 2423 5860 4 WL[6]
rlabel metal3 2423 4960 2423 4960 4 WL[5]
rlabel metal3 2423 4060 2423 4060 4 WL[4]
rlabel metal3 s 3066 918 3066 918 4 VSS
rlabel metal3 s 3066 -11 3066 -11 4 VDD
rlabel metal3 s 3666 918 3666 918 4 VSS
rlabel metal3 1823 3160 1823 3160 4 WL[3]
rlabel metal3 s 2934 5 2934 5 4 VDD
rlabel metal3 1823 2260 1823 2260 4 WL[2]
rlabel metal3 1823 1360 1823 1360 4 WL[1]
rlabel metal3 1823 460 1823 460 4 WL[0]
rlabel metal3 1721 460 1721 460 4 WL[0]
rlabel metal3 1721 3160 1721 3160 4 WL[3]
rlabel metal3 2423 1360 2423 1360 4 WL[1]
rlabel metal3 1721 1360 1721 1360 4 WL[1]
rlabel metal3 1721 2260 1721 2260 4 WL[2]
rlabel metal3 s 4134 907 4134 907 4 VSS
rlabel metal3 4121 460 4121 460 4 WL[0]
rlabel metal3 2921 1360 2921 1360 4 WL[1]
rlabel metal3 2921 2260 2921 2260 4 WL[2]
rlabel metal3 4121 3160 4121 3160 4 WL[3]
rlabel metal3 s 1734 5 1734 5 4 VDD
rlabel metal3 s 2934 907 2934 907 4 VSS
rlabel metal3 s 1866 -11 1866 -11 4 VDD
rlabel metal3 s 2466 918 2466 918 4 VSS
rlabel metal3 3623 3160 3623 3160 4 WL[3]
rlabel metal3 3623 2260 3623 2260 4 WL[2]
rlabel metal3 3623 1360 3623 1360 4 WL[1]
rlabel metal3 3623 460 3623 460 4 WL[0]
rlabel metal3 2921 3160 2921 3160 4 WL[3]
rlabel metal3 s 1866 918 1866 918 4 VSS
rlabel metal3 2423 460 2423 460 4 WL[0]
rlabel metal3 4121 2260 4121 2260 4 WL[2]
rlabel metal3 s 4134 5 4134 5 4 VDD
rlabel metal3 s 3666 -11 3666 -11 4 VDD
rlabel metal3 2921 460 2921 460 4 WL[0]
rlabel metal3 3023 3160 3023 3160 4 WL[3]
rlabel metal3 3023 2260 3023 2260 4 WL[2]
rlabel metal3 3023 1360 3023 1360 4 WL[1]
rlabel metal3 3023 460 3023 460 4 WL[0]
rlabel metal3 s 1734 907 1734 907 4 VSS
rlabel metal3 4121 1360 4121 1360 4 WL[1]
rlabel metal3 s 2466 -11 2466 -11 4 VDD
rlabel metal3 2423 3160 2423 3160 4 WL[3]
rlabel metal3 2423 2260 2423 2260 4 WL[2]
rlabel metal3 6079 1360 6079 1360 4 WL[1]
rlabel metal3 6079 460 6079 460 4 WL[0]
rlabel metal3 4223 3160 4223 3160 4 WL[3]
rlabel metal3 4223 2260 4223 2260 4 WL[2]
rlabel metal3 6577 3160 6577 3160 4 WL[3]
rlabel metal3 4223 1360 4223 1360 4 WL[1]
rlabel metal3 s 5334 5 5334 5 4 VDD
rlabel metal3 6577 2260 6577 2260 4 WL[2]
rlabel metal3 6577 1360 6577 1360 4 WL[1]
rlabel metal3 6577 460 6577 460 4 WL[0]
rlabel metal3 s 5334 907 5334 907 4 VSS
rlabel metal3 s 6066 5 6066 5 4 VDD
rlabel metal3 s 4266 -11 4266 -11 4 VDD
rlabel metal3 4223 460 4223 460 4 WL[0]
rlabel metal3 s 4866 -11 4866 -11 4 VDD
rlabel metal3 s 6534 918 6534 918 4 VSS
rlabel metal3 s 4866 918 4866 918 4 VSS
rlabel metal3 4823 2260 4823 2260 4 WL[2]
rlabel metal3 s 4266 918 4266 918 4 VSS
rlabel metal3 5321 3160 5321 3160 4 WL[3]
rlabel metal3 5321 2260 5321 2260 4 WL[2]
rlabel metal3 5321 1360 5321 1360 4 WL[1]
rlabel metal3 5321 460 5321 460 4 WL[0]
rlabel metal3 4823 3160 4823 3160 4 WL[3]
rlabel metal3 s 6066 907 6066 907 4 VSS
rlabel metal3 6079 3160 6079 3160 4 WL[3]
rlabel metal3 s 6534 -11 6534 -11 4 VDD
rlabel metal3 6079 2260 6079 2260 4 WL[2]
rlabel metal3 4823 1360 4823 1360 4 WL[1]
rlabel metal3 4823 460 4823 460 4 WL[0]
rlabel metal3 11423 4060 11423 4060 4 WL[4]
rlabel metal3 10719 4960 10719 4960 4 WL[5]
rlabel metal3 10719 6760 10719 6760 4 WL[7]
rlabel metal3 9577 6760 9577 6760 4 WL[7]
rlabel metal3 9577 5860 9577 5860 4 WL[6]
rlabel metal3 9577 4960 9577 4960 4 WL[5]
rlabel metal3 9577 4060 9577 4060 4 WL[4]
rlabel metal3 11423 4960 11423 4960 4 WL[5]
rlabel metal3 11423 6760 11423 6760 4 WL[7]
rlabel metal3 9679 4060 9679 4060 4 WL[4]
rlabel metal3 9679 4960 9679 4960 4 WL[5]
rlabel metal3 9679 5860 9679 5860 4 WL[6]
rlabel metal3 10177 6760 10177 6760 4 WL[7]
rlabel metal3 10177 5860 10177 5860 4 WL[6]
rlabel metal3 10177 4960 10177 4960 4 WL[5]
rlabel metal3 10177 4060 10177 4060 4 WL[4]
rlabel metal3 10719 4060 10719 4060 4 WL[4]
rlabel metal3 10719 5860 10719 5860 4 WL[6]
rlabel metal3 9679 6760 9679 6760 4 WL[7]
rlabel metal3 11423 5860 11423 5860 4 WL[6]
rlabel metal3 11481 6760 11481 6760 4 WL[7]
rlabel metal3 11481 5860 11481 5860 4 WL[6]
rlabel metal3 11481 4960 11481 4960 4 WL[5]
rlabel metal3 11481 4060 11481 4060 4 WL[4]
rlabel metal3 10777 6760 10777 6760 4 WL[7]
rlabel metal3 10777 5860 10777 5860 4 WL[6]
rlabel metal3 10777 4960 10777 4960 4 WL[5]
rlabel metal3 10777 4060 10777 4060 4 WL[4]
rlabel metal3 7177 4060 7177 4060 4 WL[4]
rlabel metal3 8977 6760 8977 6760 4 WL[7]
rlabel metal3 8977 5860 8977 5860 4 WL[6]
rlabel metal3 8977 4960 8977 4960 4 WL[5]
rlabel metal3 8977 4060 8977 4060 4 WL[4]
rlabel metal3 7777 5860 7777 5860 4 WL[6]
rlabel metal3 7777 4960 7777 4960 4 WL[5]
rlabel metal3 7279 4060 7279 4060 4 WL[4]
rlabel metal3 7279 4960 7279 4960 4 WL[5]
rlabel metal3 7279 5860 7279 5860 4 WL[6]
rlabel metal3 7279 6760 7279 6760 4 WL[7]
rlabel metal3 7777 4060 7777 4060 4 WL[4]
rlabel metal3 8377 5860 8377 5860 4 WL[6]
rlabel metal3 8377 4960 8377 4960 4 WL[5]
rlabel metal3 8377 4060 8377 4060 4 WL[4]
rlabel metal3 8377 6760 8377 6760 4 WL[7]
rlabel metal3 7177 6760 7177 6760 4 WL[7]
rlabel metal3 7177 5860 7177 5860 4 WL[6]
rlabel metal3 7777 6760 7777 6760 4 WL[7]
rlabel metal3 7177 4960 7177 4960 4 WL[5]
rlabel metal3 8479 4060 8479 4060 4 WL[4]
rlabel metal3 8479 4960 8479 4960 4 WL[5]
rlabel metal3 8479 5860 8479 5860 4 WL[6]
rlabel metal3 8479 6760 8479 6760 4 WL[7]
rlabel metal3 8377 460 8377 460 4 WL[0]
rlabel metal3 8977 3160 8977 3160 4 WL[3]
rlabel metal3 8977 2260 8977 2260 4 WL[2]
rlabel metal3 8977 1360 8977 1360 4 WL[1]
rlabel metal3 8977 460 8977 460 4 WL[0]
rlabel metal3 7177 2260 7177 2260 4 WL[2]
rlabel metal3 7177 1360 7177 1360 4 WL[1]
rlabel metal3 s 7734 -11 7734 -11 4 VDD
rlabel metal3 s 8334 918 8334 918 4 VSS
rlabel metal3 s 7266 5 7266 5 4 VDD
rlabel metal3 7177 460 7177 460 4 WL[0]
rlabel metal3 s 7734 918 7734 918 4 VSS
rlabel metal3 7777 3160 7777 3160 4 WL[3]
rlabel metal3 7777 2260 7777 2260 4 WL[2]
rlabel metal3 s 7134 918 7134 918 4 VSS
rlabel metal3 s 7266 907 7266 907 4 VSS
rlabel metal3 8377 3160 8377 3160 4 WL[3]
rlabel metal3 s 8934 -11 8934 -11 4 VDD
rlabel metal3 8377 2260 8377 2260 4 WL[2]
rlabel metal3 s 7134 -11 7134 -11 4 VDD
rlabel metal3 s 8334 -11 8334 -11 4 VDD
rlabel metal3 7777 1360 7777 1360 4 WL[1]
rlabel metal3 7777 460 7777 460 4 WL[0]
rlabel metal3 s 8934 918 8934 918 4 VSS
rlabel metal3 s 8466 907 8466 907 4 VSS
rlabel metal3 s 8466 5 8466 5 4 VDD
rlabel metal3 7279 460 7279 460 4 WL[0]
rlabel metal3 7279 1360 7279 1360 4 WL[1]
rlabel metal3 8479 460 8479 460 4 WL[0]
rlabel metal3 8479 1360 8479 1360 4 WL[1]
rlabel metal3 8479 2260 8479 2260 4 WL[2]
rlabel metal3 8479 3160 8479 3160 4 WL[3]
rlabel metal3 7177 3160 7177 3160 4 WL[3]
rlabel metal3 7279 2260 7279 2260 4 WL[2]
rlabel metal3 7279 3160 7279 3160 4 WL[3]
rlabel metal3 8377 1360 8377 1360 4 WL[1]
rlabel metal3 9679 3160 9679 3160 4 WL[3]
rlabel metal3 11423 2260 11423 2260 4 WL[2]
rlabel metal3 10719 2260 10719 2260 4 WL[2]
rlabel metal3 11423 3160 11423 3160 4 WL[3]
rlabel metal3 10719 3160 10719 3160 4 WL[3]
rlabel metal3 10177 3160 10177 3160 4 WL[3]
rlabel metal3 10177 2260 10177 2260 4 WL[2]
rlabel metal3 10177 1360 10177 1360 4 WL[1]
rlabel metal3 10177 460 10177 460 4 WL[0]
rlabel metal3 s 11466 -11 11466 -11 4 VDD
rlabel metal3 11423 460 11423 460 4 WL[0]
rlabel metal3 s 9534 918 9534 918 4 VSS
rlabel metal3 s 10734 920 10734 920 4 VSS
rlabel metal3 10719 460 10719 460 4 WL[0]
rlabel metal3 11423 1360 11423 1360 4 WL[1]
rlabel metal3 s 9666 907 9666 907 4 VSS
rlabel metal3 s 9666 5 9666 5 4 VDD
rlabel metal3 10719 1360 10719 1360 4 WL[1]
rlabel metal3 s 11466 920 11466 920 4 VSS
rlabel metal3 s 11466 2 11466 2 4 VDD
rlabel metal3 9577 3160 9577 3160 4 WL[3]
rlabel metal3 9577 2260 9577 2260 4 WL[2]
rlabel metal3 11481 3160 11481 3160 4 WL[3]
rlabel metal3 9577 1360 9577 1360 4 WL[1]
rlabel metal3 9577 460 9577 460 4 WL[0]
rlabel metal3 9679 460 9679 460 4 WL[0]
rlabel metal3 9679 1360 9679 1360 4 WL[1]
rlabel metal3 10777 3160 10777 3160 4 WL[3]
rlabel metal3 10777 2260 10777 2260 4 WL[2]
rlabel metal3 10777 1360 10777 1360 4 WL[1]
rlabel metal3 10777 460 10777 460 4 WL[0]
rlabel metal3 9679 2260 9679 2260 4 WL[2]
rlabel metal3 s 10134 -11 10134 -11 4 VDD
rlabel metal3 s 10734 918 10734 918 4 VSS
rlabel metal3 s 9534 -11 9534 -11 4 VDD
rlabel metal3 s 11466 918 11466 918 4 VSS
rlabel metal3 s 10134 918 10134 918 4 VSS
rlabel metal3 11481 1360 11481 1360 4 WL[1]
rlabel metal3 11481 460 11481 460 4 WL[0]
rlabel metal3 11481 2260 11481 2260 4 WL[2]
rlabel metal3 s 10734 -11 10734 -11 4 VDD
rlabel metal3 21519 13060 21519 13060 4 WL[14]
rlabel metal3 21519 13960 21519 13960 4 WL[15]
rlabel metal3 20977 11260 20977 11260 4 WL[12]
rlabel metal3 20977 12160 20977 12160 4 WL[13]
rlabel metal3 20977 13060 20977 13060 4 WL[14]
rlabel metal3 20977 13960 20977 13960 4 WL[15]
rlabel metal3 19177 13960 19177 13960 4 WL[15]
rlabel metal3 19177 13060 19177 13060 4 WL[14]
rlabel metal3 19177 12160 19177 12160 4 WL[13]
rlabel metal3 19177 11260 19177 11260 4 WL[12]
rlabel metal3 21519 11260 21519 11260 4 WL[12]
rlabel metal3 21519 12160 21519 12160 4 WL[13]
rlabel metal3 19777 13960 19777 13960 4 WL[15]
rlabel metal3 19777 13060 19777 13060 4 WL[14]
rlabel metal3 19777 12160 19777 12160 4 WL[13]
rlabel metal3 19777 11260 19777 11260 4 WL[12]
rlabel metal3 21577 13960 21577 13960 4 WL[15]
rlabel metal3 21577 13060 21577 13060 4 WL[14]
rlabel metal3 21577 12160 21577 12160 4 WL[13]
rlabel metal3 21577 11260 21577 11260 4 WL[12]
rlabel metal3 19279 11260 19279 11260 4 WL[12]
rlabel metal3 19279 12160 19279 12160 4 WL[13]
rlabel metal3 19279 13060 19279 13060 4 WL[14]
rlabel metal3 19279 13960 19279 13960 4 WL[15]
rlabel metal3 20479 11260 20479 11260 4 WL[12]
rlabel metal3 20479 12160 20479 12160 4 WL[13]
rlabel metal3 20479 13060 20479 13060 4 WL[14]
rlabel metal3 20479 13960 20479 13960 4 WL[15]
rlabel metal3 20377 13960 20377 13960 4 WL[15]
rlabel metal3 20377 13060 20377 13060 4 WL[14]
rlabel metal3 20377 12160 20377 12160 4 WL[13]
rlabel metal3 20377 11260 20377 11260 4 WL[12]
rlabel metal3 18079 12160 18079 12160 4 WL[13]
rlabel metal3 18079 13060 18079 13060 4 WL[14]
rlabel metal3 18079 13960 18079 13960 4 WL[15]
rlabel metal3 16879 12160 16879 12160 4 WL[13]
rlabel metal3 17977 13060 17977 13060 4 WL[14]
rlabel metal3 17977 13960 17977 13960 4 WL[15]
rlabel metal3 17977 12160 17977 12160 4 WL[13]
rlabel metal3 17977 11260 17977 11260 4 WL[12]
rlabel metal3 16879 13060 16879 13060 4 WL[14]
rlabel metal3 16879 13960 16879 13960 4 WL[15]
rlabel metal3 18577 13960 18577 13960 4 WL[15]
rlabel metal3 18577 13060 18577 13060 4 WL[14]
rlabel metal3 18577 12160 18577 12160 4 WL[13]
rlabel metal3 18577 11260 18577 11260 4 WL[12]
rlabel metal3 16879 11260 16879 11260 4 WL[12]
rlabel metal3 17377 13960 17377 13960 4 WL[15]
rlabel metal3 17377 13060 17377 13060 4 WL[14]
rlabel metal3 17377 12160 17377 12160 4 WL[13]
rlabel metal3 18079 11260 18079 11260 4 WL[12]
rlabel metal3 17377 11260 17377 11260 4 WL[12]
rlabel metal3 18577 10360 18577 10360 4 WL[11]
rlabel metal3 17377 7660 17377 7660 4 WL[8]
rlabel metal3 18577 9460 18577 9460 4 WL[10]
rlabel metal3 17977 10360 17977 10360 4 WL[11]
rlabel metal3 17977 9460 17977 9460 4 WL[10]
rlabel metal3 17977 8560 17977 8560 4 WL[9]
rlabel metal3 17977 7660 17977 7660 4 WL[8]
rlabel metal3 18577 8560 18577 8560 4 WL[9]
rlabel metal3 18577 7660 18577 7660 4 WL[8]
rlabel metal3 17377 9460 17377 9460 4 WL[10]
rlabel metal3 16879 7660 16879 7660 4 WL[8]
rlabel metal3 18079 7660 18079 7660 4 WL[8]
rlabel metal3 18079 8560 18079 8560 4 WL[9]
rlabel metal3 18079 9460 18079 9460 4 WL[10]
rlabel metal3 18079 10360 18079 10360 4 WL[11]
rlabel metal3 16879 8560 16879 8560 4 WL[9]
rlabel metal3 17377 8560 17377 8560 4 WL[9]
rlabel metal3 16879 9460 16879 9460 4 WL[10]
rlabel metal3 16879 10360 16879 10360 4 WL[11]
rlabel metal3 17377 10360 17377 10360 4 WL[11]
rlabel metal3 21577 10360 21577 10360 4 WL[11]
rlabel metal3 21577 9460 21577 9460 4 WL[10]
rlabel metal3 19777 7660 19777 7660 4 WL[8]
rlabel metal3 19177 9460 19177 9460 4 WL[10]
rlabel metal3 21577 7660 21577 7660 4 WL[8]
rlabel metal3 21519 10360 21519 10360 4 WL[11]
rlabel metal3 19177 8560 19177 8560 4 WL[9]
rlabel metal3 19177 7660 19177 7660 4 WL[8]
rlabel metal3 20977 7660 20977 7660 4 WL[8]
rlabel metal3 19777 10360 19777 10360 4 WL[11]
rlabel metal3 19777 9460 19777 9460 4 WL[10]
rlabel metal3 20479 7660 20479 7660 4 WL[8]
rlabel metal3 20479 8560 20479 8560 4 WL[9]
rlabel metal3 20479 9460 20479 9460 4 WL[10]
rlabel metal3 20479 10360 20479 10360 4 WL[11]
rlabel metal3 19777 8560 19777 8560 4 WL[9]
rlabel metal3 19279 7660 19279 7660 4 WL[8]
rlabel metal3 19279 8560 19279 8560 4 WL[9]
rlabel metal3 20977 8560 20977 8560 4 WL[9]
rlabel metal3 20977 9460 20977 9460 4 WL[10]
rlabel metal3 20977 10360 20977 10360 4 WL[11]
rlabel metal3 21519 8560 21519 8560 4 WL[9]
rlabel metal3 19279 9460 19279 9460 4 WL[10]
rlabel metal3 19279 10360 19279 10360 4 WL[11]
rlabel metal3 21519 9460 21519 9460 4 WL[10]
rlabel metal3 19177 10360 19177 10360 4 WL[11]
rlabel metal3 20377 10360 20377 10360 4 WL[11]
rlabel metal3 20377 9460 20377 9460 4 WL[10]
rlabel metal3 20377 8560 20377 8560 4 WL[9]
rlabel metal3 20377 7660 20377 7660 4 WL[8]
rlabel metal3 21519 7660 21519 7660 4 WL[8]
rlabel metal3 21577 8560 21577 8560 4 WL[9]
rlabel metal3 12521 12160 12521 12160 4 WL[13]
rlabel metal3 12521 13060 12521 13060 4 WL[14]
rlabel metal3 13823 7660 13823 7660 4 WL[8]
rlabel metal3 13223 9460 13223 9460 4 WL[10]
rlabel metal3 13223 11260 13223 11260 4 WL[12]
rlabel metal3 13223 13060 13223 13060 4 WL[14]
rlabel metal3 12023 13060 12023 13060 4 WL[14]
rlabel metal3 13721 13960 13721 13960 4 WL[15]
rlabel metal3 12623 11260 12623 11260 4 WL[12]
rlabel metal3 13823 8560 13823 8560 4 WL[9]
rlabel metal3 13721 12160 13721 12160 4 WL[13]
rlabel metal3 12521 9460 12521 9460 4 WL[10]
rlabel metal3 15623 8560 15623 8560 4 WL[9]
rlabel metal3 15623 7660 15623 7660 4 WL[8]
rlabel metal3 12521 7660 12521 7660 4 WL[8]
rlabel metal3 13823 12160 13823 12160 4 WL[13]
rlabel metal3 12623 7660 12623 7660 4 WL[8]
rlabel metal3 13721 7660 13721 7660 4 WL[8]
rlabel metal3 12623 8560 12623 8560 4 WL[9]
rlabel metal3 15023 13960 15023 13960 4 WL[15]
rlabel metal3 15023 13060 15023 13060 4 WL[14]
rlabel metal3 13223 8560 13223 8560 4 WL[9]
rlabel metal3 14921 7660 14921 7660 4 WL[8]
rlabel metal3 14921 8560 14921 8560 4 WL[9]
rlabel metal3 14921 9460 14921 9460 4 WL[10]
rlabel metal3 14921 10360 14921 10360 4 WL[11]
rlabel metal3 14921 11260 14921 11260 4 WL[12]
rlabel metal3 14921 12160 14921 12160 4 WL[13]
rlabel metal3 12023 13960 12023 13960 4 WL[15]
rlabel metal3 13223 10360 13223 10360 4 WL[11]
rlabel metal3 12623 12160 12623 12160 4 WL[13]
rlabel metal3 13223 12160 13223 12160 4 WL[13]
rlabel metal3 13223 13960 13223 13960 4 WL[15]
rlabel metal3 12023 11260 12023 11260 4 WL[12]
rlabel metal3 14423 9460 14423 9460 4 WL[10]
rlabel metal3 14423 7660 14423 7660 4 WL[8]
rlabel metal3 16121 7660 16121 7660 4 WL[8]
rlabel metal3 16121 8560 16121 8560 4 WL[9]
rlabel metal3 16121 9460 16121 9460 4 WL[10]
rlabel metal3 16121 10360 16121 10360 4 WL[11]
rlabel metal3 16121 11260 16121 11260 4 WL[12]
rlabel metal3 16121 12160 16121 12160 4 WL[13]
rlabel metal3 16121 13060 16121 13060 4 WL[14]
rlabel metal3 16121 13960 16121 13960 4 WL[15]
rlabel metal3 15023 12160 15023 12160 4 WL[13]
rlabel metal3 13823 9460 13823 9460 4 WL[10]
rlabel metal3 13823 11260 13823 11260 4 WL[12]
rlabel metal3 14921 13060 14921 13060 4 WL[14]
rlabel metal3 12023 8560 12023 8560 4 WL[9]
rlabel metal3 14921 13960 14921 13960 4 WL[15]
rlabel metal3 13721 13060 13721 13060 4 WL[14]
rlabel metal3 15023 11260 15023 11260 4 WL[12]
rlabel metal3 14423 8560 14423 8560 4 WL[9]
rlabel metal3 14423 10360 14423 10360 4 WL[11]
rlabel metal3 14423 12160 14423 12160 4 WL[13]
rlabel metal3 14423 13960 14423 13960 4 WL[15]
rlabel metal3 15023 10360 15023 10360 4 WL[11]
rlabel metal3 15023 9460 15023 9460 4 WL[10]
rlabel metal3 15023 8560 15023 8560 4 WL[9]
rlabel metal3 15023 7660 15023 7660 4 WL[8]
rlabel metal3 12623 13060 12623 13060 4 WL[14]
rlabel metal3 12023 7660 12023 7660 4 WL[8]
rlabel metal3 12521 13960 12521 13960 4 WL[15]
rlabel metal3 13721 8560 13721 8560 4 WL[9]
rlabel metal3 13823 10360 13823 10360 4 WL[11]
rlabel metal3 12521 10360 12521 10360 4 WL[11]
rlabel metal3 12521 11260 12521 11260 4 WL[12]
rlabel metal3 13721 9460 13721 9460 4 WL[10]
rlabel metal3 13823 13960 13823 13960 4 WL[15]
rlabel metal3 13721 10360 13721 10360 4 WL[11]
rlabel metal3 12023 10360 12023 10360 4 WL[11]
rlabel metal3 13721 11260 13721 11260 4 WL[12]
rlabel metal3 12023 12160 12023 12160 4 WL[13]
rlabel metal3 13823 13060 13823 13060 4 WL[14]
rlabel metal3 12623 10360 12623 10360 4 WL[11]
rlabel metal3 12521 8560 12521 8560 4 WL[9]
rlabel metal3 12623 13960 12623 13960 4 WL[15]
rlabel metal3 15623 13960 15623 13960 4 WL[15]
rlabel metal3 14423 11260 14423 11260 4 WL[12]
rlabel metal3 14423 13060 14423 13060 4 WL[14]
rlabel metal3 15623 13060 15623 13060 4 WL[14]
rlabel metal3 15623 12160 15623 12160 4 WL[13]
rlabel metal3 13223 7660 13223 7660 4 WL[8]
rlabel metal3 15623 11260 15623 11260 4 WL[12]
rlabel metal3 12623 9460 12623 9460 4 WL[10]
rlabel metal3 15623 10360 15623 10360 4 WL[11]
rlabel metal3 15623 9460 15623 9460 4 WL[10]
rlabel metal3 12023 9460 12023 9460 4 WL[10]
rlabel metal3 14921 4060 14921 4060 4 WL[4]
rlabel metal3 15623 5860 15623 5860 4 WL[6]
rlabel metal3 14921 6760 14921 6760 4 WL[7]
rlabel metal3 15623 4960 15623 4960 4 WL[5]
rlabel metal3 15623 6760 15623 6760 4 WL[7]
rlabel metal3 15623 4060 15623 4060 4 WL[4]
rlabel metal3 14921 4960 14921 4960 4 WL[5]
rlabel metal3 14423 4060 14423 4060 4 WL[4]
rlabel metal3 14423 6760 14423 6760 4 WL[7]
rlabel metal3 15023 6760 15023 6760 4 WL[7]
rlabel metal3 15023 5860 15023 5860 4 WL[6]
rlabel metal3 16121 4060 16121 4060 4 WL[4]
rlabel metal3 16121 4960 16121 4960 4 WL[5]
rlabel metal3 16121 5860 16121 5860 4 WL[6]
rlabel metal3 14423 4960 14423 4960 4 WL[5]
rlabel metal3 16121 6760 16121 6760 4 WL[7]
rlabel metal3 15023 4960 15023 4960 4 WL[5]
rlabel metal3 15023 4060 15023 4060 4 WL[4]
rlabel metal3 14423 5860 14423 5860 4 WL[6]
rlabel metal3 14921 5860 14921 5860 4 WL[6]
rlabel metal3 13823 6760 13823 6760 4 WL[7]
rlabel metal3 13823 4060 13823 4060 4 WL[4]
rlabel metal3 13721 6760 13721 6760 4 WL[7]
rlabel metal3 13823 5860 13823 5860 4 WL[6]
rlabel metal3 12023 4960 12023 4960 4 WL[5]
rlabel metal3 12623 5860 12623 5860 4 WL[6]
rlabel metal3 12023 5860 12023 5860 4 WL[6]
rlabel metal3 12623 4060 12623 4060 4 WL[4]
rlabel metal3 12023 6760 12023 6760 4 WL[7]
rlabel metal3 12623 4960 12623 4960 4 WL[5]
rlabel metal3 13721 4060 13721 4060 4 WL[4]
rlabel metal3 13223 4060 13223 4060 4 WL[4]
rlabel metal3 13223 5860 13223 5860 4 WL[6]
rlabel metal3 13823 4960 13823 4960 4 WL[5]
rlabel metal3 13223 6760 13223 6760 4 WL[7]
rlabel metal3 12521 6760 12521 6760 4 WL[7]
rlabel metal3 12521 4060 12521 4060 4 WL[4]
rlabel metal3 12521 4960 12521 4960 4 WL[5]
rlabel metal3 12521 5860 12521 5860 4 WL[6]
rlabel metal3 13721 4960 13721 4960 4 WL[5]
rlabel metal3 13721 5860 13721 5860 4 WL[6]
rlabel metal3 12623 6760 12623 6760 4 WL[7]
rlabel metal3 12023 4060 12023 4060 4 WL[4]
rlabel metal3 13223 4960 13223 4960 4 WL[5]
rlabel metal3 13721 2260 13721 2260 4 WL[2]
rlabel metal3 13721 3160 13721 3160 4 WL[3]
rlabel metal3 12023 460 12023 460 4 WL[0]
rlabel metal3 12521 460 12521 460 4 WL[0]
rlabel metal3 12521 1360 12521 1360 4 WL[1]
rlabel metal3 s 12666 -11 12666 -11 4 VDD
rlabel metal3 12023 1360 12023 1360 4 WL[1]
rlabel metal3 13223 460 13223 460 4 WL[0]
rlabel metal3 13223 2260 13223 2260 4 WL[2]
rlabel metal3 s 13866 -11 13866 -11 4 VDD
rlabel metal3 12623 460 12623 460 4 WL[0]
rlabel metal3 13223 1360 13223 1360 4 WL[1]
rlabel metal3 12521 3160 12521 3160 4 WL[3]
rlabel metal3 s 13734 907 13734 907 4 VSS
rlabel metal3 s 13734 5 13734 5 4 VDD
rlabel metal3 s 13266 -11 13266 -11 4 VDD
rlabel metal3 s 13266 918 13266 918 4 VSS
rlabel metal3 12023 2260 12023 2260 4 WL[2]
rlabel metal3 13721 1360 13721 1360 4 WL[1]
rlabel metal3 12023 3160 12023 3160 4 WL[3]
rlabel metal3 13823 460 13823 460 4 WL[0]
rlabel metal3 s 12534 5 12534 5 4 VDD
rlabel metal3 12623 1360 12623 1360 4 WL[1]
rlabel metal3 12521 2260 12521 2260 4 WL[2]
rlabel metal3 s 13866 918 13866 918 4 VSS
rlabel metal3 13223 3160 13223 3160 4 WL[3]
rlabel metal3 13823 2260 13823 2260 4 WL[2]
rlabel metal3 s 12066 -11 12066 -11 4 VDD
rlabel metal3 13721 460 13721 460 4 WL[0]
rlabel metal3 13823 3160 13823 3160 4 WL[3]
rlabel metal3 s 12066 918 12066 918 4 VSS
rlabel metal3 s 12666 918 12666 918 4 VSS
rlabel metal3 13823 1360 13823 1360 4 WL[1]
rlabel metal3 12623 3160 12623 3160 4 WL[3]
rlabel metal3 12623 2260 12623 2260 4 WL[2]
rlabel metal3 s 12534 907 12534 907 4 VSS
rlabel metal3 14423 460 14423 460 4 WL[0]
rlabel metal3 s 15066 -11 15066 -11 4 VDD
rlabel metal3 14921 2260 14921 2260 4 WL[2]
rlabel metal3 15623 2260 15623 2260 4 WL[2]
rlabel metal3 15623 1360 15623 1360 4 WL[1]
rlabel metal3 15623 460 15623 460 4 WL[0]
rlabel metal3 15023 2260 15023 2260 4 WL[2]
rlabel metal3 16121 460 16121 460 4 WL[0]
rlabel metal3 s 14934 907 14934 907 4 VSS
rlabel metal3 14423 3160 14423 3160 4 WL[3]
rlabel metal3 s 14934 5 14934 5 4 VDD
rlabel metal3 15023 1360 15023 1360 4 WL[1]
rlabel metal3 16121 2260 16121 2260 4 WL[2]
rlabel metal3 s 15666 918 15666 918 4 VSS
rlabel metal3 15023 3160 15023 3160 4 WL[3]
rlabel metal3 14423 1360 14423 1360 4 WL[1]
rlabel metal3 16121 3160 16121 3160 4 WL[3]
rlabel metal3 14921 1360 14921 1360 4 WL[1]
rlabel metal3 16121 1360 16121 1360 4 WL[1]
rlabel metal3 14921 460 14921 460 4 WL[0]
rlabel metal3 s 16134 907 16134 907 4 VSS
rlabel metal3 s 16134 5 16134 5 4 VDD
rlabel metal3 s 15666 -11 15666 -11 4 VDD
rlabel metal3 s 14466 -11 14466 -11 4 VDD
rlabel metal3 s 15066 918 15066 918 4 VSS
rlabel metal3 14921 3160 14921 3160 4 WL[3]
rlabel metal3 15023 460 15023 460 4 WL[0]
rlabel metal3 s 14466 918 14466 918 4 VSS
rlabel metal3 14423 2260 14423 2260 4 WL[2]
rlabel metal3 15623 3160 15623 3160 4 WL[3]
rlabel metal3 21519 6760 21519 6760 4 WL[7]
rlabel metal3 19279 4060 19279 4060 4 WL[4]
rlabel metal3 19279 4960 19279 4960 4 WL[5]
rlabel metal3 19279 5860 19279 5860 4 WL[6]
rlabel metal3 19279 6760 19279 6760 4 WL[7]
rlabel metal3 20977 4960 20977 4960 4 WL[5]
rlabel metal3 21519 5860 21519 5860 4 WL[6]
rlabel metal3 19177 6760 19177 6760 4 WL[7]
rlabel metal3 19177 5860 19177 5860 4 WL[6]
rlabel metal3 19177 4960 19177 4960 4 WL[5]
rlabel metal3 19177 4060 19177 4060 4 WL[4]
rlabel metal3 19777 6760 19777 6760 4 WL[7]
rlabel metal3 21519 4060 21519 4060 4 WL[4]
rlabel metal3 19777 5860 19777 5860 4 WL[6]
rlabel metal3 19777 4960 19777 4960 4 WL[5]
rlabel metal3 19777 4060 19777 4060 4 WL[4]
rlabel metal3 20377 5860 20377 5860 4 WL[6]
rlabel metal3 21577 4960 21577 4960 4 WL[5]
rlabel metal3 20377 4960 20377 4960 4 WL[5]
rlabel metal3 20377 4060 20377 4060 4 WL[4]
rlabel metal3 21577 5860 21577 5860 4 WL[6]
rlabel metal3 20479 4060 20479 4060 4 WL[4]
rlabel metal3 20479 4960 20479 4960 4 WL[5]
rlabel metal3 20479 5860 20479 5860 4 WL[6]
rlabel metal3 20479 6760 20479 6760 4 WL[7]
rlabel metal3 20977 4060 20977 4060 4 WL[4]
rlabel metal3 20977 5860 20977 5860 4 WL[6]
rlabel metal3 21519 4960 21519 4960 4 WL[5]
rlabel metal3 21577 4060 21577 4060 4 WL[4]
rlabel metal3 20977 6760 20977 6760 4 WL[7]
rlabel metal3 21577 6760 21577 6760 4 WL[7]
rlabel metal3 20377 6760 20377 6760 4 WL[7]
rlabel metal3 18577 4960 18577 4960 4 WL[5]
rlabel metal3 17377 6760 17377 6760 4 WL[7]
rlabel metal3 16879 4960 16879 4960 4 WL[5]
rlabel metal3 17377 4060 17377 4060 4 WL[4]
rlabel metal3 16879 5860 16879 5860 4 WL[6]
rlabel metal3 16879 4060 16879 4060 4 WL[4]
rlabel metal3 16879 6760 16879 6760 4 WL[7]
rlabel metal3 17377 5860 17377 5860 4 WL[6]
rlabel metal3 18577 6760 18577 6760 4 WL[7]
rlabel metal3 17977 6760 17977 6760 4 WL[7]
rlabel metal3 18577 4060 18577 4060 4 WL[4]
rlabel metal3 18079 4060 18079 4060 4 WL[4]
rlabel metal3 18079 4960 18079 4960 4 WL[5]
rlabel metal3 18079 5860 18079 5860 4 WL[6]
rlabel metal3 17377 4960 17377 4960 4 WL[5]
rlabel metal3 18079 6760 18079 6760 4 WL[7]
rlabel metal3 17977 5860 17977 5860 4 WL[6]
rlabel metal3 18577 5860 18577 5860 4 WL[6]
rlabel metal3 17977 4960 17977 4960 4 WL[5]
rlabel metal3 17977 4060 17977 4060 4 WL[4]
rlabel metal3 16879 2260 16879 2260 4 WL[2]
rlabel metal3 s 17334 -11 17334 -11 4 VDD
rlabel metal3 17377 3160 17377 3160 4 WL[3]
rlabel metal3 18577 3160 18577 3160 4 WL[3]
rlabel metal3 18577 2260 18577 2260 4 WL[2]
rlabel metal3 17377 460 17377 460 4 WL[0]
rlabel metal3 s 17934 918 17934 918 4 VSS
rlabel metal3 s 18534 918 18534 918 4 VSS
rlabel metal3 s 16866 907 16866 907 4 VSS
rlabel metal3 s 16866 5 16866 5 4 VDD
rlabel metal3 17977 3160 17977 3160 4 WL[3]
rlabel metal3 18577 1360 18577 1360 4 WL[1]
rlabel metal3 18577 460 18577 460 4 WL[0]
rlabel metal3 16879 3160 16879 3160 4 WL[3]
rlabel metal3 17977 1360 17977 1360 4 WL[1]
rlabel metal3 17977 2260 17977 2260 4 WL[2]
rlabel metal3 s 18534 -11 18534 -11 4 VDD
rlabel metal3 s 17334 918 17334 918 4 VSS
rlabel metal3 s 18066 907 18066 907 4 VSS
rlabel metal3 18079 460 18079 460 4 WL[0]
rlabel metal3 18079 1360 18079 1360 4 WL[1]
rlabel metal3 s 17934 -11 17934 -11 4 VDD
rlabel metal3 17377 2260 17377 2260 4 WL[2]
rlabel metal3 17377 1360 17377 1360 4 WL[1]
rlabel metal3 18079 2260 18079 2260 4 WL[2]
rlabel metal3 18079 3160 18079 3160 4 WL[3]
rlabel metal3 s 18066 5 18066 5 4 VDD
rlabel metal3 17977 460 17977 460 4 WL[0]
rlabel metal3 16879 460 16879 460 4 WL[0]
rlabel metal3 16879 1360 16879 1360 4 WL[1]
rlabel metal3 s 19266 5 19266 5 4 VDD
rlabel metal3 20377 460 20377 460 4 WL[0]
rlabel metal3 19177 1360 19177 1360 4 WL[1]
rlabel metal3 s 20934 918 20934 918 4 VSS
rlabel metal3 19177 460 19177 460 4 WL[0]
rlabel metal3 s 20934 -11 20934 -11 4 VDD
rlabel metal3 19279 2260 19279 2260 4 WL[2]
rlabel metal3 20377 2260 20377 2260 4 WL[2]
rlabel metal3 s 21534 918 21534 918 4 VSS
rlabel metal3 s 21534 -11 21534 -11 4 VDD
rlabel metal3 20479 460 20479 460 4 WL[0]
rlabel metal3 20479 1360 20479 1360 4 WL[1]
rlabel metal3 20479 2260 20479 2260 4 WL[2]
rlabel metal3 20479 3160 20479 3160 4 WL[3]
rlabel metal3 19177 3160 19177 3160 4 WL[3]
rlabel metal3 s 19134 918 19134 918 4 VSS
rlabel metal3 s 20466 907 20466 907 4 VSS
rlabel metal3 20977 3160 20977 3160 4 WL[3]
rlabel metal3 s 20466 5 20466 5 4 VDD
rlabel metal3 21519 1360 21519 1360 4 WL[1]
rlabel metal3 21519 3160 21519 3160 4 WL[3]
rlabel metal3 21577 3160 21577 3160 4 WL[3]
rlabel metal3 20377 1360 20377 1360 4 WL[1]
rlabel metal3 19279 3160 19279 3160 4 WL[3]
rlabel metal3 21577 460 21577 460 4 WL[0]
rlabel metal3 21519 460 21519 460 4 WL[0]
rlabel metal3 21577 1360 21577 1360 4 WL[1]
rlabel metal3 s 20334 -11 20334 -11 4 VDD
rlabel metal3 20977 2260 20977 2260 4 WL[2]
rlabel metal3 s 21534 920 21534 920 4 VSS
rlabel metal3 20977 1360 20977 1360 4 WL[1]
rlabel metal3 20977 460 20977 460 4 WL[0]
rlabel metal3 s 19734 -11 19734 -11 4 VDD
rlabel metal3 s 19134 -11 19134 -11 4 VDD
rlabel metal3 19177 2260 19177 2260 4 WL[2]
rlabel metal3 s 19734 918 19734 918 4 VSS
rlabel metal3 s 20334 918 20334 918 4 VSS
rlabel metal3 19279 460 19279 460 4 WL[0]
rlabel metal3 19279 1360 19279 1360 4 WL[1]
rlabel metal3 21577 2260 21577 2260 4 WL[2]
rlabel metal3 21519 2260 21519 2260 4 WL[2]
rlabel metal3 19777 3160 19777 3160 4 WL[3]
rlabel metal3 19777 2260 19777 2260 4 WL[2]
rlabel metal3 19777 1360 19777 1360 4 WL[1]
rlabel metal3 19777 460 19777 460 4 WL[0]
rlabel metal3 20377 3160 20377 3160 4 WL[3]
rlabel metal3 s 19266 907 19266 907 4 VSS
rlabel metal3 s 701 8562 701 8562 4 WL[9]
port 1 nsew
rlabel metal3 s 701 25662 701 25662 4 WL[28]
port 2 nsew
rlabel metal3 s 701 20262 701 20262 4 WL[22]
port 3 nsew
rlabel metal3 s 701 26562 701 26562 4 WL[29]
port 4 nsew
rlabel metal3 s 701 21162 701 21162 4 WL[23]
port 5 nsew
rlabel metal3 s 701 27462 701 27462 4 WL[30]
port 6 nsew
rlabel metal3 s 701 23862 701 23862 4 WL[26]
port 7 nsew
rlabel metal3 s 701 18462 701 18462 4 WL[20]
port 8 nsew
rlabel metal3 s 701 24762 701 24762 4 WL[27]
port 9 nsew
rlabel metal3 s 701 22062 701 22062 4 WL[24]
port 10 nsew
rlabel metal3 s 701 22962 701 22962 4 WL[25]
port 11 nsew
rlabel metal3 s 701 26562 701 26562 4 WL[29]
port 4 nsew
rlabel metal3 s 701 22962 701 22962 4 WL[25]
port 11 nsew
rlabel metal3 s 701 22062 701 22062 4 WL[24]
port 10 nsew
rlabel metal3 s 701 21162 701 21162 4 WL[23]
port 5 nsew
rlabel metal3 s 701 20262 701 20262 4 WL[22]
port 3 nsew
rlabel metal3 s 701 18462 701 18462 4 WL[20]
port 8 nsew
rlabel metal3 s 701 24762 701 24762 4 WL[27]
port 9 nsew
rlabel metal3 s 701 27462 701 27462 4 WL[30]
port 6 nsew
rlabel metal3 s 701 16662 701 16662 4 WL[18]
port 12 nsew
rlabel metal3 s 701 7662 701 7662 4 WL[8]
port 13 nsew
rlabel metal3 s 701 10362 701 10362 4 WL[11]
port 14 nsew
rlabel metal3 s 701 13962 701 13962 4 WL[15]
port 15 nsew
rlabel metal3 s 701 462 701 462 4 WL[0]
port 16 nsew
rlabel metal3 s 701 2262 701 2262 4 WL[2]
port 17 nsew
rlabel metal3 s 701 11262 701 11262 4 WL[12]
port 18 nsew
rlabel metal3 s 701 9462 701 9462 4 WL[10]
port 19 nsew
rlabel metal3 s 701 10362 701 10362 4 WL[11]
port 14 nsew
rlabel metal3 s 701 5862 701 5862 4 WL[6]
port 20 nsew
rlabel metal3 s 701 4062 701 4062 4 WL[4]
port 21 nsew
rlabel metal3 s 701 3162 701 3162 4 WL[3]
port 22 nsew
rlabel metal3 s 701 4062 701 4062 4 WL[4]
port 21 nsew
rlabel metal3 s 701 13062 701 13062 4 WL[14]
port 23 nsew
rlabel metal3 s 701 16662 701 16662 4 WL[18]
port 12 nsew
rlabel metal3 s 701 11262 701 11262 4 WL[12]
port 18 nsew
rlabel metal3 s 701 4962 701 4962 4 WL[5]
port 24 nsew
rlabel metal3 s 701 5862 701 5862 4 WL[6]
port 20 nsew
rlabel metal3 s 701 17562 701 17562 4 WL[19]
port 25 nsew
rlabel metal3 s 701 6762 701 6762 4 WL[7]
port 26 nsew
rlabel metal3 s 701 7662 701 7662 4 WL[8]
port 13 nsew
rlabel metal3 s 701 8562 701 8562 4 WL[9]
port 1 nsew
rlabel metal3 s 701 1362 701 1362 4 WL[1]
port 27 nsew
rlabel metal3 s 701 28362 701 28362 4 WL[31]
port 28 nsew
rlabel metal3 s 701 9462 701 9462 4 WL[10]
port 19 nsew
rlabel metal3 s 701 12162 701 12162 4 WL[13]
port 29 nsew
rlabel metal3 s 701 13062 701 13062 4 WL[14]
port 23 nsew
rlabel metal3 s 701 14862 701 14862 4 WL[16]
port 30 nsew
rlabel metal3 s 701 15762 701 15762 4 WL[17]
port 31 nsew
rlabel metal3 s 701 23862 701 23862 4 WL[26]
port 7 nsew
rlabel metal3 s 701 17562 701 17562 4 WL[19]
port 25 nsew
rlabel metal3 s 701 25662 701 25662 4 WL[28]
port 2 nsew
rlabel metal3 s 701 19362 701 19362 4 WL[21]
port 32 nsew
rlabel metal3 s 701 13962 701 13962 4 WL[15]
port 15 nsew
rlabel metal3 s 701 1362 701 1362 4 WL[1]
port 27 nsew
rlabel metal3 s 701 462 701 462 4 WL[0]
port 16 nsew
rlabel metal3 s 701 2262 701 2262 4 WL[2]
port 17 nsew
rlabel metal3 s 701 3162 701 3162 4 WL[3]
port 22 nsew
rlabel metal3 s 701 4962 701 4962 4 WL[5]
port 24 nsew
rlabel metal3 s 701 28362 701 28362 4 WL[31]
port 28 nsew
rlabel metal3 s 701 12162 701 12162 4 WL[13]
port 29 nsew
rlabel metal3 s 701 14862 701 14862 4 WL[16]
port 30 nsew
rlabel metal3 s 701 19362 701 19362 4 WL[21]
port 32 nsew
rlabel metal3 s 701 15762 701 15762 4 WL[17]
port 31 nsew
rlabel metal3 s 701 6762 701 6762 4 WL[7]
port 26 nsew
<< properties >>
string GDS_END 2046258
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1924278
<< end >>
