magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 355 3222 870
rect -86 352 952 355
rect 1550 352 3222 355
<< pwell >>
rect 952 352 1550 355
rect -86 -86 3222 352
<< mvnmos >>
rect 124 137 244 216
rect 348 137 468 216
rect 572 137 692 216
rect 799 137 919 216
rect 1059 156 1179 235
rect 1315 156 1435 235
rect 1815 91 1935 169
rect 2039 91 2159 169
rect 2407 91 2527 169
rect 2591 91 2711 169
rect 2851 91 2971 217
<< mvpmos >>
rect 144 475 244 660
rect 348 475 448 660
rect 588 507 688 660
rect 887 507 987 660
rect 1127 475 1227 628
rect 1335 475 1435 628
rect 1809 475 1909 659
rect 2014 475 2114 659
rect 2407 472 2507 656
rect 2611 472 2711 656
rect 2851 472 2951 716
<< mvndiff >>
rect 979 216 1059 235
rect 36 199 124 216
rect 36 153 49 199
rect 95 153 124 199
rect 36 137 124 153
rect 244 199 348 216
rect 244 153 273 199
rect 319 153 348 199
rect 244 137 348 153
rect 468 199 572 216
rect 468 153 497 199
rect 543 153 572 199
rect 468 137 572 153
rect 692 199 799 216
rect 692 153 721 199
rect 767 153 799 199
rect 692 137 799 153
rect 919 156 1059 216
rect 1179 215 1315 235
rect 1179 169 1224 215
rect 1270 169 1315 215
rect 1179 156 1315 169
rect 1435 215 1523 235
rect 1435 169 1464 215
rect 1510 169 1523 215
rect 2771 169 2851 217
rect 1435 156 1523 169
rect 919 137 999 156
rect 1727 152 1815 169
rect 1727 106 1740 152
rect 1786 106 1815 152
rect 1727 91 1815 106
rect 1935 152 2039 169
rect 1935 106 1964 152
rect 2010 106 2039 152
rect 1935 91 2039 106
rect 2159 152 2247 169
rect 2159 106 2188 152
rect 2234 106 2247 152
rect 2159 91 2247 106
rect 2319 152 2407 169
rect 2319 106 2332 152
rect 2378 106 2407 152
rect 2319 91 2407 106
rect 2527 91 2591 169
rect 2711 150 2851 169
rect 2711 104 2740 150
rect 2786 104 2851 150
rect 2711 91 2851 104
rect 2971 189 3059 217
rect 2971 143 3000 189
rect 3046 143 3059 189
rect 2971 91 3059 143
<< mvpdiff >>
rect 56 647 144 660
rect 56 507 69 647
rect 115 507 144 647
rect 56 475 144 507
rect 244 475 348 660
rect 448 507 588 660
rect 688 614 887 660
rect 688 568 762 614
rect 808 568 887 614
rect 688 507 887 568
rect 987 628 1067 660
rect 987 507 1127 628
rect 448 475 528 507
rect 1047 475 1127 507
rect 1227 615 1335 628
rect 1227 569 1260 615
rect 1306 569 1335 615
rect 1227 475 1335 569
rect 1435 544 1523 628
rect 1435 498 1464 544
rect 1510 498 1523 544
rect 1435 475 1523 498
rect 1721 559 1809 659
rect 1721 513 1734 559
rect 1780 513 1809 559
rect 1721 475 1809 513
rect 1909 641 2014 659
rect 1909 595 1938 641
rect 1984 595 2014 641
rect 1909 475 2014 595
rect 2114 559 2202 659
rect 2771 656 2851 716
rect 2114 513 2143 559
rect 2189 513 2202 559
rect 2114 475 2202 513
rect 2314 643 2407 656
rect 2314 503 2327 643
rect 2373 503 2407 643
rect 2314 472 2407 503
rect 2507 639 2611 656
rect 2507 499 2536 639
rect 2582 499 2611 639
rect 2507 472 2611 499
rect 2711 640 2851 656
rect 2711 594 2740 640
rect 2786 594 2851 640
rect 2711 472 2851 594
rect 2951 625 3039 716
rect 2951 485 2980 625
rect 3026 485 3039 625
rect 2951 472 3039 485
<< mvndiffc >>
rect 49 153 95 199
rect 273 153 319 199
rect 497 153 543 199
rect 721 153 767 199
rect 1224 169 1270 215
rect 1464 169 1510 215
rect 1740 106 1786 152
rect 1964 106 2010 152
rect 2188 106 2234 152
rect 2332 106 2378 152
rect 2740 104 2786 150
rect 3000 143 3046 189
<< mvpdiffc >>
rect 69 507 115 647
rect 762 568 808 614
rect 1260 569 1306 615
rect 1464 498 1510 544
rect 1734 513 1780 559
rect 1938 595 1984 641
rect 2143 513 2189 559
rect 2327 503 2373 643
rect 2536 499 2582 639
rect 2740 594 2786 640
rect 2980 485 3026 625
<< polysilicon >>
rect 887 720 1909 760
rect 144 660 244 704
rect 348 660 448 704
rect 588 660 688 704
rect 887 660 987 720
rect 1127 628 1227 672
rect 1335 628 1435 672
rect 1809 659 1909 720
rect 2851 716 2951 760
rect 2014 659 2114 706
rect 144 415 244 475
rect 144 369 159 415
rect 205 369 244 415
rect 144 260 244 369
rect 124 216 244 260
rect 348 415 448 475
rect 348 369 387 415
rect 433 369 448 415
rect 588 447 688 507
rect 588 407 839 447
rect 348 260 448 369
rect 572 346 751 359
rect 572 300 692 346
rect 738 300 751 346
rect 572 287 751 300
rect 348 216 468 260
rect 572 216 692 287
rect 799 260 839 407
rect 887 420 987 507
rect 2407 656 2507 703
rect 2611 656 2711 703
rect 887 374 913 420
rect 959 374 987 420
rect 887 361 987 374
rect 1127 407 1227 475
rect 1127 361 1150 407
rect 1196 361 1227 407
rect 1127 348 1227 361
rect 1127 279 1179 348
rect 1335 314 1435 475
rect 1335 279 1355 314
rect 799 216 919 260
rect 1059 235 1179 279
rect 1315 268 1355 279
rect 1401 268 1435 314
rect 1315 235 1435 268
rect 1809 411 1909 475
rect 1809 365 1850 411
rect 1896 365 1909 411
rect 1809 286 1909 365
rect 1809 240 1850 286
rect 1896 240 1909 286
rect 1809 229 1909 240
rect 2014 353 2114 475
rect 2014 307 2054 353
rect 2100 307 2114 353
rect 2014 229 2114 307
rect 1815 214 1909 229
rect 2039 214 2114 229
rect 2407 303 2507 472
rect 2407 257 2425 303
rect 2471 257 2507 303
rect 1815 169 1935 214
rect 2039 169 2159 214
rect 2407 213 2507 257
rect 2611 439 2711 472
rect 2611 393 2626 439
rect 2672 393 2711 439
rect 2611 213 2711 393
rect 2851 394 2951 472
rect 2851 348 2864 394
rect 2910 348 2951 394
rect 2851 288 2951 348
rect 2851 217 2971 288
rect 2407 169 2527 213
rect 2591 169 2711 213
rect 124 93 244 137
rect 348 93 468 137
rect 572 93 692 137
rect 799 64 919 137
rect 1059 112 1179 156
rect 1315 112 1435 156
rect 1583 152 1655 165
rect 1583 106 1596 152
rect 1642 106 1655 152
rect 1583 64 1655 106
rect 799 24 1655 64
rect 1815 46 1935 91
rect 2039 46 2159 91
rect 2407 47 2527 91
rect 2591 47 2711 91
rect 2851 44 2971 91
<< polycontact >>
rect 159 369 205 415
rect 387 369 433 415
rect 692 300 738 346
rect 913 374 959 420
rect 1150 361 1196 407
rect 1355 268 1401 314
rect 1850 365 1896 411
rect 1850 240 1896 286
rect 2054 307 2100 353
rect 2425 257 2471 303
rect 2626 393 2672 439
rect 2864 348 2910 394
rect 1596 106 1642 152
<< metal1 >>
rect 0 724 3136 844
rect 69 647 115 724
rect 69 496 115 507
rect 468 430 550 674
rect 762 614 808 625
rect 1249 615 1317 724
rect 1249 569 1260 615
rect 1306 569 1317 615
rect 1464 632 1879 678
rect 762 512 808 568
rect 1464 544 1510 632
rect 58 415 318 430
rect 58 369 159 415
rect 205 369 318 415
rect 58 354 318 369
rect 373 415 550 430
rect 373 369 387 415
rect 433 369 550 415
rect 373 354 550 369
rect 600 466 1087 512
rect 38 245 423 292
rect 38 199 106 245
rect 377 199 423 245
rect 600 199 646 466
rect 692 374 913 420
rect 959 374 987 420
rect 692 346 738 374
rect 692 289 738 300
rect 1041 315 1087 466
rect 1464 407 1510 498
rect 1729 559 1786 570
rect 1729 513 1734 559
rect 1780 513 1786 559
rect 1729 407 1786 513
rect 1833 538 1879 632
rect 1938 641 1984 724
rect 1938 584 1984 595
rect 2040 632 2281 678
rect 2040 538 2086 632
rect 1833 491 2086 538
rect 2143 559 2189 570
rect 2143 445 2189 513
rect 1137 361 1150 407
rect 1196 361 1510 407
rect 1041 314 1416 315
rect 1041 268 1355 314
rect 1401 268 1416 314
rect 1464 215 1510 361
rect 38 153 49 199
rect 95 153 106 199
rect 262 153 273 199
rect 319 153 330 199
rect 377 153 497 199
rect 543 153 554 199
rect 600 153 721 199
rect 767 153 778 199
rect 1213 169 1224 215
rect 1270 169 1281 215
rect 262 60 330 153
rect 1213 60 1281 169
rect 1464 156 1510 169
rect 1583 361 1786 407
rect 1849 411 2189 445
rect 1849 365 1850 411
rect 1896 399 2189 411
rect 2235 445 2281 632
rect 2327 643 2373 724
rect 2327 492 2373 503
rect 2536 639 2582 650
rect 2740 640 2786 724
rect 2740 580 2786 594
rect 2832 625 3046 654
rect 2582 499 2775 534
rect 2536 488 2775 499
rect 2235 442 2453 445
rect 2235 439 2683 442
rect 2235 399 2626 439
rect 1896 365 1897 399
rect 2402 393 2626 399
rect 2672 393 2683 439
rect 2729 405 2775 488
rect 2832 485 2980 625
rect 3026 485 3046 625
rect 2832 466 3046 485
rect 2729 394 2910 405
rect 1583 152 1655 361
rect 1849 286 1897 365
rect 2043 307 2054 353
rect 2100 318 2213 353
rect 2729 348 2864 394
rect 2729 337 2910 348
rect 2100 307 2551 318
rect 2729 307 2775 337
rect 1849 240 1850 286
rect 1896 261 1897 286
rect 2157 303 2551 307
rect 1896 240 2102 261
rect 2157 257 2425 303
rect 2471 257 2551 303
rect 2157 242 2551 257
rect 2602 253 2775 307
rect 1849 215 2102 240
rect 1964 152 2010 169
rect 1583 106 1596 152
rect 1642 106 1740 152
rect 1786 106 1815 152
rect 2056 152 2102 215
rect 2602 152 2648 253
rect 2956 224 3046 466
rect 2940 189 3046 224
rect 2056 106 2188 152
rect 2234 106 2247 152
rect 2319 106 2332 152
rect 2378 106 2648 152
rect 2740 150 2786 161
rect 1964 60 2010 106
rect 2940 143 3000 189
rect 2940 112 3046 143
rect 2740 60 2786 104
rect 0 -60 3136 60
<< labels >>
flabel metal1 s 2832 466 3046 654 0 FreeSans 400 0 0 0 Q
port 4 nsew default output
flabel metal1 s 58 354 318 430 0 FreeSans 400 0 0 0 TE
port 3 nsew default input
flabel metal1 s 0 724 3136 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1213 199 1281 215 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 2043 318 2213 353 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel metal1 s 468 430 550 674 0 FreeSans 400 0 0 0 E
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 2043 307 2551 318 1 CLK
port 1 nsew clock input
rlabel metal1 s 2157 242 2551 307 1 CLK
port 1 nsew clock input
rlabel metal1 s 373 354 550 430 1 E
port 2 nsew default input
rlabel metal1 s 2956 224 3046 466 1 Q
port 4 nsew default output
rlabel metal1 s 2940 112 3046 224 1 Q
port 4 nsew default output
rlabel metal1 s 2740 584 2786 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 584 2373 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1938 584 1984 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1249 584 1317 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 584 115 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2740 580 2786 584 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 580 2373 584 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1249 580 1317 584 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 580 115 584 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 569 2373 580 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1249 569 1317 580 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 569 115 580 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 496 2373 569 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 496 115 569 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 492 2373 496 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1213 169 1281 199 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 169 330 199 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1964 161 2010 169 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1213 161 1281 169 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 161 330 169 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2740 60 2786 161 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1964 60 2010 161 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1213 60 1281 161 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 161 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3136 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3136 784
string GDS_END 458006
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 450740
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
