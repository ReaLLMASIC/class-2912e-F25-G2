magic
tech gf180mcuD
timestamp 1749799538
<< properties >>
string gencell npn_00p54x10p00_0
string library gf180mcu
string parameter m=1
<< end >>
