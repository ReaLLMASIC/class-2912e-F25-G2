magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 453 982 1094
<< pwell >>
rect -86 -86 982 453
<< mvnmos >>
rect 124 126 244 272
rect 348 126 468 272
rect 572 126 692 272
<< mvpmos >>
rect 124 573 224 939
rect 348 573 448 939
rect 572 573 672 939
<< mvndiff >>
rect 36 193 124 272
rect 36 147 49 193
rect 95 147 124 193
rect 36 126 124 147
rect 244 193 348 272
rect 244 147 273 193
rect 319 147 348 193
rect 244 126 348 147
rect 468 185 572 272
rect 468 139 497 185
rect 543 139 572 185
rect 468 126 572 139
rect 692 193 780 272
rect 692 147 721 193
rect 767 147 780 193
rect 692 126 780 147
<< mvpdiff >>
rect 36 861 124 939
rect 36 721 49 861
rect 95 721 124 861
rect 36 573 124 721
rect 224 861 348 939
rect 224 721 273 861
rect 319 721 348 861
rect 224 573 348 721
rect 448 861 572 939
rect 448 721 477 861
rect 523 721 572 861
rect 448 573 572 721
rect 672 861 760 939
rect 672 721 701 861
rect 747 721 760 861
rect 672 573 760 721
<< mvndiffc >>
rect 49 147 95 193
rect 273 147 319 193
rect 497 139 543 185
rect 721 147 767 193
<< mvpdiffc >>
rect 49 721 95 861
rect 273 721 319 861
rect 477 721 523 861
rect 701 721 747 861
<< polysilicon >>
rect 124 939 224 983
rect 348 939 448 983
rect 572 939 672 983
rect 124 513 224 573
rect 348 513 448 573
rect 572 513 672 573
rect 124 500 672 513
rect 124 454 137 500
rect 465 454 672 500
rect 124 441 672 454
rect 124 272 244 441
rect 348 272 468 441
rect 572 316 672 441
rect 572 272 692 316
rect 124 82 244 126
rect 348 82 468 126
rect 572 82 692 126
<< polycontact >>
rect 137 454 465 500
<< metal1 >>
rect 0 918 896 1098
rect 49 861 95 918
rect 49 710 95 721
rect 273 861 319 872
rect 273 664 319 721
rect 477 861 523 918
rect 477 710 523 721
rect 701 861 767 872
rect 747 721 767 861
rect 701 664 767 721
rect 273 618 767 664
rect 137 500 465 542
rect 137 443 465 454
rect 366 354 418 443
rect 702 288 767 618
rect 273 242 767 288
rect 49 193 95 204
rect 49 90 95 147
rect 273 193 319 242
rect 273 136 319 147
rect 497 185 543 196
rect 497 90 543 139
rect 721 193 767 242
rect 721 136 767 147
rect 0 -90 896 90
<< labels >>
flabel metal1 s 137 443 465 542 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 896 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 49 196 95 204 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 701 664 767 872 0 FreeSans 200 0 0 0 ZN
port 2 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 366 354 418 443 1 I
port 1 nsew default input
rlabel metal1 s 273 664 319 872 1 ZN
port 2 nsew default output
rlabel metal1 s 273 618 767 664 1 ZN
port 2 nsew default output
rlabel metal1 s 702 288 767 618 1 ZN
port 2 nsew default output
rlabel metal1 s 273 242 767 288 1 ZN
port 2 nsew default output
rlabel metal1 s 721 136 767 242 1 ZN
port 2 nsew default output
rlabel metal1 s 273 136 319 242 1 ZN
port 2 nsew default output
rlabel metal1 s 477 710 523 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 497 90 543 196 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 196 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 896 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 896 1008
string GDS_END 1449310
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1446280
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
