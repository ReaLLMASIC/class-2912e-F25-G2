magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 352 1430 870
<< pwell >>
rect -86 -86 1430 352
<< metal1 >>
rect 0 724 1344 844
rect 244 428 312 676
rect 168 346 312 428
rect 358 322 428 676
rect 580 322 652 676
rect 743 506 789 724
rect 968 531 1092 676
rect 1185 587 1231 724
rect 968 476 1208 531
rect 1149 307 1208 476
rect 974 253 1208 307
rect 273 60 319 179
rect 721 60 767 179
rect 974 106 1098 253
rect 1205 60 1251 184
rect 0 -60 1344 60
<< obsm1 >>
rect 49 272 115 678
rect 792 353 1103 399
rect 792 272 838 353
rect 49 225 838 272
rect 49 106 95 225
rect 497 106 543 225
<< labels >>
rlabel metal1 s 168 346 312 428 6 A1
port 1 nsew default input
rlabel metal1 s 244 428 312 676 6 A1
port 1 nsew default input
rlabel metal1 s 358 322 428 676 6 A2
port 2 nsew default input
rlabel metal1 s 580 322 652 676 6 A3
port 3 nsew default input
rlabel metal1 s 974 106 1098 253 6 Z
port 4 nsew default output
rlabel metal1 s 974 253 1208 307 6 Z
port 4 nsew default output
rlabel metal1 s 1149 307 1208 476 6 Z
port 4 nsew default output
rlabel metal1 s 968 476 1208 531 6 Z
port 4 nsew default output
rlabel metal1 s 968 531 1092 676 6 Z
port 4 nsew default output
rlabel metal1 s 1185 587 1231 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 743 506 789 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 724 1344 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel nwell s -86 352 1430 870 6 VNW
port 6 nsew power bidirectional
rlabel pwell s -86 -86 1430 352 6 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 0 -60 1344 60 8 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1205 60 1251 184 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 721 60 767 179 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 179 6 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1344 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 162208
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 158400
<< end >>
