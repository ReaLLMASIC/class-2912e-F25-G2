magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 377 4006 870
rect -86 352 219 377
rect 2916 352 4006 377
<< pwell >>
rect -86 -86 4006 352
<< mvnmos >>
rect 124 68 244 232
rect 392 93 512 257
rect 616 93 736 257
rect 840 93 960 257
rect 1064 93 1184 257
rect 1288 93 1408 257
rect 1512 93 1632 257
rect 1736 93 1856 257
rect 1960 93 2080 257
rect 2184 93 2304 257
rect 2408 93 2528 257
rect 2632 93 2752 257
rect 2960 68 3080 232
rect 3184 68 3304 232
rect 3408 68 3528 232
rect 3632 68 3752 232
<< mvpmos >>
rect 144 497 244 716
rect 392 497 492 716
rect 636 497 736 716
rect 840 497 940 716
rect 1084 497 1184 716
rect 1308 497 1408 716
rect 1512 497 1612 716
rect 1756 497 1856 716
rect 1960 497 2060 716
rect 2204 497 2304 716
rect 2408 497 2508 716
rect 2632 497 2732 716
rect 2980 497 3080 716
rect 3184 497 3284 716
rect 3428 497 3528 716
rect 3632 497 3732 716
<< mvndiff >>
rect 304 244 392 257
rect 304 232 317 244
rect 36 152 124 232
rect 36 106 49 152
rect 95 106 124 152
rect 36 68 124 106
rect 244 198 317 232
rect 363 198 392 244
rect 244 93 392 198
rect 512 152 616 257
rect 512 106 541 152
rect 587 106 616 152
rect 512 93 616 106
rect 736 244 840 257
rect 736 198 765 244
rect 811 198 840 244
rect 736 93 840 198
rect 960 152 1064 257
rect 960 106 989 152
rect 1035 106 1064 152
rect 960 93 1064 106
rect 1184 244 1288 257
rect 1184 198 1213 244
rect 1259 198 1288 244
rect 1184 93 1288 198
rect 1408 152 1512 257
rect 1408 106 1437 152
rect 1483 106 1512 152
rect 1408 93 1512 106
rect 1632 244 1736 257
rect 1632 198 1661 244
rect 1707 198 1736 244
rect 1632 93 1736 198
rect 1856 152 1960 257
rect 1856 106 1885 152
rect 1931 106 1960 152
rect 1856 93 1960 106
rect 2080 244 2184 257
rect 2080 198 2109 244
rect 2155 198 2184 244
rect 2080 93 2184 198
rect 2304 152 2408 257
rect 2304 106 2333 152
rect 2379 106 2408 152
rect 2304 93 2408 106
rect 2528 244 2632 257
rect 2528 198 2557 244
rect 2603 198 2632 244
rect 2528 93 2632 198
rect 2752 232 2832 257
rect 2752 152 2960 232
rect 2752 106 2885 152
rect 2931 106 2960 152
rect 2752 93 2960 106
rect 244 68 324 93
rect 2812 68 2960 93
rect 3080 127 3184 232
rect 3080 81 3109 127
rect 3155 81 3184 127
rect 3080 68 3184 81
rect 3304 219 3408 232
rect 3304 173 3333 219
rect 3379 173 3408 219
rect 3304 68 3408 173
rect 3528 127 3632 232
rect 3528 81 3557 127
rect 3603 81 3632 127
rect 3528 68 3632 81
rect 3752 219 3840 232
rect 3752 173 3781 219
rect 3827 173 3840 219
rect 3752 68 3840 173
<< mvpdiff >>
rect 56 665 144 716
rect 56 525 69 665
rect 115 525 144 665
rect 56 497 144 525
rect 244 703 392 716
rect 244 657 317 703
rect 363 657 392 703
rect 244 497 392 657
rect 492 665 636 716
rect 492 525 541 665
rect 587 525 636 665
rect 492 497 636 525
rect 736 703 840 716
rect 736 657 765 703
rect 811 657 840 703
rect 736 497 840 657
rect 940 497 1084 716
rect 1184 497 1308 716
rect 1408 586 1512 716
rect 1408 540 1437 586
rect 1483 540 1512 586
rect 1408 497 1512 540
rect 1612 497 1756 716
rect 1856 678 1960 716
rect 1856 632 1885 678
rect 1931 632 1960 678
rect 1856 497 1960 632
rect 2060 497 2204 716
rect 2304 586 2408 716
rect 2304 540 2333 586
rect 2379 540 2408 586
rect 2304 497 2408 540
rect 2508 497 2632 716
rect 2732 678 2820 716
rect 2732 632 2761 678
rect 2807 632 2820 678
rect 2732 497 2820 632
rect 2892 703 2980 716
rect 2892 657 2905 703
rect 2951 657 2980 703
rect 2892 497 2980 657
rect 3080 586 3184 716
rect 3080 540 3109 586
rect 3155 540 3184 586
rect 3080 497 3184 540
rect 3284 703 3428 716
rect 3284 657 3333 703
rect 3379 657 3428 703
rect 3284 497 3428 657
rect 3528 586 3632 716
rect 3528 540 3557 586
rect 3603 540 3632 586
rect 3528 497 3632 540
rect 3732 665 3830 716
rect 3732 525 3771 665
rect 3817 525 3830 665
rect 3732 497 3830 525
<< mvndiffc >>
rect 49 106 95 152
rect 317 198 363 244
rect 541 106 587 152
rect 765 198 811 244
rect 989 106 1035 152
rect 1213 198 1259 244
rect 1437 106 1483 152
rect 1661 198 1707 244
rect 1885 106 1931 152
rect 2109 198 2155 244
rect 2333 106 2379 152
rect 2557 198 2603 244
rect 2885 106 2931 152
rect 3109 81 3155 127
rect 3333 173 3379 219
rect 3557 81 3603 127
rect 3781 173 3827 219
<< mvpdiffc >>
rect 69 525 115 665
rect 317 657 363 703
rect 541 525 587 665
rect 765 657 811 703
rect 1437 540 1483 586
rect 1885 632 1931 678
rect 2333 540 2379 586
rect 2761 632 2807 678
rect 2905 657 2951 703
rect 3109 540 3155 586
rect 3333 657 3379 703
rect 3557 540 3603 586
rect 3771 525 3817 665
<< polysilicon >>
rect 144 716 244 760
rect 392 716 492 760
rect 636 716 736 760
rect 840 716 940 760
rect 1084 716 1184 760
rect 1308 716 1408 760
rect 1512 716 1612 760
rect 1756 716 1856 760
rect 1960 716 2060 760
rect 2204 716 2304 760
rect 2408 716 2508 760
rect 2632 716 2732 760
rect 2980 716 3080 760
rect 3184 716 3284 760
rect 3428 716 3528 760
rect 3632 716 3732 760
rect 144 408 244 497
rect 392 408 492 497
rect 636 408 736 497
rect 840 408 940 497
rect 1084 433 1184 497
rect 124 395 960 408
rect 1084 402 1111 433
rect 124 349 161 395
rect 207 349 265 395
rect 311 349 369 395
rect 415 349 473 395
rect 519 349 577 395
rect 623 349 960 395
rect 124 336 960 349
rect 124 232 244 336
rect 392 257 512 336
rect 616 257 736 336
rect 840 257 960 336
rect 1064 387 1111 402
rect 1157 387 1184 433
rect 1308 402 1408 497
rect 1064 257 1184 387
rect 1288 394 1408 402
rect 1512 402 1612 497
rect 1756 433 1856 497
rect 1756 402 1783 433
rect 1512 394 1632 402
rect 1288 348 1632 394
rect 1288 336 1408 348
rect 1288 290 1325 336
rect 1371 290 1408 336
rect 1288 257 1408 290
rect 1512 336 1632 348
rect 1512 290 1549 336
rect 1595 290 1632 336
rect 1512 257 1632 290
rect 1736 387 1783 402
rect 1829 394 1856 433
rect 1960 433 2060 497
rect 1960 394 1987 433
rect 1829 387 1987 394
rect 2033 402 2060 433
rect 2204 402 2304 497
rect 2033 387 2080 402
rect 1736 348 2080 387
rect 1736 257 1856 348
rect 1960 257 2080 348
rect 2184 394 2304 402
rect 2408 402 2508 497
rect 2632 433 2732 497
rect 2408 394 2528 402
rect 2184 348 2528 394
rect 2184 336 2304 348
rect 2184 290 2221 336
rect 2267 290 2304 336
rect 2184 257 2304 290
rect 2408 336 2528 348
rect 2408 290 2427 336
rect 2473 290 2528 336
rect 2408 257 2528 290
rect 2632 387 2651 433
rect 2697 402 2732 433
rect 2980 415 3080 497
rect 2980 402 3007 415
rect 2697 387 2752 402
rect 2632 257 2752 387
rect 2960 369 3007 402
rect 3053 402 3080 415
rect 3184 415 3284 497
rect 3184 402 3211 415
rect 3053 369 3211 402
rect 3257 402 3284 415
rect 3428 415 3528 497
rect 3428 402 3455 415
rect 3257 369 3455 402
rect 3501 402 3528 415
rect 3632 415 3732 497
rect 3632 402 3659 415
rect 3501 369 3659 402
rect 3705 402 3732 415
rect 3705 369 3752 402
rect 2960 348 3752 369
rect 2960 232 3080 348
rect 3184 232 3304 348
rect 3408 232 3528 348
rect 3632 232 3752 348
rect 124 24 244 68
rect 392 24 512 93
rect 616 24 736 93
rect 840 24 960 93
rect 1064 24 1184 93
rect 1288 24 1408 93
rect 1512 24 1632 93
rect 1736 24 1856 93
rect 1960 24 2080 93
rect 2184 24 2304 93
rect 2408 24 2528 93
rect 2632 24 2752 93
rect 2960 24 3080 68
rect 3184 24 3304 68
rect 3408 24 3528 68
rect 3632 24 3752 68
<< polycontact >>
rect 161 349 207 395
rect 265 349 311 395
rect 369 349 415 395
rect 473 349 519 395
rect 577 349 623 395
rect 1111 387 1157 433
rect 1325 290 1371 336
rect 1549 290 1595 336
rect 1783 387 1829 433
rect 1987 387 2033 433
rect 2221 290 2267 336
rect 2427 290 2473 336
rect 2651 387 2697 433
rect 3007 369 3053 415
rect 3211 369 3257 415
rect 3455 369 3501 415
rect 3659 369 3705 415
<< metal1 >>
rect 0 724 3920 844
rect 306 703 374 724
rect 69 665 115 676
rect 306 657 317 703
rect 363 657 374 703
rect 754 703 822 724
rect 541 665 587 676
rect 115 525 541 560
rect 754 657 765 703
rect 811 657 822 703
rect 2894 703 2962 724
rect 872 632 1885 678
rect 1931 632 2761 678
rect 2807 632 2820 678
rect 2894 657 2905 703
rect 2951 657 2962 703
rect 3322 703 3390 724
rect 3322 657 3333 703
rect 3379 657 3390 703
rect 3771 665 3817 724
rect 872 560 918 632
rect 587 525 918 560
rect 69 514 918 525
rect 1030 490 1355 542
rect 1426 540 1437 586
rect 1483 540 2333 586
rect 2379 540 3109 586
rect 3155 540 3557 586
rect 3603 540 3686 586
rect 1030 444 2778 490
rect 1084 433 1184 444
rect 124 395 648 430
rect 124 349 161 395
rect 207 349 265 395
rect 311 349 369 395
rect 415 349 473 395
rect 519 349 577 395
rect 623 349 648 395
rect 696 354 984 430
rect 1084 387 1111 433
rect 1157 387 1184 433
rect 1084 382 1184 387
rect 1772 433 2044 444
rect 1772 387 1783 433
rect 1829 387 1987 433
rect 2033 387 2044 433
rect 1772 382 2044 387
rect 2594 433 2778 444
rect 2594 387 2651 433
rect 2697 387 2778 433
rect 124 336 648 349
rect 938 336 984 354
rect 2594 345 2778 387
rect 2824 472 3686 540
rect 3771 514 3817 525
rect 938 290 1325 336
rect 1371 290 1549 336
rect 1595 290 2221 336
rect 2267 290 2427 336
rect 2473 290 2484 336
rect 2824 244 2888 472
rect 2978 415 3830 424
rect 2978 369 3007 415
rect 3053 369 3211 415
rect 3257 369 3455 415
rect 3501 369 3659 415
rect 3705 369 3830 415
rect 2978 357 3830 369
rect 262 198 317 244
rect 363 198 765 244
rect 811 198 1213 244
rect 1259 198 1661 244
rect 1707 198 2109 244
rect 2155 198 2557 244
rect 2603 198 2888 244
rect 2996 173 3333 219
rect 3379 173 3781 219
rect 3827 173 3840 219
rect 2996 152 3042 173
rect 36 106 49 152
rect 95 106 541 152
rect 587 106 989 152
rect 1035 106 1437 152
rect 1483 106 1885 152
rect 1931 106 2333 152
rect 2379 106 2885 152
rect 2931 106 3042 152
rect 3098 81 3109 127
rect 3155 81 3166 127
rect 3098 60 3166 81
rect 3546 81 3557 127
rect 3603 81 3614 127
rect 3546 60 3614 81
rect 0 -60 3920 60
<< labels >>
flabel metal1 s 124 336 648 430 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 2978 357 3830 424 0 FreeSans 400 0 0 0 B
port 4 nsew default input
flabel metal1 s 0 724 3920 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 3546 60 3614 127 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 1426 540 3686 586 0 FreeSans 400 0 0 0 ZN
port 5 nsew default output
flabel metal1 s 696 354 984 430 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1030 490 1355 542 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 938 336 984 354 1 A1
port 1 nsew default input
rlabel metal1 s 938 290 2484 336 1 A1
port 1 nsew default input
rlabel metal1 s 1030 444 2778 490 1 A2
port 2 nsew default input
rlabel metal1 s 2594 382 2778 444 1 A2
port 2 nsew default input
rlabel metal1 s 1772 382 2044 444 1 A2
port 2 nsew default input
rlabel metal1 s 1084 382 1184 444 1 A2
port 2 nsew default input
rlabel metal1 s 2594 345 2778 382 1 A2
port 2 nsew default input
rlabel metal1 s 2824 472 3686 540 1 ZN
port 5 nsew default output
rlabel metal1 s 2824 244 2888 472 1 ZN
port 5 nsew default output
rlabel metal1 s 262 198 2888 244 1 ZN
port 5 nsew default output
rlabel metal1 s 3771 657 3817 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3322 657 3390 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2894 657 2962 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 754 657 822 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 306 657 374 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3771 514 3817 657 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3098 60 3166 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3920 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3920 784
string GDS_END 51476
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 44342
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
