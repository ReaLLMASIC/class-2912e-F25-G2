magic
tech gf180mcuD
magscale 1 10
timestamp 1749760379
<< nwell >>
rect -86 352 1654 870
<< pwell >>
rect -86 -86 1654 352
<< metal1 >>
rect 0 724 1568 844
rect 69 518 115 724
rect 165 588 768 647
rect 165 450 211 588
rect 29 404 211 450
rect 261 476 1326 531
rect 1373 526 1419 724
rect 29 223 84 404
rect 261 333 316 476
rect 387 354 542 419
rect 591 365 878 419
rect 141 278 316 333
rect 477 318 542 354
rect 925 354 1130 430
rect 925 318 979 354
rect 1250 346 1326 476
rect 477 272 979 318
rect 29 177 1450 223
rect 29 106 106 177
rect 260 60 332 131
rect 378 106 662 177
rect 708 60 780 131
rect 826 106 1110 177
rect 1156 60 1228 131
rect 1381 106 1450 177
rect 0 -60 1568 60
<< labels >>
rlabel metal1 s 591 365 878 419 6 A1
port 1 nsew default input
rlabel metal1 s 477 272 979 318 6 A2
port 2 nsew default input
rlabel metal1 s 925 318 979 354 6 A2
port 2 nsew default input
rlabel metal1 s 925 354 1130 430 6 A2
port 2 nsew default input
rlabel metal1 s 477 318 542 354 6 A2
port 2 nsew default input
rlabel metal1 s 387 354 542 419 6 A2
port 2 nsew default input
rlabel metal1 s 141 278 316 333 6 A3
port 3 nsew default input
rlabel metal1 s 1250 346 1326 476 6 A3
port 3 nsew default input
rlabel metal1 s 261 333 316 476 6 A3
port 3 nsew default input
rlabel metal1 s 261 476 1326 531 6 A3
port 3 nsew default input
rlabel metal1 s 1381 106 1450 177 6 ZN
port 4 nsew default output
rlabel metal1 s 826 106 1110 177 6 ZN
port 4 nsew default output
rlabel metal1 s 378 106 662 177 6 ZN
port 4 nsew default output
rlabel metal1 s 29 106 106 177 6 ZN
port 4 nsew default output
rlabel metal1 s 29 177 1450 223 6 ZN
port 4 nsew default output
rlabel metal1 s 29 223 84 404 6 ZN
port 4 nsew default output
rlabel metal1 s 29 404 211 450 6 ZN
port 4 nsew default output
rlabel metal1 s 165 450 211 588 6 ZN
port 4 nsew default output
rlabel metal1 s 165 588 768 647 6 ZN
port 4 nsew default output
rlabel metal1 s 1373 526 1419 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 518 115 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 724 1568 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel nwell s -86 352 1654 870 6 VNW
port 6 nsew power bidirectional
rlabel pwell s -86 -86 1654 352 6 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 0 -60 1568 60 8 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1156 60 1228 131 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 708 60 780 131 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 260 60 332 131 6 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1568 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 754848
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 750976
<< end >>
